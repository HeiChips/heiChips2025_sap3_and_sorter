* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_lgcp_1 abstract view
.subckt sg13g2_lgcp_1 GATE CLK GCLK VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
X_3155_ VPWR VGND _0677_ _0682_ _1703_ _1607_ _0683_ _1622_ sg13g2_a221oi_1
X_3086_ _0603_ _0605_ _0608_ _0613_ _0614_ VPWR VGND sg13g2_nor4_1
X_2106_ net774 net772 _1526_ VPWR VGND sg13g2_nor2_1
XFILLER_27_428 VPWR VGND sg13g2_fill_1
X_2037_ VPWR _1459_ net805 VGND sg13g2_inv_1
XFILLER_36_962 VPWR VGND sg13g2_decap_8
XFILLER_23_645 VPWR VGND sg13g2_decap_8
X_3988_ _1402_ sap_3_inst.alu.act\[3\] net582 VPWR VGND sg13g2_nand2_1
XFILLER_11_818 VPWR VGND sg13g2_decap_8
X_2939_ VGND VPWR net796 _1473_ _0495_ _0462_ sg13g2_a21oi_1
Xfanout831 net832 net831 VPWR VGND sg13g2_buf_8
Xfanout820 net822 net820 VPWR VGND sg13g2_buf_8
Xfanout842 net845 net842 VPWR VGND sg13g2_buf_8
XFILLER_46_737 VPWR VGND sg13g2_decap_8
XFILLER_27_973 VPWR VGND sg13g2_decap_8
XFILLER_26_450 VPWR VGND sg13g2_decap_8
XFILLER_42_954 VPWR VGND sg13g2_decap_8
XFILLER_14_667 VPWR VGND sg13g2_decap_8
XFILLER_41_497 VPWR VGND sg13g2_decap_8
XFILLER_13_177 VPWR VGND sg13g2_fill_1
XFILLER_10_851 VPWR VGND sg13g2_decap_8
XFILLER_6_866 VPWR VGND sg13g2_decap_8
XFILLER_49_575 VPWR VGND sg13g2_decap_8
XFILLER_37_737 VPWR VGND sg13g2_decap_8
XFILLER_18_973 VPWR VGND sg13g2_decap_8
XFILLER_45_781 VPWR VGND sg13g2_decap_8
XFILLER_33_910 VPWR VGND sg13g2_decap_8
XFILLER_17_494 VPWR VGND sg13g2_decap_8
X_3911_ _1341_ VPWR _0163_ VGND _1502_ _0154_ sg13g2_o21ai_1
X_3842_ _1281_ _1278_ _1280_ VPWR VGND sg13g2_nand2_1
XFILLER_33_987 VPWR VGND sg13g2_decap_8
XFILLER_20_626 VPWR VGND sg13g2_decap_8
X_3773_ _1184_ net613 net713 _1234_ VPWR VGND sg13g2_a21o_1
XFILLER_8_170 VPWR VGND sg13g2_fill_2
X_2724_ _0295_ _0294_ _1601_ _0291_ _0290_ VPWR VGND sg13g2_a22oi_1
XFILLER_9_693 VPWR VGND sg13g2_decap_8
X_2655_ _0242_ net629 _0241_ VPWR VGND sg13g2_nand2_1
X_2586_ VGND VPWR _1996_ net628 net802 sg13g2_or2_1
X_3207_ _0735_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] net677 VPWR
+ VGND sg13g2_nand2_1
X_4187_ net824 VGND VPWR _0151_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\]
+ clknet_5_10__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3138_ VPWR _0666_ net676 VGND sg13g2_inv_1
XFILLER_43_707 VPWR VGND sg13g2_decap_8
X_3069_ net738 net32 _0601_ VPWR VGND sg13g2_nor2_1
XFILLER_24_965 VPWR VGND sg13g2_decap_8
XFILLER_11_615 VPWR VGND sg13g2_decap_8
XFILLER_23_442 VPWR VGND sg13g2_decap_8
XFILLER_6_129 VPWR VGND sg13g2_fill_2
XFILLER_5_4 VPWR VGND sg13g2_decap_4
XFILLER_3_869 VPWR VGND sg13g2_decap_8
Xfanout650 _1800_ net650 VPWR VGND sg13g2_buf_8
Xfanout672 net673 net672 VPWR VGND sg13g2_buf_1
Xfanout683 _0338_ net683 VPWR VGND sg13g2_buf_8
Xfanout661 net662 net661 VPWR VGND sg13g2_buf_8
Xfanout694 net695 net694 VPWR VGND sg13g2_buf_2
XFILLER_46_534 VPWR VGND sg13g2_decap_8
XFILLER_19_759 VPWR VGND sg13g2_decap_8
XFILLER_15_910 VPWR VGND sg13g2_decap_8
XFILLER_27_770 VPWR VGND sg13g2_decap_8
XFILLER_42_751 VPWR VGND sg13g2_decap_8
XFILLER_15_987 VPWR VGND sg13g2_decap_8
XFILLER_18_1015 VPWR VGND sg13g2_decap_8
XFILLER_30_968 VPWR VGND sg13g2_decap_8
XFILLER_6_663 VPWR VGND sg13g2_decap_8
X_2440_ _1860_ _1809_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\] net637
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_184 VPWR VGND sg13g2_fill_1
X_2371_ _1742_ _1790_ net756 _1791_ VPWR VGND sg13g2_nand3_1
X_4110_ net843 VGND VPWR _0074_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\]
+ clknet_5_27__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_49_372 VPWR VGND sg13g2_decap_8
XFILLER_37_534 VPWR VGND sg13g2_decap_8
XFILLER_18_770 VPWR VGND sg13g2_decap_8
XFILLER_25_729 VPWR VGND sg13g2_decap_8
XFILLER_21_935 VPWR VGND sg13g2_decap_8
XFILLER_33_784 VPWR VGND sg13g2_decap_8
X_3825_ net13 net608 _1269_ VPWR VGND sg13g2_nor2_1
X_3756_ net711 VPWR _1219_ VGND net651 _0898_ sg13g2_o21ai_1
X_2707_ _1644_ _0284_ _0286_ _0004_ VPWR VGND sg13g2_nor3_1
XFILLER_9_490 VPWR VGND sg13g2_decap_8
X_3687_ _1046_ _1047_ net579 _1175_ VPWR VGND sg13g2_nor3_1
X_2638_ _0218_ _0226_ _0214_ net18 VPWR VGND sg13g2_nand3_1
X_2569_ VGND VPWR net577 _1980_ _1981_ _1973_ sg13g2_a21oi_1
X_4239_ regFile_serial net29 VPWR VGND sg13g2_buf_8
XFILLER_28_567 VPWR VGND sg13g2_decap_8
XFILLER_43_504 VPWR VGND sg13g2_decap_8
XFILLER_24_762 VPWR VGND sg13g2_decap_8
XFILLER_12_924 VPWR VGND sg13g2_decap_8
XFILLER_11_489 VPWR VGND sg13g2_decap_8
XFILLER_20_990 VPWR VGND sg13g2_decap_8
XFILLER_3_666 VPWR VGND sg13g2_decap_8
XFILLER_2_143 VPWR VGND sg13g2_fill_1
XFILLER_47_865 VPWR VGND sg13g2_decap_8
XFILLER_19_556 VPWR VGND sg13g2_decap_8
XFILLER_15_784 VPWR VGND sg13g2_decap_8
XFILLER_30_765 VPWR VGND sg13g2_decap_8
X_3610_ _0088_ _1110_ _1115_ net619 _1492_ VPWR VGND sg13g2_a22oi_1
XFILLER_7_950 VPWR VGND sg13g2_decap_8
X_3541_ net32 _0850_ _1057_ VPWR VGND sg13g2_nor2_1
X_3472_ _0993_ _0994_ net651 _0995_ VPWR VGND sg13g2_mux2_1
X_2423_ _1597_ _1646_ net777 _1843_ VPWR VGND sg13g2_nand3_1
X_2354_ net736 _1717_ net774 _1774_ VPWR VGND sg13g2_nand3_1
XFILLER_29_0 VPWR VGND sg13g2_fill_1
X_2285_ _1575_ net726 _1705_ VPWR VGND sg13g2_nor2_1
XFILLER_38_821 VPWR VGND sg13g2_decap_8
X_4024_ _1429_ net74 _0189_ VPWR VGND sg13g2_xor2_1
XFILLER_38_898 VPWR VGND sg13g2_decap_8
XFILLER_25_526 VPWR VGND sg13g2_decap_8
XFILLER_21_732 VPWR VGND sg13g2_decap_8
XFILLER_33_581 VPWR VGND sg13g2_decap_8
X_3808_ VGND VPWR _1486_ net612 _0144_ _1257_ sg13g2_a21oi_1
X_3739_ _1177_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] net593 _0123_
+ VPWR VGND sg13g2_mux2_1
XFILLER_0_647 VPWR VGND sg13g2_decap_8
XFILLER_29_832 VPWR VGND sg13g2_decap_8
XFILLER_44_813 VPWR VGND sg13g2_decap_8
XFILLER_31_507 VPWR VGND sg13g2_decap_8
XFILLER_43_378 VPWR VGND sg13g2_decap_8
XFILLER_12_721 VPWR VGND sg13g2_decap_8
XFILLER_8_747 VPWR VGND sg13g2_decap_8
XFILLER_12_798 VPWR VGND sg13g2_decap_8
XFILLER_7_246 VPWR VGND sg13g2_fill_1
XFILLER_4_942 VPWR VGND sg13g2_decap_8
XFILLER_39_607 VPWR VGND sg13g2_decap_8
X_2070_ VPWR _1492_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_47_662 VPWR VGND sg13g2_decap_8
XFILLER_35_857 VPWR VGND sg13g2_decap_8
X_2972_ VGND VPWR _0489_ _0525_ _0527_ _0328_ sg13g2_a21oi_1
XFILLER_15_581 VPWR VGND sg13g2_decap_8
XFILLER_30_562 VPWR VGND sg13g2_decap_8
X_3524_ _0700_ net596 _1044_ VPWR VGND sg13g2_and2_1
X_3455_ _0930_ _0953_ _0908_ _0978_ VPWR VGND _0977_ sg13g2_nand4_1
X_2406_ VGND VPWR _1826_ _1825_ net777 sg13g2_or2_1
X_3386_ _0912_ _0910_ net586 VPWR VGND sg13g2_nand2b_1
X_2337_ _1757_ _1747_ net736 _1705_ _1593_ VPWR VGND sg13g2_a22oi_1
X_2268_ _1688_ _1686_ _1687_ _1604_ net735 VPWR VGND sg13g2_a22oi_1
XFILLER_44_109 VPWR VGND sg13g2_fill_2
X_4007_ _1416_ u_ser.bit_pos\[1\] net814 VPWR VGND sg13g2_nand2_1
X_2199_ _1525_ _1562_ _1444_ _1619_ VPWR VGND sg13g2_nand3_1
XFILLER_26_835 VPWR VGND sg13g2_decap_8
XFILLER_38_695 VPWR VGND sg13g2_decap_8
XFILLER_41_805 VPWR VGND sg13g2_decap_8
XFILLER_13_529 VPWR VGND sg13g2_decap_8
XFILLER_5_728 VPWR VGND sg13g2_decap_8
XFILLER_1_934 VPWR VGND sg13g2_decap_8
Xhold30 u_ser.bit_pos\[0\] VPWR VGND net79 sg13g2_dlygate4sd3_1
XFILLER_48_437 VPWR VGND sg13g2_decap_8
XFILLER_17_802 VPWR VGND sg13g2_decap_8
XFILLER_44_610 VPWR VGND sg13g2_decap_8
XFILLER_16_345 VPWR VGND sg13g2_fill_2
XFILLER_17_879 VPWR VGND sg13g2_decap_8
XFILLER_44_687 VPWR VGND sg13g2_decap_8
XFILLER_31_304 VPWR VGND sg13g2_fill_1
XFILLER_25_890 VPWR VGND sg13g2_decap_8
XFILLER_8_544 VPWR VGND sg13g2_decap_8
XFILLER_12_595 VPWR VGND sg13g2_decap_8
X_3240_ net703 net690 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] _0768_
+ VPWR VGND sg13g2_nand3_1
XFILLER_6_1027 VPWR VGND sg13g2_fill_2
X_3171_ net704 net701 net693 net688 _0699_ VPWR VGND sg13g2_nor4_1
X_2122_ net779 _1444_ net786 net783 _1542_ VPWR VGND sg13g2_nor4_1
X_2053_ VPWR _1475_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_35_654 VPWR VGND sg13g2_decap_8
XFILLER_23_827 VPWR VGND sg13g2_decap_8
X_2955_ sap_3_inst.alu.tmp\[6\] net790 _0510_ VPWR VGND sg13g2_xor2_1
XFILLER_31_871 VPWR VGND sg13g2_decap_8
X_2886_ net580 net799 _0443_ _0036_ VPWR VGND sg13g2_a21o_1
X_3507_ _1028_ _0992_ _1007_ _1027_ VPWR VGND sg13g2_and3_1
X_3438_ _0962_ _0936_ _0953_ VPWR VGND sg13g2_xnor2_1
X_3369_ _0896_ _0843_ _0883_ VPWR VGND sg13g2_xnor2_1
XFILLER_46_919 VPWR VGND sg13g2_decap_8
XFILLER_39_971 VPWR VGND sg13g2_decap_8
XFILLER_26_632 VPWR VGND sg13g2_decap_8
XFILLER_38_492 VPWR VGND sg13g2_decap_8
XFILLER_41_602 VPWR VGND sg13g2_decap_8
XFILLER_14_849 VPWR VGND sg13g2_decap_8
XFILLER_13_348 VPWR VGND sg13g2_fill_1
XFILLER_41_679 VPWR VGND sg13g2_decap_8
XFILLER_22_860 VPWR VGND sg13g2_decap_8
XFILLER_5_525 VPWR VGND sg13g2_decap_8
Xoutput20 net20 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_731 VPWR VGND sg13g2_decap_8
XFILLER_49_757 VPWR VGND sg13g2_decap_8
XFILLER_37_919 VPWR VGND sg13g2_decap_8
XFILLER_45_963 VPWR VGND sg13g2_decap_8
XFILLER_44_484 VPWR VGND sg13g2_decap_8
XFILLER_17_676 VPWR VGND sg13g2_decap_8
XFILLER_32_657 VPWR VGND sg13g2_decap_8
XFILLER_20_808 VPWR VGND sg13g2_decap_8
X_2740_ VGND VPWR _1549_ _1717_ _0301_ _1551_ sg13g2_a21oi_1
XFILLER_13_893 VPWR VGND sg13g2_decap_8
XFILLER_9_875 VPWR VGND sg13g2_decap_8
X_2671_ _0253_ _0256_ _1868_ _0257_ VPWR VGND sg13g2_nand3_1
X_3223_ net698 net694 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] _0751_
+ VPWR VGND net689 sg13g2_nand4_1
X_3154_ _0679_ _0680_ _1787_ _0682_ VPWR VGND _0681_ sg13g2_nand4_1
X_3085_ _0609_ _0611_ _1770_ _0613_ VPWR VGND _0612_ sg13g2_nand4_1
X_2105_ net785 net782 _1525_ VPWR VGND sg13g2_nor2_2
X_2036_ _1458_ net803 VPWR VGND sg13g2_inv_2
XFILLER_36_941 VPWR VGND sg13g2_decap_8
XFILLER_23_624 VPWR VGND sg13g2_decap_8
X_3987_ VGND VPWR _0434_ net709 _1401_ _1400_ sg13g2_a21oi_1
XFILLER_10_329 VPWR VGND sg13g2_fill_2
X_2938_ VPWR VGND net790 _0493_ net682 net796 _0494_ net683 sg13g2_a221oi_1
XFILLER_11_1021 VPWR VGND sg13g2_decap_8
X_2869_ _0427_ _0400_ _0426_ VPWR VGND sg13g2_nand2_2
XFILLER_2_539 VPWR VGND sg13g2_decap_8
Xfanout843 net844 net843 VPWR VGND sg13g2_buf_8
Xfanout832 net835 net832 VPWR VGND sg13g2_buf_8
Xfanout821 net822 net821 VPWR VGND sg13g2_buf_8
Xfanout810 _1304_ net810 VPWR VGND sg13g2_buf_8
XFILLER_46_716 VPWR VGND sg13g2_decap_8
XFILLER_45_237 VPWR VGND sg13g2_fill_1
XFILLER_27_952 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_42_933 VPWR VGND sg13g2_decap_8
XFILLER_41_421 VPWR VGND sg13g2_fill_1
XFILLER_14_646 VPWR VGND sg13g2_decap_8
XFILLER_41_476 VPWR VGND sg13g2_decap_8
XFILLER_10_830 VPWR VGND sg13g2_decap_8
XFILLER_6_845 VPWR VGND sg13g2_decap_8
XFILLER_49_554 VPWR VGND sg13g2_decap_8
XFILLER_37_716 VPWR VGND sg13g2_decap_8
XFILLER_18_952 VPWR VGND sg13g2_decap_8
XFILLER_45_760 VPWR VGND sg13g2_decap_8
XFILLER_44_281 VPWR VGND sg13g2_fill_2
X_3910_ _1339_ _1333_ _1340_ _1341_ VPWR VGND sg13g2_a21o_1
XFILLER_20_605 VPWR VGND sg13g2_decap_8
X_3841_ _1280_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\] _1279_ VPWR
+ VGND sg13g2_nand2_1
XFILLER_33_966 VPWR VGND sg13g2_decap_8
X_3772_ _0937_ _1232_ net651 _1233_ VPWR VGND sg13g2_mux2_1
X_2723_ net744 _1683_ _0293_ _0294_ VPWR VGND sg13g2_or3_1
XFILLER_13_690 VPWR VGND sg13g2_decap_8
XFILLER_9_672 VPWR VGND sg13g2_decap_8
X_2654_ _0241_ sap_3_inst.alu.flags\[0\] _1839_ VPWR VGND sg13g2_nand2_1
X_2585_ VGND VPWR _1995_ _1994_ _1723_ sg13g2_or2_1
X_3206_ _0734_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] net674 VPWR
+ VGND sg13g2_nand2_1
X_4186_ net842 VGND VPWR _0150_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\]
+ clknet_5_30__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_749 VPWR VGND sg13g2_decap_8
X_3137_ _0665_ net705 net699 _0658_ VPWR VGND sg13g2_and3_1
X_3068_ _0600_ VPWR _0061_ VGND net738 net572 sg13g2_o21ai_1
X_2019_ net777 _1441_ VPWR VGND sg13g2_inv_4
XFILLER_23_421 VPWR VGND sg13g2_decap_8
XFILLER_24_944 VPWR VGND sg13g2_decap_8
XFILLER_10_115 VPWR VGND sg13g2_fill_2
XFILLER_23_498 VPWR VGND sg13g2_decap_8
XFILLER_3_848 VPWR VGND sg13g2_decap_8
Xfanout651 _0821_ net651 VPWR VGND sg13g2_buf_8
Xfanout640 net641 net640 VPWR VGND sg13g2_buf_8
Xfanout684 net685 net684 VPWR VGND sg13g2_buf_8
Xfanout662 _0702_ net662 VPWR VGND sg13g2_buf_8
Xfanout673 _0692_ net673 VPWR VGND sg13g2_buf_8
XFILLER_46_513 VPWR VGND sg13g2_decap_8
XFILLER_19_738 VPWR VGND sg13g2_decap_8
Xfanout695 net696 net695 VPWR VGND sg13g2_buf_1
XFILLER_37_52 VPWR VGND sg13g2_fill_2
XFILLER_42_730 VPWR VGND sg13g2_decap_8
XFILLER_15_966 VPWR VGND sg13g2_decap_8
XFILLER_30_947 VPWR VGND sg13g2_decap_8
XFILLER_6_642 VPWR VGND sg13g2_decap_8
X_2370_ net745 net763 net777 _1790_ VPWR VGND _1549_ sg13g2_nand4_1
XFILLER_25_1009 VPWR VGND sg13g2_decap_8
XFILLER_49_351 VPWR VGND sg13g2_decap_8
XFILLER_37_513 VPWR VGND sg13g2_decap_8
XFILLER_25_708 VPWR VGND sg13g2_decap_8
XFILLER_21_914 VPWR VGND sg13g2_decap_8
XFILLER_33_763 VPWR VGND sg13g2_decap_8
XFILLER_20_446 VPWR VGND sg13g2_fill_2
X_3824_ _1268_ VPWR _0149_ VGND _1447_ net655 sg13g2_o21ai_1
X_3755_ net614 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] _1218_ _0130_
+ VPWR VGND sg13g2_a21o_1
X_2706_ VGND VPWR sap_3_inst.controller.stage\[2\] _1507_ _0286_ sap_3_inst.controller.stage\[3\]
+ sg13g2_a21oi_1
X_3686_ net677 _1137_ _1174_ VPWR VGND sg13g2_nor2_2
X_2637_ net576 VPWR _0226_ VGND _0221_ _0225_ sg13g2_o21ai_1
XFILLER_0_829 VPWR VGND sg13g2_decap_8
X_2568_ _1977_ _1979_ _1976_ _1980_ VPWR VGND sg13g2_nand3_1
X_2499_ _1913_ net639 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] net641
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4238_ sap_3_outputReg_start_sync net28 VPWR VGND sg13g2_buf_1
X_4169_ net821 VGND VPWR _0133_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\]
+ clknet_5_7__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_546 VPWR VGND sg13g2_decap_8
XFILLER_12_903 VPWR VGND sg13g2_decap_8
XFILLER_24_741 VPWR VGND sg13g2_decap_8
XFILLER_8_929 VPWR VGND sg13g2_decap_8
Xclkbuf_4_12_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_12_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_3_645 VPWR VGND sg13g2_decap_8
XFILLER_47_844 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_fill_2
XFILLER_19_535 VPWR VGND sg13g2_decap_8
XFILLER_46_387 VPWR VGND sg13g2_decap_8
XFILLER_34_549 VPWR VGND sg13g2_decap_8
XFILLER_9_12 VPWR VGND sg13g2_fill_2
XFILLER_15_763 VPWR VGND sg13g2_decap_8
XFILLER_30_744 VPWR VGND sg13g2_decap_8
X_3540_ VGND VPWR _1453_ net584 _0077_ _1056_ sg13g2_a21oi_1
X_3471_ _0994_ _0955_ _0977_ VPWR VGND sg13g2_xnor2_1
X_2422_ _1530_ VPWR _1842_ VGND _1517_ net729 sg13g2_o21ai_1
X_2353_ _1773_ _1772_ _1637_ _1767_ _1625_ VPWR VGND sg13g2_a22oi_1
X_2284_ _1575_ _1639_ _1704_ VPWR VGND sg13g2_nor2_1
X_4023_ _1440_ _1285_ _1429_ VPWR VGND sg13g2_nor2_2
XFILLER_38_800 VPWR VGND sg13g2_decap_8
XFILLER_25_505 VPWR VGND sg13g2_decap_8
XFILLER_38_877 VPWR VGND sg13g2_decap_8
XFILLER_21_711 VPWR VGND sg13g2_decap_8
XFILLER_33_560 VPWR VGND sg13g2_decap_8
XFILLER_20_210 VPWR VGND sg13g2_fill_2
X_3807_ net612 _1066_ _1132_ _1257_ VPWR VGND sg13g2_nor3_1
XFILLER_21_788 VPWR VGND sg13g2_decap_8
X_3738_ net593 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] _1209_ _0122_
+ VPWR VGND sg13g2_a21o_1
X_3669_ net623 _1158_ _1159_ _1160_ VPWR VGND sg13g2_or3_1
XFILLER_0_626 VPWR VGND sg13g2_decap_8
Xclkbuf_4_4_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_4_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_48_619 VPWR VGND sg13g2_decap_8
XFILLER_29_811 VPWR VGND sg13g2_decap_8
XFILLER_28_332 VPWR VGND sg13g2_fill_1
XFILLER_29_888 VPWR VGND sg13g2_decap_8
XFILLER_16_549 VPWR VGND sg13g2_decap_8
XFILLER_44_869 VPWR VGND sg13g2_decap_8
XFILLER_12_700 VPWR VGND sg13g2_decap_8
XFILLER_15_1008 VPWR VGND sg13g2_decap_8
XFILLER_8_726 VPWR VGND sg13g2_decap_8
XFILLER_7_203 VPWR VGND sg13g2_fill_1
XFILLER_12_777 VPWR VGND sg13g2_decap_8
XFILLER_4_921 VPWR VGND sg13g2_decap_8
XFILLER_4_998 VPWR VGND sg13g2_decap_8
XFILLER_22_8 VPWR VGND sg13g2_fill_2
XFILLER_47_641 VPWR VGND sg13g2_decap_8
XFILLER_35_836 VPWR VGND sg13g2_decap_8
X_2971_ VGND VPWR _0526_ _0525_ _0489_ sg13g2_or2_1
XFILLER_15_560 VPWR VGND sg13g2_decap_8
XFILLER_30_541 VPWR VGND sg13g2_decap_8
X_3523_ _0073_ _1039_ _1043_ net586 _1494_ VPWR VGND sg13g2_a22oi_1
X_3454_ _0977_ _0973_ _0976_ net670 _1480_ VPWR VGND sg13g2_a22oi_1
XFILLER_41_0 VPWR VGND sg13g2_fill_1
X_2405_ _1825_ _1685_ _1602_ _1646_ _1597_ VPWR VGND sg13g2_a22oi_1
X_3385_ _0911_ _0775_ _0897_ VPWR VGND sg13g2_xnor2_1
X_2336_ _1743_ _1745_ _1750_ _1755_ _1756_ VPWR VGND sg13g2_or4_1
X_2267_ VGND VPWR _1536_ net746 _1687_ net735 sg13g2_a21oi_1
X_4006_ _1437_ u_ser.state\[0\] _1415_ VPWR VGND sg13g2_nor2_2
XFILLER_26_814 VPWR VGND sg13g2_decap_8
XFILLER_38_674 VPWR VGND sg13g2_decap_8
X_2198_ net780 net785 net782 _1618_ VGND VPWR _1563_ sg13g2_nor4_2
XFILLER_13_508 VPWR VGND sg13g2_decap_8
XFILLER_25_379 VPWR VGND sg13g2_decap_8
XFILLER_21_585 VPWR VGND sg13g2_decap_8
XFILLER_5_707 VPWR VGND sg13g2_decap_8
XFILLER_1_913 VPWR VGND sg13g2_decap_8
XFILLER_0_423 VPWR VGND sg13g2_fill_2
XFILLER_49_939 VPWR VGND sg13g2_decap_8
XFILLER_48_416 VPWR VGND sg13g2_decap_8
Xhold20 u_ser.shadow_reg\[0\] VPWR VGND net69 sg13g2_dlygate4sd3_1
XFILLER_29_53 VPWR VGND sg13g2_fill_1
XFILLER_21_1012 VPWR VGND sg13g2_decap_8
XFILLER_29_685 VPWR VGND sg13g2_decap_8
XFILLER_44_666 VPWR VGND sg13g2_decap_8
XFILLER_17_858 VPWR VGND sg13g2_decap_8
XFILLER_32_839 VPWR VGND sg13g2_decap_8
XFILLER_8_523 VPWR VGND sg13g2_decap_8
XFILLER_12_574 VPWR VGND sg13g2_decap_8
XFILLER_4_795 VPWR VGND sg13g2_decap_8
XFILLER_3_294 VPWR VGND sg13g2_fill_2
XFILLER_6_1006 VPWR VGND sg13g2_decap_8
X_3170_ _0698_ net706 _0694_ VPWR VGND sg13g2_nand2_1
XFILLER_0_990 VPWR VGND sg13g2_decap_8
X_2121_ _1523_ _1525_ net765 _1541_ VPWR VGND _1540_ sg13g2_nand4_1
X_2052_ _1474_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[4\] VPWR VGND
+ sg13g2_inv_2
XFILLER_48_983 VPWR VGND sg13g2_decap_8
XFILLER_35_633 VPWR VGND sg13g2_decap_8
XFILLER_23_806 VPWR VGND sg13g2_decap_8
X_2954_ net791 sap_3_inst.alu.tmp\[6\] _0509_ VPWR VGND sg13g2_and2_1
XFILLER_31_850 VPWR VGND sg13g2_decap_8
X_2885_ VPWR VGND _0442_ net580 _0441_ net572 _0443_ net627 sg13g2_a221oi_1
X_3506_ _1027_ _1022_ _1026_ net672 _1494_ VPWR VGND sg13g2_a22oi_1
X_3437_ _0907_ _0931_ _0885_ _0961_ VPWR VGND _0954_ sg13g2_nand4_1
XFILLER_44_1023 VPWR VGND sg13g2_decap_4
X_3368_ net586 _0887_ _0892_ _0894_ _0895_ VPWR VGND sg13g2_nor4_1
X_2319_ _1739_ _1738_ VPWR VGND sg13g2_inv_2
X_3299_ _0822_ _0824_ _0816_ _0827_ VPWR VGND _0825_ sg13g2_nand4_1
XFILLER_39_950 VPWR VGND sg13g2_decap_8
XFILLER_26_611 VPWR VGND sg13g2_decap_8
XFILLER_14_828 VPWR VGND sg13g2_decap_8
XFILLER_26_688 VPWR VGND sg13g2_decap_8
XFILLER_41_658 VPWR VGND sg13g2_decap_8
XFILLER_40_157 VPWR VGND sg13g2_fill_1
XFILLER_21_382 VPWR VGND sg13g2_fill_1
XFILLER_5_504 VPWR VGND sg13g2_decap_8
Xoutput21 net32 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_710 VPWR VGND sg13g2_decap_8
Xoutput10 net10 uio_oe[1] VPWR VGND sg13g2_buf_1
XFILLER_1_787 VPWR VGND sg13g2_decap_8
Xclkbuf_5_6__f_sap_3_inst.alu.clk_regs clknet_4_3_0_sap_3_inst.alu.clk_regs clknet_5_6__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_49_736 VPWR VGND sg13g2_decap_8
XFILLER_29_482 VPWR VGND sg13g2_decap_8
XFILLER_45_942 VPWR VGND sg13g2_decap_8
XFILLER_17_655 VPWR VGND sg13g2_decap_8
XFILLER_44_463 VPWR VGND sg13g2_decap_8
XFILLER_32_636 VPWR VGND sg13g2_decap_8
XFILLER_13_872 VPWR VGND sg13g2_decap_8
XFILLER_9_854 VPWR VGND sg13g2_decap_8
X_2670_ _1959_ _0254_ _1950_ _0256_ VPWR VGND _0255_ sg13g2_nand4_1
XFILLER_4_592 VPWR VGND sg13g2_decap_8
X_3222_ net704 net698 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] _0750_
+ VPWR VGND net691 sg13g2_nand4_1
X_3153_ net730 net734 net753 _0681_ VPWR VGND sg13g2_a21o_1
X_2104_ VGND VPWR _1524_ net770 net769 sg13g2_or2_1
XFILLER_48_780 VPWR VGND sg13g2_decap_8
X_3084_ _1549_ net735 net773 _0612_ VPWR VGND sg13g2_nand3_1
XFILLER_36_920 VPWR VGND sg13g2_decap_8
XFILLER_47_290 VPWR VGND sg13g2_fill_2
X_2035_ VPWR _1457_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_35_441 VPWR VGND sg13g2_fill_1
XFILLER_23_603 VPWR VGND sg13g2_decap_8
XFILLER_36_997 VPWR VGND sg13g2_decap_8
X_3986_ _1445_ net709 _1400_ VPWR VGND sg13g2_nor2_1
X_2937_ net793 _0324_ _0493_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1000 VPWR VGND sg13g2_decap_8
X_2868_ VPWR _0426_ _0425_ VGND sg13g2_inv_1
X_2799_ _0359_ _0356_ _0358_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_518 VPWR VGND sg13g2_decap_8
Xfanout800 sap_3_inst.alu.acc\[3\] net800 VPWR VGND sg13g2_buf_8
Xclkbuf_5_13__f_sap_3_inst.alu.clk_regs clknet_4_6_0_sap_3_inst.alu.clk_regs clknet_5_13__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
Xfanout833 net835 net833 VPWR VGND sg13g2_buf_8
Xfanout822 rst_n net822 VPWR VGND sg13g2_buf_8
Xfanout811 net812 net811 VPWR VGND sg13g2_buf_8
Xfanout844 net845 net844 VPWR VGND sg13g2_buf_8
XFILLER_27_931 VPWR VGND sg13g2_decap_8
XFILLER_42_912 VPWR VGND sg13g2_decap_8
XFILLER_14_625 VPWR VGND sg13g2_decap_8
XFILLER_26_485 VPWR VGND sg13g2_decap_8
XFILLER_42_989 VPWR VGND sg13g2_decap_8
XFILLER_41_455 VPWR VGND sg13g2_decap_8
XFILLER_13_157 VPWR VGND sg13g2_fill_1
XFILLER_6_824 VPWR VGND sg13g2_decap_8
XFILLER_10_886 VPWR VGND sg13g2_decap_8
XFILLER_49_533 VPWR VGND sg13g2_decap_8
XFILLER_1_584 VPWR VGND sg13g2_decap_8
XFILLER_3_1009 VPWR VGND sg13g2_decap_8
XFILLER_18_931 VPWR VGND sg13g2_decap_8
XFILLER_36_249 VPWR VGND sg13g2_fill_1
XFILLER_33_945 VPWR VGND sg13g2_decap_8
X_3840_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\] net817 _1279_ VPWR
+ VGND sg13g2_and2_1
X_3771_ _1232_ _0908_ _0931_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_1011 VPWR VGND sg13g2_decap_8
X_2722_ net752 net750 _1634_ _0293_ VPWR VGND sg13g2_nor3_1
XFILLER_9_651 VPWR VGND sg13g2_decap_8
X_2653_ VGND VPWR _0240_ net628 net806 sg13g2_or2_1
X_2584_ _1993_ _1989_ _1986_ _1994_ VPWR VGND sg13g2_a21o_2
X_3205_ _0724_ _0727_ _0729_ _0731_ _0733_ VPWR VGND sg13g2_or4_1
XFILLER_41_1015 VPWR VGND sg13g2_decap_8
X_4185_ net821 VGND VPWR _0149_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\]
+ clknet_5_7__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_728 VPWR VGND sg13g2_decap_8
X_3136_ _0664_ net705 _0662_ VPWR VGND sg13g2_nand2_2
X_3067_ _0600_ net776 net739 VPWR VGND sg13g2_nand2_1
X_2018_ VPWR _1440_ net77 VGND sg13g2_inv_1
XFILLER_23_400 VPWR VGND sg13g2_decap_8
XFILLER_24_923 VPWR VGND sg13g2_decap_8
XFILLER_36_794 VPWR VGND sg13g2_decap_8
XFILLER_23_477 VPWR VGND sg13g2_decap_8
X_3969_ _1387_ net658 _1197_ VPWR VGND sg13g2_nand2_1
XFILLER_12_45 VPWR VGND sg13g2_fill_2
XFILLER_3_827 VPWR VGND sg13g2_decap_8
Xfanout630 _1812_ net630 VPWR VGND sg13g2_buf_8
Xfanout641 _1806_ net641 VPWR VGND sg13g2_buf_8
Xfanout685 _0867_ net685 VPWR VGND sg13g2_buf_8
Xfanout652 _0821_ net652 VPWR VGND sg13g2_buf_1
Xfanout663 _0699_ net663 VPWR VGND sg13g2_buf_8
Xfanout674 _0689_ net674 VPWR VGND sg13g2_buf_8
Xfanout696 _0657_ net696 VPWR VGND sg13g2_buf_2
XFILLER_19_717 VPWR VGND sg13g2_decap_8
XFILLER_46_569 VPWR VGND sg13g2_decap_8
XFILLER_15_945 VPWR VGND sg13g2_decap_8
XFILLER_42_786 VPWR VGND sg13g2_decap_8
XFILLER_14_499 VPWR VGND sg13g2_decap_8
XFILLER_30_926 VPWR VGND sg13g2_decap_8
XFILLER_6_621 VPWR VGND sg13g2_decap_8
XFILLER_10_683 VPWR VGND sg13g2_decap_8
XFILLER_6_698 VPWR VGND sg13g2_decap_8
XFILLER_2_882 VPWR VGND sg13g2_decap_8
XFILLER_49_330 VPWR VGND sg13g2_decap_8
XFILLER_37_569 VPWR VGND sg13g2_decap_8
XFILLER_33_742 VPWR VGND sg13g2_decap_8
X_3823_ _1267_ VPWR _1268_ VGND _1233_ _1266_ sg13g2_o21ai_1
XFILLER_20_458 VPWR VGND sg13g2_fill_1
X_3754_ VPWR VGND _1217_ net612 _1215_ net603 _1218_ _0847_ sg13g2_a221oi_1
X_3685_ _0105_ _1172_ _1173_ net624 _1498_ VPWR VGND sg13g2_a22oi_1
X_2705_ _0284_ _0285_ _0003_ VPWR VGND sg13g2_nor2_1
X_2636_ _0223_ _0224_ _0222_ _0225_ VPWR VGND sg13g2_nand3_1
XFILLER_0_808 VPWR VGND sg13g2_decap_8
X_2567_ _1805_ _1974_ _1975_ _1978_ _1979_ VPWR VGND sg13g2_and4_1
X_2498_ _1912_ net635 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\] net642
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4237_ sap_3_outputReg_serial net27 VPWR VGND sg13g2_buf_1
XFILLER_28_525 VPWR VGND sg13g2_decap_8
X_4168_ net823 VGND VPWR _0132_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3119_ _0647_ net727 _0646_ _1615_ net751 VPWR VGND sg13g2_a22oi_1
X_4099_ net818 VGND VPWR _0063_ sap_3_inst.controller.opcode\[5\] clknet_5_0__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_43_539 VPWR VGND sg13g2_decap_8
XFILLER_24_720 VPWR VGND sg13g2_decap_8
XFILLER_36_591 VPWR VGND sg13g2_decap_8
XFILLER_24_797 VPWR VGND sg13g2_decap_8
XFILLER_8_908 VPWR VGND sg13g2_decap_8
XFILLER_11_447 VPWR VGND sg13g2_fill_2
XFILLER_12_959 VPWR VGND sg13g2_decap_8
XFILLER_7_418 VPWR VGND sg13g2_fill_2
XFILLER_3_624 VPWR VGND sg13g2_decap_8
XFILLER_2_134 VPWR VGND sg13g2_fill_2
XFILLER_24_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_823 VPWR VGND sg13g2_decap_8
XFILLER_19_514 VPWR VGND sg13g2_decap_8
XFILLER_0_26 VPWR VGND sg13g2_fill_1
XFILLER_46_366 VPWR VGND sg13g2_decap_8
XFILLER_0_59 VPWR VGND sg13g2_decap_8
XFILLER_34_528 VPWR VGND sg13g2_decap_8
XFILLER_15_742 VPWR VGND sg13g2_decap_8
XFILLER_42_583 VPWR VGND sg13g2_decap_8
XFILLER_30_723 VPWR VGND sg13g2_decap_8
XFILLER_10_480 VPWR VGND sg13g2_decap_8
XFILLER_31_1025 VPWR VGND sg13g2_decap_4
XFILLER_7_985 VPWR VGND sg13g2_decap_8
XFILLER_6_495 VPWR VGND sg13g2_decap_8
X_3470_ _0993_ _0961_ _0977_ VPWR VGND sg13g2_xnor2_1
X_2421_ VGND VPWR net628 _1840_ _1841_ _1838_ sg13g2_a21oi_1
X_2352_ _1751_ _1754_ _1768_ _1771_ _1772_ VPWR VGND sg13g2_and4_1
XFILLER_9_1015 VPWR VGND sg13g2_decap_8
X_2283_ VPWR _1703_ net726 VGND sg13g2_inv_1
X_4022_ net72 u_ser.state\[1\] net813 _0188_ VPWR VGND sg13g2_a21o_1
XFILLER_38_856 VPWR VGND sg13g2_decap_8
X_3806_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] _1193_ net660 _0143_
+ VPWR VGND sg13g2_mux2_1
XFILLER_21_767 VPWR VGND sg13g2_decap_8
X_3737_ _1046_ _1047_ net594 _1209_ VPWR VGND sg13g2_nor3_1
X_3668_ net599 _0980_ _1159_ VPWR VGND sg13g2_nor2_1
X_2619_ _0206_ _0207_ _0208_ VPWR VGND sg13g2_and2_1
X_3599_ VGND VPWR _1106_ net685 net14 sg13g2_or2_1
XFILLER_0_605 VPWR VGND sg13g2_decap_8
XFILLER_29_867 VPWR VGND sg13g2_decap_8
XFILLER_44_848 VPWR VGND sg13g2_decap_8
XFILLER_16_528 VPWR VGND sg13g2_decap_8
XFILLER_12_756 VPWR VGND sg13g2_decap_8
XFILLER_24_594 VPWR VGND sg13g2_decap_8
XFILLER_34_65 VPWR VGND sg13g2_fill_1
XFILLER_8_705 VPWR VGND sg13g2_decap_8
XFILLER_4_900 VPWR VGND sg13g2_decap_8
XFILLER_4_977 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_3_498 VPWR VGND sg13g2_decap_8
XFILLER_47_620 VPWR VGND sg13g2_decap_8
XFILLER_35_815 VPWR VGND sg13g2_decap_8
XFILLER_47_697 VPWR VGND sg13g2_decap_8
XFILLER_46_163 VPWR VGND sg13g2_fill_2
X_2970_ _0525_ _0510_ _0524_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_520 VPWR VGND sg13g2_decap_8
XFILLER_30_597 VPWR VGND sg13g2_decap_8
XFILLER_7_782 VPWR VGND sg13g2_decap_8
X_3522_ VPWR VGND net602 net621 _1040_ net597 _1043_ _0862_ sg13g2_a221oi_1
X_3453_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] _0975_
+ net656 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] _0976_ net679 sg13g2_a221oi_1
X_2404_ VPWR _1824_ _1823_ VGND sg13g2_inv_1
X_3384_ _0910_ net600 _0909_ VPWR VGND sg13g2_nand2_1
X_2335_ VPWR VGND _1657_ net748 _1748_ _1594_ _1755_ net728 sg13g2_a221oi_1
X_2266_ VPWR _1686_ _1685_ VGND sg13g2_inv_1
X_4005_ _1413_ VPWR _0184_ VGND net583 _1414_ sg13g2_o21ai_1
X_2197_ _1617_ _1523_ VPWR VGND net767 sg13g2_nand2b_2
XFILLER_38_653 VPWR VGND sg13g2_decap_8
XFILLER_34_892 VPWR VGND sg13g2_decap_8
XFILLER_21_564 VPWR VGND sg13g2_decap_8
XFILLER_1_969 VPWR VGND sg13g2_decap_8
XFILLER_49_918 VPWR VGND sg13g2_decap_8
XFILLER_0_479 VPWR VGND sg13g2_decap_8
Xhold10 u_ser.shadow_reg\[1\] VPWR VGND net59 sg13g2_dlygate4sd3_1
Xhold21 u_ser.bit_pos\[1\] VPWR VGND net70 sg13g2_dlygate4sd3_1
XFILLER_29_664 VPWR VGND sg13g2_decap_8
XFILLER_17_837 VPWR VGND sg13g2_decap_8
XFILLER_44_645 VPWR VGND sg13g2_decap_8
XFILLER_16_347 VPWR VGND sg13g2_fill_1
XFILLER_32_818 VPWR VGND sg13g2_decap_8
XFILLER_8_502 VPWR VGND sg13g2_decap_8
XFILLER_12_553 VPWR VGND sg13g2_decap_8
XFILLER_24_391 VPWR VGND sg13g2_decap_8
XFILLER_40_884 VPWR VGND sg13g2_decap_8
XFILLER_8_579 VPWR VGND sg13g2_decap_8
XFILLER_4_774 VPWR VGND sg13g2_decap_8
X_2120_ net776 net781 _1540_ VPWR VGND sg13g2_nor2b_1
XFILLER_48_962 VPWR VGND sg13g2_decap_8
X_2051_ VPWR _1473_ sap_3_inst.alu.tmp\[4\] VGND sg13g2_inv_1
XFILLER_35_612 VPWR VGND sg13g2_decap_8
XFILLER_47_494 VPWR VGND sg13g2_decap_8
XFILLER_35_689 VPWR VGND sg13g2_decap_8
X_2953_ VGND VPWR _0508_ sap_3_inst.alu.tmp\[6\] net791 sg13g2_or2_1
XFILLER_16_892 VPWR VGND sg13g2_decap_8
X_2884_ VGND VPWR sap_3_inst.alu.act\[3\] net708 _0442_ net626 sg13g2_a21oi_1
X_3505_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] _1025_
+ net658 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] _1026_ net675 sg13g2_a221oi_1
XFILLER_44_1002 VPWR VGND sg13g2_decap_8
X_3436_ _0959_ VPWR _0960_ VGND net622 _0957_ sg13g2_o21ai_1
X_3367_ _0894_ _0869_ _0893_ net595 net18 VPWR VGND sg13g2_a22oi_1
X_2318_ _1737_ VPWR _1738_ VGND _1625_ _1736_ sg13g2_o21ai_1
X_3298_ _0816_ _0822_ _0824_ _0825_ _0826_ VPWR VGND sg13g2_and4_1
X_2249_ _1626_ VPWR _1669_ VGND _1652_ _1668_ sg13g2_o21ai_1
XFILLER_14_807 VPWR VGND sg13g2_decap_8
XFILLER_25_155 VPWR VGND sg13g2_fill_1
XFILLER_26_667 VPWR VGND sg13g2_decap_8
XFILLER_41_637 VPWR VGND sg13g2_decap_8
XFILLER_13_339 VPWR VGND sg13g2_fill_1
XFILLER_25_199 VPWR VGND sg13g2_fill_2
XFILLER_22_895 VPWR VGND sg13g2_decap_8
Xoutput11 net11 uio_oe[2] VPWR VGND sg13g2_buf_1
Xoutput22 net22 uio_out[5] VPWR VGND sg13g2_buf_1
Xoutput9 net9 uio_oe[0] VPWR VGND sg13g2_buf_1
XFILLER_49_715 VPWR VGND sg13g2_decap_8
XFILLER_1_766 VPWR VGND sg13g2_decap_8
XFILLER_48_269 VPWR VGND sg13g2_decap_8
XFILLER_45_921 VPWR VGND sg13g2_decap_8
XFILLER_17_634 VPWR VGND sg13g2_decap_8
XFILLER_45_998 VPWR VGND sg13g2_decap_8
XFILLER_44_442 VPWR VGND sg13g2_decap_8
XFILLER_32_615 VPWR VGND sg13g2_decap_8
XFILLER_13_851 VPWR VGND sg13g2_decap_8
XFILLER_31_158 VPWR VGND sg13g2_fill_1
XFILLER_40_681 VPWR VGND sg13g2_decap_8
XFILLER_9_833 VPWR VGND sg13g2_decap_8
XFILLER_12_350 VPWR VGND sg13g2_fill_1
XFILLER_8_343 VPWR VGND sg13g2_fill_2
XFILLER_28_1008 VPWR VGND sg13g2_decap_8
XFILLER_4_571 VPWR VGND sg13g2_decap_8
X_3221_ net701 net694 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] _0749_
+ VPWR VGND net689 sg13g2_nand4_1
X_3152_ net764 net753 _1639_ _0680_ VPWR VGND sg13g2_or3_1
X_2103_ net768 net770 _1523_ VPWR VGND sg13g2_nor2_2
X_3083_ _1645_ net733 _1605_ _0611_ VPWR VGND sg13g2_a21o_1
X_2034_ VPWR _1456_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_36_976 VPWR VGND sg13g2_decap_8
XFILLER_35_486 VPWR VGND sg13g2_decap_8
X_3985_ _1399_ VPWR _0179_ VGND net582 _1398_ sg13g2_o21ai_1
XFILLER_23_659 VPWR VGND sg13g2_decap_8
X_2936_ _0492_ _0485_ _0335_ _0484_ _0342_ VPWR VGND sg13g2_a22oi_1
X_2867_ _0425_ _0423_ _0424_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_180 VPWR VGND sg13g2_fill_2
X_2798_ _0358_ sap_3_inst.alu.tmp\[0\] net806 VPWR VGND sg13g2_nand2b_1
Xclkbuf_1_0__f_clk_div_out clknet_0_clk_div_out clknet_1_0__leaf_clk_div_out VPWR
+ VGND sg13g2_buf_8
Xfanout801 sap_3_inst.alu.acc\[2\] net801 VPWR VGND sg13g2_buf_8
Xfanout834 net835 net834 VPWR VGND sg13g2_buf_8
Xfanout823 net830 net823 VPWR VGND sg13g2_buf_8
X_3419_ _0766_ net592 _0835_ _0944_ VPWR VGND sg13g2_nor3_1
Xfanout812 _1277_ net812 VPWR VGND sg13g2_buf_8
Xfanout845 net849 net845 VPWR VGND sg13g2_buf_8
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_14_604 VPWR VGND sg13g2_decap_8
XFILLER_26_464 VPWR VGND sg13g2_decap_8
XFILLER_27_987 VPWR VGND sg13g2_decap_8
XFILLER_42_968 VPWR VGND sg13g2_decap_8
XFILLER_41_434 VPWR VGND sg13g2_decap_8
XFILLER_6_803 VPWR VGND sg13g2_decap_8
XFILLER_22_692 VPWR VGND sg13g2_decap_8
XFILLER_10_865 VPWR VGND sg13g2_decap_8
XFILLER_49_512 VPWR VGND sg13g2_decap_8
XFILLER_1_563 VPWR VGND sg13g2_decap_8
XFILLER_49_589 VPWR VGND sg13g2_decap_8
XFILLER_18_910 VPWR VGND sg13g2_decap_8
XFILLER_18_987 VPWR VGND sg13g2_decap_8
XFILLER_45_795 VPWR VGND sg13g2_decap_8
XFILLER_33_924 VPWR VGND sg13g2_decap_8
X_3770_ VPWR VGND net601 net611 _0934_ _0287_ _1231_ _0849_ sg13g2_a221oi_1
X_2721_ _1661_ _1662_ _1696_ _0292_ VPWR VGND sg13g2_nor3_1
XFILLER_9_630 VPWR VGND sg13g2_decap_8
XFILLER_12_180 VPWR VGND sg13g2_fill_1
X_2652_ VPWR VGND _0238_ _1723_ _0235_ _1468_ _0239_ net650 sg13g2_a221oi_1
X_2583_ _1993_ _1990_ _1991_ _1992_ VPWR VGND sg13g2_and3_1
X_3204_ _0724_ _0727_ _0729_ _0732_ VGND VPWR _0731_ sg13g2_nor4_2
X_4184_ net833 VGND VPWR _0148_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\]
+ clknet_5_28__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_707 VPWR VGND sg13g2_decap_8
X_3135_ _0663_ net703 net697 net692 VPWR VGND sg13g2_and3_2
X_3066_ VGND VPWR _1444_ net738 _0060_ _0599_ sg13g2_a21oi_1
X_2017_ VPWR _1439_ u_ser.bit_pos\[2\] VGND sg13g2_inv_1
XFILLER_24_902 VPWR VGND sg13g2_decap_8
XFILLER_36_773 VPWR VGND sg13g2_decap_8
XFILLER_23_456 VPWR VGND sg13g2_decap_8
XFILLER_24_979 VPWR VGND sg13g2_decap_8
X_3968_ _1386_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] net609 VPWR
+ VGND sg13g2_nand2_1
XFILLER_11_629 VPWR VGND sg13g2_decap_8
X_2919_ net581 net797 _0475_ _0037_ VPWR VGND sg13g2_a21o_1
XFILLER_12_35 VPWR VGND sg13g2_fill_2
X_3899_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] _1330_
+ _1314_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] _1331_ _1307_ sg13g2_a221oi_1
XFILLER_3_806 VPWR VGND sg13g2_decap_8
Xfanout642 _1804_ net642 VPWR VGND sg13g2_buf_8
Xfanout620 _0696_ net620 VPWR VGND sg13g2_buf_8
Xfanout631 _1812_ net631 VPWR VGND sg13g2_buf_8
Xfanout664 _0699_ net664 VPWR VGND sg13g2_buf_1
Xfanout653 _0820_ net653 VPWR VGND sg13g2_buf_8
Xfanout675 _0689_ net675 VPWR VGND sg13g2_buf_2
Xfanout697 net700 net697 VPWR VGND sg13g2_buf_8
Xfanout686 net687 net686 VPWR VGND sg13g2_buf_8
XFILLER_46_548 VPWR VGND sg13g2_decap_8
XFILLER_37_54 VPWR VGND sg13g2_fill_1
XFILLER_15_924 VPWR VGND sg13g2_decap_8
XFILLER_26_261 VPWR VGND sg13g2_fill_1
XFILLER_27_784 VPWR VGND sg13g2_decap_8
XFILLER_42_765 VPWR VGND sg13g2_decap_8
XFILLER_30_905 VPWR VGND sg13g2_decap_8
XFILLER_6_600 VPWR VGND sg13g2_decap_8
XFILLER_10_662 VPWR VGND sg13g2_decap_8
XFILLER_6_677 VPWR VGND sg13g2_decap_8
XFILLER_2_861 VPWR VGND sg13g2_decap_8
XFILLER_49_386 VPWR VGND sg13g2_decap_8
XFILLER_37_548 VPWR VGND sg13g2_decap_8
XFILLER_18_784 VPWR VGND sg13g2_decap_8
XFILLER_33_721 VPWR VGND sg13g2_decap_8
XFILLER_45_592 VPWR VGND sg13g2_decap_8
XFILLER_32_220 VPWR VGND sg13g2_fill_2
X_3822_ VPWR VGND net601 net610 _0934_ _0287_ _1267_ _0849_ sg13g2_a221oi_1
XFILLER_33_798 VPWR VGND sg13g2_decap_8
XFILLER_21_949 VPWR VGND sg13g2_decap_8
X_3753_ VGND VPWR _0843_ _1216_ _1217_ _1045_ sg13g2_a21oi_1
X_3684_ VGND VPWR net602 _1040_ _1173_ net624 sg13g2_a21oi_1
X_2704_ _0285_ net759 _1507_ VPWR VGND sg13g2_xnor2_1
X_2635_ _0224_ net646 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] net649
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2566_ _1978_ net635 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\] net644
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2497_ sap_3_inst.alu.flags\[5\] net573 _1867_ _0030_ VPWR VGND sg13g2_mux2_1
X_4236_ mem_mar_we net26 VPWR VGND sg13g2_buf_1
X_4167_ net819 VGND VPWR _0131_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_504 VPWR VGND sg13g2_decap_8
X_3118_ VGND VPWR _0646_ _1792_ _1441_ sg13g2_or2_1
X_4098_ net818 VGND VPWR _0062_ sap_3_inst.controller.opcode\[4\] clknet_5_4__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_43_518 VPWR VGND sg13g2_decap_8
X_3049_ _0593_ _1849_ _0592_ _1780_ net736 VPWR VGND sg13g2_a22oi_1
XFILLER_36_570 VPWR VGND sg13g2_decap_8
XFILLER_12_938 VPWR VGND sg13g2_decap_8
XFILLER_24_776 VPWR VGND sg13g2_decap_8
XFILLER_23_67 VPWR VGND sg13g2_fill_1
XFILLER_3_603 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_24_1000 VPWR VGND sg13g2_decap_8
XFILLER_47_802 VPWR VGND sg13g2_decap_8
XFILLER_47_879 VPWR VGND sg13g2_decap_8
XFILLER_46_345 VPWR VGND sg13g2_decap_8
XFILLER_0_38 VPWR VGND sg13g2_decap_8
XFILLER_34_507 VPWR VGND sg13g2_decap_8
XFILLER_15_721 VPWR VGND sg13g2_decap_8
XFILLER_27_581 VPWR VGND sg13g2_decap_8
XFILLER_14_220 VPWR VGND sg13g2_fill_2
XFILLER_42_562 VPWR VGND sg13g2_decap_8
XFILLER_14_242 VPWR VGND sg13g2_fill_2
XFILLER_14_253 VPWR VGND sg13g2_fill_1
XFILLER_30_702 VPWR VGND sg13g2_decap_8
XFILLER_15_798 VPWR VGND sg13g2_decap_8
XFILLER_30_779 VPWR VGND sg13g2_decap_8
XFILLER_31_1004 VPWR VGND sg13g2_decap_8
XFILLER_11_993 VPWR VGND sg13g2_decap_8
XFILLER_7_964 VPWR VGND sg13g2_decap_8
X_2420_ _1840_ sap_3_inst.alu.flags\[7\] _1839_ VPWR VGND sg13g2_nand2_1
X_2351_ net775 VPWR _1771_ VGND _1732_ _1769_ sg13g2_o21ai_1
X_2282_ _1702_ net746 net758 net754 net755 VPWR VGND sg13g2_a22oi_1
X_4021_ VPWR _0187_ _1428_ VGND sg13g2_inv_1
XFILLER_38_835 VPWR VGND sg13g2_decap_8
XFILLER_18_581 VPWR VGND sg13g2_decap_8
XFILLER_20_212 VPWR VGND sg13g2_fill_1
XFILLER_21_746 VPWR VGND sg13g2_decap_8
XFILLER_33_595 VPWR VGND sg13g2_decap_8
X_3805_ VGND VPWR _1476_ net613 _0142_ _1256_ sg13g2_a21oi_1
X_3736_ VGND VPWR net680 _1208_ _1656_ _1595_ sg13g2_a21oi_2
X_3667_ _1158_ _0984_ _1149_ net684 net22 VPWR VGND sg13g2_a22oi_1
X_2618_ _0207_ net635 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] net646
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] VPWR VGND sg13g2_a22oi_1
X_3598_ _1105_ _1076_ net22 VPWR VGND sg13g2_nand2b_1
X_2549_ _1961_ _1946_ _1960_ VPWR VGND sg13g2_nand2_2
X_4219_ net837 VGND VPWR _0182_ sap_3_inst.alu.act\[5\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_29_846 VPWR VGND sg13g2_decap_8
XFILLER_16_507 VPWR VGND sg13g2_decap_8
XFILLER_44_827 VPWR VGND sg13g2_decap_8
XFILLER_24_573 VPWR VGND sg13g2_decap_8
XFILLER_11_212 VPWR VGND sg13g2_fill_1
XFILLER_12_735 VPWR VGND sg13g2_decap_8
XFILLER_4_956 VPWR VGND sg13g2_decap_8
XFILLER_47_676 VPWR VGND sg13g2_decap_8
XFILLER_43_882 VPWR VGND sg13g2_decap_8
XFILLER_15_595 VPWR VGND sg13g2_decap_8
XFILLER_30_576 VPWR VGND sg13g2_decap_8
X_3521_ _1042_ _1041_ VPWR VGND _0846_ sg13g2_nand2b_2
XFILLER_7_761 VPWR VGND sg13g2_decap_8
XFILLER_11_790 VPWR VGND sg13g2_decap_8
X_3452_ _0975_ _0971_ _0974_ VPWR VGND sg13g2_nand2_1
X_2403_ _1550_ net734 _1823_ VPWR VGND sg13g2_nor2_2
X_3383_ _0907_ _0889_ _0909_ VPWR VGND sg13g2_xor2_1
X_2334_ _1754_ _1638_ _1753_ VPWR VGND sg13g2_nand2_1
X_2265_ _1508_ _1558_ _1685_ VPWR VGND sg13g2_nor2_2
XFILLER_38_632 VPWR VGND sg13g2_decap_8
X_4004_ VGND VPWR _0552_ _1389_ _1414_ _1412_ sg13g2_a21oi_1
X_2196_ net766 _1524_ _1616_ VPWR VGND sg13g2_nor2_1
XFILLER_37_131 VPWR VGND sg13g2_fill_1
XFILLER_26_849 VPWR VGND sg13g2_decap_8
XFILLER_41_819 VPWR VGND sg13g2_decap_8
XFILLER_34_871 VPWR VGND sg13g2_decap_8
XFILLER_21_543 VPWR VGND sg13g2_decap_8
XFILLER_14_1010 VPWR VGND sg13g2_decap_8
X_3719_ net616 _1046_ _1083_ _1199_ VPWR VGND sg13g2_nor3_1
XFILLER_1_948 VPWR VGND sg13g2_decap_8
Xhold11 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[2\] VPWR VGND net60
+ sg13g2_dlygate4sd3_1
Xhold22 regFile_serial VPWR VGND net71 sg13g2_dlygate4sd3_1
X_4039__4 VPWR net40 clknet_leaf_0_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_29_643 VPWR VGND sg13g2_decap_8
XFILLER_44_624 VPWR VGND sg13g2_decap_8
XFILLER_17_816 VPWR VGND sg13g2_decap_8
XFILLER_40_863 VPWR VGND sg13g2_decap_8
XFILLER_12_532 VPWR VGND sg13g2_decap_8
XFILLER_8_558 VPWR VGND sg13g2_decap_8
XFILLER_4_753 VPWR VGND sg13g2_decap_8
XFILLER_48_941 VPWR VGND sg13g2_decap_8
X_2050_ VPWR _1472_ sap_3_inst.alu.tmp\[3\] VGND sg13g2_inv_1
XFILLER_47_473 VPWR VGND sg13g2_decap_8
Xclkbuf_5_21__f_sap_3_inst.alu.clk_regs clknet_4_10_0_sap_3_inst.alu.clk_regs clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_16_871 VPWR VGND sg13g2_decap_8
XFILLER_35_668 VPWR VGND sg13g2_decap_8
XFILLER_37_1010 VPWR VGND sg13g2_decap_8
X_2952_ net33 _0311_ _0507_ VPWR VGND sg13g2_nor2b_1
X_2883_ _0441_ _0440_ _0439_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_885 VPWR VGND sg13g2_decap_8
X_3504_ _1023_ _1024_ _1021_ _1025_ VPWR VGND sg13g2_nand3_1
X_3435_ VGND VPWR net622 _0958_ _0959_ net598 sg13g2_a21oi_1
X_3366_ _0893_ net597 net10 VPWR VGND sg13g2_nand2b_1
X_2317_ _1737_ net743 _1565_ _1505_ net758 VPWR VGND sg13g2_a22oi_1
X_3297_ net743 _1711_ net776 _0825_ VPWR VGND sg13g2_nand3_1
Xheichips25_template_35 VPWR VGND uo_out[6] sg13g2_tielo
X_2248_ _1641_ _1665_ _1637_ _1668_ VPWR VGND _1667_ sg13g2_nand4_1
XFILLER_39_985 VPWR VGND sg13g2_decap_8
X_2179_ _1527_ _1564_ _1580_ _1599_ VPWR VGND sg13g2_nor3_2
XFILLER_26_646 VPWR VGND sg13g2_decap_8
XFILLER_41_616 VPWR VGND sg13g2_decap_8
XFILLER_22_874 VPWR VGND sg13g2_decap_8
XFILLER_5_539 VPWR VGND sg13g2_decap_8
Xoutput23 net33 uio_out[6] VPWR VGND sg13g2_buf_1
Xoutput12 net12 uio_oe[3] VPWR VGND sg13g2_buf_1
XFILLER_1_745 VPWR VGND sg13g2_decap_8
XFILLER_0_288 VPWR VGND sg13g2_fill_2
XFILLER_45_900 VPWR VGND sg13g2_decap_8
XFILLER_17_613 VPWR VGND sg13g2_decap_8
XFILLER_44_421 VPWR VGND sg13g2_decap_8
XFILLER_45_977 VPWR VGND sg13g2_decap_8
XFILLER_44_498 VPWR VGND sg13g2_decap_8
XFILLER_13_830 VPWR VGND sg13g2_decap_8
XFILLER_40_660 VPWR VGND sg13g2_decap_8
XFILLER_9_812 VPWR VGND sg13g2_decap_8
XFILLER_9_889 VPWR VGND sg13g2_decap_8
XFILLER_4_550 VPWR VGND sg13g2_decap_8
X_3220_ _1479_ _0690_ _0748_ VPWR VGND sg13g2_nor2_1
X_3151_ _0679_ net752 net726 VPWR VGND sg13g2_nand2b_1
X_2102_ net766 net756 _1522_ VPWR VGND sg13g2_nor2_1
X_3082_ VGND VPWR net731 _1657_ _0610_ _1596_ sg13g2_a21oi_1
X_2033_ VPWR _1455_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_36_955 VPWR VGND sg13g2_decap_8
XFILLER_23_638 VPWR VGND sg13g2_decap_8
X_3984_ _1399_ sap_3_inst.alu.act\[2\] net582 VPWR VGND sg13g2_nand2_1
X_2935_ sap_3_inst.alu.tmp\[5\] _0344_ net794 _0491_ VPWR VGND sg13g2_nand3_1
X_2866_ VGND VPWR _0384_ _0398_ _0424_ _0382_ sg13g2_a21oi_1
XFILLER_31_682 VPWR VGND sg13g2_decap_8
X_2797_ _0357_ net804 sap_3_inst.alu.tmp\[1\] VPWR VGND sg13g2_xnor2_1
Xfanout824 net827 net824 VPWR VGND sg13g2_buf_8
Xfanout813 _0185_ net813 VPWR VGND sg13g2_buf_8
Xfanout802 sap_3_inst.alu.acc\[2\] net802 VPWR VGND sg13g2_buf_2
X_3418_ VGND VPWR _0943_ _0942_ _0802_ sg13g2_or2_1
Xfanout835 net849 net835 VPWR VGND sg13g2_buf_8
X_3349_ _0876_ net677 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] net679
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] VPWR VGND sg13g2_a22oi_1
Xfanout846 net847 net846 VPWR VGND sg13g2_buf_8
XFILLER_39_782 VPWR VGND sg13g2_decap_8
XFILLER_26_443 VPWR VGND sg13g2_decap_8
XFILLER_27_966 VPWR VGND sg13g2_decap_8
XFILLER_42_947 VPWR VGND sg13g2_decap_8
XFILLER_13_115 VPWR VGND sg13g2_fill_2
XFILLER_22_671 VPWR VGND sg13g2_decap_8
XFILLER_10_844 VPWR VGND sg13g2_decap_8
XFILLER_21_170 VPWR VGND sg13g2_fill_2
XFILLER_6_859 VPWR VGND sg13g2_decap_8
XFILLER_1_542 VPWR VGND sg13g2_decap_8
XFILLER_49_568 VPWR VGND sg13g2_decap_8
XFILLER_29_270 VPWR VGND sg13g2_fill_1
XFILLER_18_966 VPWR VGND sg13g2_decap_8
XFILLER_33_903 VPWR VGND sg13g2_decap_8
XFILLER_45_774 VPWR VGND sg13g2_decap_8
XFILLER_17_487 VPWR VGND sg13g2_decap_8
XFILLER_41_980 VPWR VGND sg13g2_decap_8
XFILLER_20_619 VPWR VGND sg13g2_decap_8
X_2720_ _1573_ VPWR _0291_ VGND _1609_ _1648_ sg13g2_o21ai_1
XFILLER_9_686 VPWR VGND sg13g2_decap_8
X_2651_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] _0237_
+ net640 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] _0238_ net645 sg13g2_a221oi_1
X_2582_ _1992_ net642 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] net646
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] VPWR VGND sg13g2_a22oi_1
X_3203_ _0731_ _0728_ _0730_ VPWR VGND sg13g2_nand2_1
X_4183_ net823 VGND VPWR _0147_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3134_ net702 net691 _0662_ VPWR VGND sg13g2_nor2_2
X_3065_ net738 net19 _0599_ VPWR VGND sg13g2_nor2_1
X_2016_ VPWR _1438_ u_ser.state\[0\] VGND sg13g2_inv_1
XFILLER_36_752 VPWR VGND sg13g2_decap_8
Xclkbuf_5_18__f_sap_3_inst.alu.clk_regs clknet_4_9_0_sap_3_inst.alu.clk_regs clknet_5_18__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_23_435 VPWR VGND sg13g2_decap_8
XFILLER_24_958 VPWR VGND sg13g2_decap_8
X_3967_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] _1212_ net656 _0175_
+ VPWR VGND sg13g2_mux2_1
XFILLER_11_608 VPWR VGND sg13g2_decap_8
X_2918_ net581 _0444_ _0474_ _0475_ VPWR VGND sg13g2_nor3_1
X_3898_ _1327_ _1328_ _1325_ _1330_ VPWR VGND _1329_ sg13g2_nand4_1
X_2849_ _0399_ net574 _0408_ VPWR VGND sg13g2_nor2b_1
XFILLER_5_8 VPWR VGND sg13g2_fill_1
Xfanout632 net633 net632 VPWR VGND sg13g2_buf_8
Xfanout621 _0693_ net621 VPWR VGND sg13g2_buf_8
Xfanout610 _0705_ net610 VPWR VGND sg13g2_buf_8
Xfanout654 _0820_ net654 VPWR VGND sg13g2_buf_1
Xfanout676 net677 net676 VPWR VGND sg13g2_buf_8
Xfanout665 _0697_ net665 VPWR VGND sg13g2_buf_8
Xfanout643 _1804_ net643 VPWR VGND sg13g2_buf_8
Xfanout687 _0688_ net687 VPWR VGND sg13g2_buf_8
Xfanout698 net699 net698 VPWR VGND sg13g2_buf_2
XFILLER_46_527 VPWR VGND sg13g2_decap_8
XFILLER_2_1022 VPWR VGND sg13g2_decap_8
XFILLER_15_903 VPWR VGND sg13g2_decap_8
XFILLER_27_763 VPWR VGND sg13g2_decap_8
XFILLER_42_744 VPWR VGND sg13g2_decap_8
XFILLER_18_1008 VPWR VGND sg13g2_decap_8
XFILLER_10_641 VPWR VGND sg13g2_decap_8
XFILLER_6_656 VPWR VGND sg13g2_decap_8
XFILLER_2_840 VPWR VGND sg13g2_decap_8
XFILLER_49_365 VPWR VGND sg13g2_decap_8
XFILLER_37_527 VPWR VGND sg13g2_decap_8
XFILLER_18_763 VPWR VGND sg13g2_decap_8
XFILLER_45_571 VPWR VGND sg13g2_decap_8
XFILLER_33_700 VPWR VGND sg13g2_decap_8
XFILLER_21_928 VPWR VGND sg13g2_decap_8
X_3821_ _1184_ net608 net713 _1266_ VPWR VGND sg13g2_a21o_1
XFILLER_33_777 VPWR VGND sg13g2_decap_8
X_3752_ VGND VPWR _0711_ _0842_ _1216_ _0873_ sg13g2_a21oi_1
X_2703_ _1536_ _0284_ _0002_ VPWR VGND sg13g2_nor2_1
XFILLER_9_483 VPWR VGND sg13g2_decap_8
X_3683_ _1170_ VPWR _1172_ VGND _1030_ _1171_ sg13g2_o21ai_1
X_2634_ _0223_ net636 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] net639
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2565_ _1977_ net630 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] net636
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2496_ net573 _1911_ VPWR VGND _1900_ sg13g2_nand2b_2
X_4235_ mem_ram_we net25 VPWR VGND sg13g2_buf_1
X_4166_ net843 VGND VPWR _0130_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\]
+ clknet_5_27__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3117_ _0640_ net757 _0643_ _0645_ VPWR VGND sg13g2_a21o_1
X_4097_ net818 VGND VPWR _0061_ sap_3_inst.controller.opcode\[3\] clknet_5_4__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3048_ net736 _1553_ _1732_ _0592_ VPWR VGND sg13g2_nor3_1
XFILLER_24_755 VPWR VGND sg13g2_decap_8
XFILLER_12_917 VPWR VGND sg13g2_decap_8
XFILLER_20_983 VPWR VGND sg13g2_decap_8
XFILLER_3_659 VPWR VGND sg13g2_decap_8
XFILLER_2_136 VPWR VGND sg13g2_fill_1
XFILLER_47_858 VPWR VGND sg13g2_decap_8
XFILLER_19_549 VPWR VGND sg13g2_decap_8
XFILLER_15_700 VPWR VGND sg13g2_decap_8
XFILLER_27_560 VPWR VGND sg13g2_decap_8
XFILLER_42_541 VPWR VGND sg13g2_decap_8
XFILLER_15_777 VPWR VGND sg13g2_decap_8
XFILLER_30_758 VPWR VGND sg13g2_decap_8
XFILLER_7_943 VPWR VGND sg13g2_decap_8
XFILLER_11_972 VPWR VGND sg13g2_decap_8
Xsap_3_inst.clock.clock_gate_inst sap_3_inst.clock.hlt clknet_1_0__leaf_clk_div_out
+ sap_3_inst.alu.clk VPWR VGND sg13g2_lgcp_1
X_2350_ _1602_ VPWR _1770_ VGND net745 net728 sg13g2_o21ai_1
X_2281_ VPWR VGND _1553_ _1660_ _1676_ _1566_ _1701_ _1571_ sg13g2_a221oi_1
X_4020_ _1427_ VPWR _1428_ VGND net78 _0186_ sg13g2_o21ai_1
XFILLER_38_814 VPWR VGND sg13g2_decap_8
XFILLER_18_560 VPWR VGND sg13g2_decap_8
XFILLER_25_519 VPWR VGND sg13g2_decap_8
XFILLER_46_891 VPWR VGND sg13g2_decap_8
XFILLER_21_725 VPWR VGND sg13g2_decap_8
XFILLER_33_574 VPWR VGND sg13g2_decap_8
X_3804_ net613 _1189_ _1255_ _1256_ VPWR VGND sg13g2_nor3_1
X_3735_ _0121_ _1069_ _1207_ net617 _1497_ VPWR VGND sg13g2_a22oi_1
X_3666_ _1157_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] net623 VPWR
+ VGND sg13g2_nand2_1
XFILLER_47_1012 VPWR VGND sg13g2_decap_8
X_2617_ _0206_ net641 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] net644
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] VPWR VGND sg13g2_a22oi_1
X_3597_ _1098_ _1104_ _0086_ VPWR VGND sg13g2_nor2b_1
X_2548_ _1960_ _1950_ _1959_ VPWR VGND sg13g2_nand2_2
X_2479_ _1895_ _1893_ _1894_ VPWR VGND sg13g2_nand2_1
X_4218_ net837 VGND VPWR _0181_ sap_3_inst.alu.act\[4\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_29_825 VPWR VGND sg13g2_decap_8
X_4149_ net828 VGND VPWR _0113_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\]
+ clknet_5_15__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_44_806 VPWR VGND sg13g2_decap_8
XFILLER_18_68 VPWR VGND sg13g2_fill_2
XFILLER_37_891 VPWR VGND sg13g2_decap_8
XFILLER_24_552 VPWR VGND sg13g2_decap_8
XFILLER_12_714 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_3_0__leaf_clk clkload0/X VPWR VGND sg13g2_buf_1
XFILLER_20_780 VPWR VGND sg13g2_decap_8
XFILLER_4_935 VPWR VGND sg13g2_decap_8
XFILLER_47_655 VPWR VGND sg13g2_decap_8
XFILLER_43_861 VPWR VGND sg13g2_decap_8
XFILLER_15_574 VPWR VGND sg13g2_decap_8
XFILLER_30_555 VPWR VGND sg13g2_decap_8
X_3520_ _0721_ VPWR _1041_ VGND net592 _0840_ sg13g2_o21ai_1
XFILLER_7_740 VPWR VGND sg13g2_decap_8
X_3451_ _0974_ net665 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] net677
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] VPWR VGND sg13g2_a22oi_1
X_2402_ _1822_ _1520_ net728 VPWR VGND sg13g2_nand2_1
X_3382_ _0711_ _0842_ _0884_ _0908_ VGND VPWR _0907_ sg13g2_nor4_2
X_2333_ net753 _1614_ _1587_ _1753_ VPWR VGND sg13g2_nand3_1
X_2264_ net744 _1681_ _1682_ _1683_ _1684_ VPWR VGND sg13g2_nor4_1
XFILLER_38_611 VPWR VGND sg13g2_decap_8
X_4003_ _1413_ sap_3_inst.alu.act\[7\] net583 VPWR VGND sg13g2_nand2_1
X_2195_ _1586_ _1599_ _1608_ _1615_ VGND VPWR _1613_ sg13g2_nor4_2
XFILLER_26_828 VPWR VGND sg13g2_decap_8
XFILLER_38_688 VPWR VGND sg13g2_decap_8
XFILLER_25_349 VPWR VGND sg13g2_fill_2
XFILLER_34_850 VPWR VGND sg13g2_decap_8
XFILLER_21_522 VPWR VGND sg13g2_decap_8
XFILLER_21_599 VPWR VGND sg13g2_decap_8
X_3718_ _1195_ VPWR _0113_ VGND _1196_ _1198_ sg13g2_o21ai_1
X_3649_ _1087_ _1143_ _1144_ VPWR VGND sg13g2_nor2_1
XFILLER_1_927 VPWR VGND sg13g2_decap_8
Xhold23 sap_3_outputReg_start_sync VPWR VGND net72 sg13g2_dlygate4sd3_1
Xhold12 u_ser.state\[0\] VPWR VGND net61 sg13g2_dlygate4sd3_1
XFILLER_29_622 VPWR VGND sg13g2_decap_8
XFILLER_21_1026 VPWR VGND sg13g2_fill_2
XFILLER_44_603 VPWR VGND sg13g2_decap_8
XFILLER_43_113 VPWR VGND sg13g2_fill_1
XFILLER_29_699 VPWR VGND sg13g2_decap_8
XFILLER_12_511 VPWR VGND sg13g2_decap_8
XFILLER_25_883 VPWR VGND sg13g2_decap_8
XFILLER_40_842 VPWR VGND sg13g2_decap_8
XFILLER_8_537 VPWR VGND sg13g2_decap_8
XFILLER_12_588 VPWR VGND sg13g2_decap_8
XFILLER_4_732 VPWR VGND sg13g2_decap_8
XFILLER_48_920 VPWR VGND sg13g2_decap_8
XFILLER_48_997 VPWR VGND sg13g2_decap_8
XFILLER_47_452 VPWR VGND sg13g2_decap_8
XFILLER_35_647 VPWR VGND sg13g2_decap_8
XFILLER_16_850 VPWR VGND sg13g2_decap_8
X_2951_ net581 net794 _0506_ _0038_ VPWR VGND sg13g2_a21o_1
XFILLER_31_864 VPWR VGND sg13g2_decap_8
X_2882_ VGND VPWR net574 _0425_ _0440_ net707 sg13g2_a21oi_1
XFILLER_30_374 VPWR VGND sg13g2_fill_2
X_3503_ _1024_ net678 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] net681
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3434_ _0844_ VPWR _0958_ VGND _0756_ _0944_ sg13g2_o21ai_1
X_3365_ net599 _0891_ _0892_ VPWR VGND sg13g2_nor2_1
X_3296_ _0823_ VPWR _0824_ VGND net750 _0622_ sg13g2_o21ai_1
X_2316_ _1624_ _1726_ _1733_ _1735_ _1736_ VPWR VGND sg13g2_and4_1
Xheichips25_template_36 VPWR VGND uo_out[7] sg13g2_tielo
X_2247_ _1653_ _1661_ _1664_ _1666_ _1667_ VPWR VGND sg13g2_nor4_1
XFILLER_39_964 VPWR VGND sg13g2_decap_8
X_2178_ net765 _1590_ _1511_ _1598_ VPWR VGND sg13g2_nand3_1
XFILLER_26_625 VPWR VGND sg13g2_decap_8
XFILLER_38_485 VPWR VGND sg13g2_decap_8
XFILLER_22_853 VPWR VGND sg13g2_decap_8
XFILLER_21_341 VPWR VGND sg13g2_fill_1
XFILLER_5_518 VPWR VGND sg13g2_decap_8
X_4041__6 VPWR net42 clknet_leaf_2_sap_3_inst.alu.clk VGND sg13g2_inv_1
Xoutput24 net34 uio_out[7] VPWR VGND sg13g2_buf_1
Xoutput13 net13 uio_oe[4] VPWR VGND sg13g2_buf_1
XFILLER_1_724 VPWR VGND sg13g2_decap_8
XFILLER_45_956 VPWR VGND sg13g2_decap_8
XFILLER_44_400 VPWR VGND sg13g2_decap_8
XFILLER_29_496 VPWR VGND sg13g2_decap_8
XFILLER_17_669 VPWR VGND sg13g2_decap_8
XFILLER_44_477 VPWR VGND sg13g2_decap_8
XFILLER_25_680 VPWR VGND sg13g2_decap_8
XFILLER_31_127 VPWR VGND sg13g2_fill_2
XFILLER_31_149 VPWR VGND sg13g2_fill_1
XFILLER_13_886 VPWR VGND sg13g2_decap_8
XFILLER_9_868 VPWR VGND sg13g2_decap_8
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
X_3150_ VGND VPWR _1587_ _0676_ _0678_ net726 sg13g2_a21oi_1
X_3081_ net752 VPWR _0609_ VGND _1576_ _1656_ sg13g2_o21ai_1
X_2101_ _1514_ _1518_ _1441_ _1521_ VPWR VGND sg13g2_nand3_1
X_2032_ VPWR _1454_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_48_794 VPWR VGND sg13g2_decap_8
XFILLER_36_934 VPWR VGND sg13g2_decap_8
XFILLER_23_617 VPWR VGND sg13g2_decap_8
X_3983_ VGND VPWR _0388_ net710 _1398_ _1397_ sg13g2_a21oi_1
X_2934_ _0490_ _0459_ _0487_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_661 VPWR VGND sg13g2_decap_8
X_2865_ _0423_ net799 sap_3_inst.alu.tmp\[3\] VPWR VGND sg13g2_xnor2_1
XFILLER_11_1014 VPWR VGND sg13g2_decap_8
X_2796_ sap_3_inst.alu.tmp\[1\] net804 _0356_ VPWR VGND sg13g2_xor2_1
Xfanout825 net827 net825 VPWR VGND sg13g2_buf_8
Xfanout814 net79 net814 VPWR VGND sg13g2_buf_8
Xfanout803 sap_3_inst.alu.acc\[1\] net803 VPWR VGND sg13g2_buf_8
X_3417_ VGND VPWR net591 _0800_ _0942_ _0766_ sg13g2_a21oi_1
Xfanout836 net837 net836 VPWR VGND sg13g2_buf_8
X_3348_ _0875_ net660 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] net668
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] VPWR VGND sg13g2_a22oi_1
Xfanout847 net848 net847 VPWR VGND sg13g2_buf_2
XFILLER_46_709 VPWR VGND sg13g2_decap_8
XFILLER_45_208 VPWR VGND sg13g2_fill_1
X_3279_ _0807_ _0711_ _0806_ VPWR VGND sg13g2_nand2_1
XFILLER_39_761 VPWR VGND sg13g2_decap_8
XFILLER_26_422 VPWR VGND sg13g2_decap_8
XFILLER_27_945 VPWR VGND sg13g2_decap_8
XFILLER_38_293 VPWR VGND sg13g2_fill_1
XFILLER_42_926 VPWR VGND sg13g2_decap_8
XFILLER_41_414 VPWR VGND sg13g2_decap_8
XFILLER_14_639 VPWR VGND sg13g2_decap_8
XFILLER_26_499 VPWR VGND sg13g2_decap_8
XFILLER_41_469 VPWR VGND sg13g2_decap_8
XFILLER_22_650 VPWR VGND sg13g2_decap_8
XFILLER_10_823 VPWR VGND sg13g2_decap_8
XFILLER_6_838 VPWR VGND sg13g2_decap_8
XFILLER_1_521 VPWR VGND sg13g2_decap_8
XFILLER_49_547 VPWR VGND sg13g2_decap_8
XFILLER_1_598 VPWR VGND sg13g2_decap_8
XFILLER_37_709 VPWR VGND sg13g2_decap_8
XFILLER_18_945 VPWR VGND sg13g2_decap_8
XFILLER_45_753 VPWR VGND sg13g2_decap_8
XFILLER_33_959 VPWR VGND sg13g2_decap_8
XFILLER_8_120 VPWR VGND sg13g2_fill_2
XFILLER_13_683 VPWR VGND sg13g2_decap_8
XFILLER_34_1025 VPWR VGND sg13g2_decap_4
X_2650_ _0232_ _0236_ net648 _0237_ VPWR VGND sg13g2_nand3_1
XFILLER_9_665 VPWR VGND sg13g2_decap_8
XFILLER_8_164 VPWR VGND sg13g2_fill_1
X_2581_ _1991_ net636 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] net641
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_882 VPWR VGND sg13g2_decap_8
X_3202_ _0730_ net677 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] net679
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] VPWR VGND sg13g2_a22oi_1
X_4182_ net843 VGND VPWR _0146_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\]
+ clknet_5_26__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3133_ _0661_ net704 net690 VPWR VGND sg13g2_nand2_1
X_3064_ _0598_ VPWR _0059_ VGND net739 _0227_ sg13g2_o21ai_1
XFILLER_48_591 VPWR VGND sg13g2_decap_8
X_2015_ VPWR _1437_ u_ser.state\[1\] VGND sg13g2_inv_1
XFILLER_36_731 VPWR VGND sg13g2_decap_8
XFILLER_23_414 VPWR VGND sg13g2_decap_8
XFILLER_24_937 VPWR VGND sg13g2_decap_8
X_3966_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] _1131_ net655 _0174_
+ VPWR VGND sg13g2_mux2_1
X_2917_ VPWR VGND _0473_ net627 _0472_ sap_3_inst.alu.act\[4\] _0474_ net707 sg13g2_a221oi_1
X_3897_ _1329_ net809 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] _1309_
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2848_ net574 _0402_ _0406_ _0407_ VPWR VGND sg13g2_nor3_1
X_2779_ _1955_ _0199_ _0340_ VPWR VGND sg13g2_nor2_2
Xfanout611 net615 net611 VPWR VGND sg13g2_buf_8
Xfanout600 net601 net600 VPWR VGND sg13g2_buf_8
Xfanout633 _1811_ net633 VPWR VGND sg13g2_buf_8
Xfanout622 _0693_ net622 VPWR VGND sg13g2_buf_1
Xfanout655 net659 net655 VPWR VGND sg13g2_buf_8
Xfanout644 _1803_ net644 VPWR VGND sg13g2_buf_8
Xfanout666 _0697_ net666 VPWR VGND sg13g2_buf_8
XFILLER_46_506 VPWR VGND sg13g2_decap_8
Xfanout688 _0687_ net688 VPWR VGND sg13g2_buf_8
Xfanout677 _0665_ net677 VPWR VGND sg13g2_buf_8
Xfanout699 net700 net699 VPWR VGND sg13g2_buf_1
XFILLER_2_1001 VPWR VGND sg13g2_decap_8
XFILLER_27_742 VPWR VGND sg13g2_decap_8
XFILLER_42_723 VPWR VGND sg13g2_decap_8
XFILLER_15_959 VPWR VGND sg13g2_decap_8
XFILLER_41_255 VPWR VGND sg13g2_fill_2
XFILLER_10_620 VPWR VGND sg13g2_decap_8
XFILLER_23_981 VPWR VGND sg13g2_decap_8
XFILLER_6_635 VPWR VGND sg13g2_decap_8
XFILLER_10_697 VPWR VGND sg13g2_decap_8
XFILLER_5_167 VPWR VGND sg13g2_fill_1
XFILLER_2_896 VPWR VGND sg13g2_decap_8
XFILLER_49_344 VPWR VGND sg13g2_decap_8
XFILLER_37_506 VPWR VGND sg13g2_decap_8
XFILLER_18_742 VPWR VGND sg13g2_decap_8
XFILLER_45_550 VPWR VGND sg13g2_decap_8
XFILLER_33_756 VPWR VGND sg13g2_decap_8
XFILLER_21_907 VPWR VGND sg13g2_decap_8
X_3820_ _0148_ _1147_ _1265_ net608 _1454_ VPWR VGND sg13g2_a22oi_1
X_3751_ net713 VPWR _1215_ VGND net9 net652 sg13g2_o21ai_1
X_2702_ sap_3_inst.controller.stage\[0\] _0284_ _0001_ VPWR VGND sg13g2_nor2_1
X_3682_ net607 VPWR _1171_ VGND net679 _1032_ sg13g2_o21ai_1
X_2633_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] net642
+ net641 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] _0222_ net723 sg13g2_a221oi_1
X_2564_ _1976_ net639 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] net641
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2495_ VPWR VGND net576 _1903_ _1910_ net6 _1911_ _1858_ sg13g2_a221oi_1
X_4165_ net828 VGND VPWR _0129_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\]
+ clknet_5_14__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3116_ VGND VPWR _0643_ _0644_ _0640_ net757 sg13g2_a21oi_2
XFILLER_28_539 VPWR VGND sg13g2_decap_8
X_4096_ net818 VGND VPWR _0060_ sap_3_inst.controller.opcode\[2\] clknet_5_4__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3047_ _0591_ VPWR _0049_ VGND _0588_ _0590_ sg13g2_o21ai_1
XFILLER_24_734 VPWR VGND sg13g2_decap_8
XFILLER_20_962 VPWR VGND sg13g2_decap_8
X_3949_ _1375_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] _1300_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_3_638 VPWR VGND sg13g2_decap_8
XFILLER_48_22 VPWR VGND sg13g2_decap_4
XFILLER_47_837 VPWR VGND sg13g2_decap_8
XFILLER_19_528 VPWR VGND sg13g2_decap_8
XFILLER_42_520 VPWR VGND sg13g2_decap_8
XFILLER_14_222 VPWR VGND sg13g2_fill_1
XFILLER_9_27 VPWR VGND sg13g2_decap_4
XFILLER_15_756 VPWR VGND sg13g2_decap_8
XFILLER_42_597 VPWR VGND sg13g2_decap_8
XFILLER_14_288 VPWR VGND sg13g2_fill_2
XFILLER_30_737 VPWR VGND sg13g2_decap_8
XFILLER_11_951 VPWR VGND sg13g2_decap_8
XFILLER_7_922 VPWR VGND sg13g2_decap_8
XFILLER_10_494 VPWR VGND sg13g2_decap_8
XFILLER_13_91 VPWR VGND sg13g2_fill_1
XFILLER_7_999 VPWR VGND sg13g2_decap_8
X_2280_ _1700_ _1566_ _1571_ VPWR VGND sg13g2_nand2_1
XFILLER_2_693 VPWR VGND sg13g2_decap_8
XFILLER_46_870 VPWR VGND sg13g2_decap_8
XFILLER_21_704 VPWR VGND sg13g2_decap_8
XFILLER_33_553 VPWR VGND sg13g2_decap_8
X_3803_ net654 net713 _0837_ _1254_ _1255_ VPWR VGND sg13g2_nor4_1
X_3734_ VGND VPWR net603 _1040_ _1207_ net616 sg13g2_a21oi_1
Xclkbuf_4_15_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_15_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3665_ _0102_ _1154_ _1156_ net624 _1479_ VPWR VGND sg13g2_a22oi_1
X_2616_ _0205_ net762 _0204_ VPWR VGND sg13g2_nand2_1
X_3596_ _1099_ _1100_ net667 _1104_ VPWR VGND _1103_ sg13g2_nand4_1
X_2547_ _1959_ _1958_ VPWR VGND _1951_ sg13g2_nand2b_2
XFILLER_0_619 VPWR VGND sg13g2_decap_8
X_2478_ _1894_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] net722
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4217_ net832 VGND VPWR _0180_ sap_3_inst.alu.act\[3\] clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_29_804 VPWR VGND sg13g2_decap_8
X_4148_ net826 VGND VPWR _0112_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\]
+ clknet_5_3__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4079_ net836 VGND VPWR _0043_ sap_3_inst.out\[2\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_37_870 VPWR VGND sg13g2_decap_8
XFILLER_24_531 VPWR VGND sg13g2_decap_8
XFILLER_8_719 VPWR VGND sg13g2_decap_8
Xclkload1 VPWR clkload1/Y clknet_3_1__leaf_clk VGND sg13g2_inv_1
XFILLER_4_914 VPWR VGND sg13g2_decap_8
XFILLER_47_634 VPWR VGND sg13g2_decap_8
XFILLER_19_336 VPWR VGND sg13g2_fill_2
XFILLER_35_829 VPWR VGND sg13g2_decap_8
XFILLER_43_840 VPWR VGND sg13g2_decap_8
XFILLER_15_553 VPWR VGND sg13g2_decap_8
XFILLER_42_394 VPWR VGND sg13g2_decap_8
XFILLER_30_534 VPWR VGND sg13g2_decap_8
XFILLER_7_796 VPWR VGND sg13g2_decap_8
X_3450_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] _0972_
+ net664 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] _0973_ net668 sg13g2_a221oi_1
X_2401_ net756 _1678_ _1821_ VPWR VGND sg13g2_nor2_1
X_3381_ _0906_ VPWR _0907_ VGND sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[2\]
+ net622 sg13g2_o21ai_1
X_2332_ _1692_ net725 _1752_ VPWR VGND sg13g2_nor2_1
XFILLER_2_490 VPWR VGND sg13g2_decap_8
X_4002_ net710 net788 _1412_ VPWR VGND sg13g2_nor2b_1
X_2263_ VGND VPWR net732 _1654_ _1683_ net751 sg13g2_a21oi_1
Xclkbuf_4_7_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_7_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2194_ _1511_ _1562_ _1444_ _1614_ VPWR VGND sg13g2_nand3_1
XFILLER_26_807 VPWR VGND sg13g2_decap_8
XFILLER_38_667 VPWR VGND sg13g2_decap_8
XFILLER_19_892 VPWR VGND sg13g2_decap_8
XFILLER_21_501 VPWR VGND sg13g2_decap_8
XFILLER_21_578 VPWR VGND sg13g2_decap_8
X_3717_ _1198_ _1197_ net578 VPWR VGND sg13g2_nand2b_1
X_3648_ net597 VPWR _1143_ VGND net10 _1138_ sg13g2_o21ai_1
XFILLER_1_906 VPWR VGND sg13g2_decap_8
X_3579_ _1086_ _1089_ _1090_ VPWR VGND sg13g2_nor2_1
XFILLER_48_409 VPWR VGND sg13g2_decap_8
Xhold13 _0195_ VPWR VGND net62 sg13g2_dlygate4sd3_1
Xhold24 _0188_ VPWR VGND net73 sg13g2_dlygate4sd3_1
XFILLER_29_601 VPWR VGND sg13g2_decap_8
XFILLER_21_1005 VPWR VGND sg13g2_decap_8
XFILLER_29_678 VPWR VGND sg13g2_decap_8
XFILLER_44_659 VPWR VGND sg13g2_decap_8
XFILLER_25_862 VPWR VGND sg13g2_decap_8
XFILLER_40_821 VPWR VGND sg13g2_decap_8
XFILLER_40_898 VPWR VGND sg13g2_decap_8
XFILLER_8_516 VPWR VGND sg13g2_decap_8
XFILLER_12_567 VPWR VGND sg13g2_decap_8
XFILLER_4_711 VPWR VGND sg13g2_decap_8
XFILLER_4_788 VPWR VGND sg13g2_decap_8
XFILLER_0_983 VPWR VGND sg13g2_decap_8
XFILLER_47_431 VPWR VGND sg13g2_decap_8
XFILLER_48_976 VPWR VGND sg13g2_decap_8
XFILLER_35_626 VPWR VGND sg13g2_decap_8
X_2950_ net581 _0476_ _0505_ _0506_ VPWR VGND sg13g2_nor3_1
X_2881_ net574 _0417_ _0438_ _0439_ VPWR VGND sg13g2_nor3_1
XFILLER_31_843 VPWR VGND sg13g2_decap_8
XFILLER_7_593 VPWR VGND sg13g2_decap_8
X_3502_ _1023_ net662 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] _0695_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3433_ _0957_ _0933_ _0953_ VPWR VGND sg13g2_xnor2_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_44_1016 VPWR VGND sg13g2_decap_8
X_3364_ _0889_ _0890_ _0891_ VPWR VGND sg13g2_nor2_1
XFILLER_32_0 VPWR VGND sg13g2_fill_1
X_2315_ _1728_ _1731_ _1734_ _1735_ VPWR VGND sg13g2_nor3_1
X_3295_ _0823_ net750 _1654_ VPWR VGND sg13g2_nand2_1
X_2246_ VGND VPWR _1573_ _1651_ _1666_ net749 sg13g2_a21oi_1
XFILLER_39_943 VPWR VGND sg13g2_decap_8
XFILLER_26_604 VPWR VGND sg13g2_decap_8
X_2177_ _1512_ net764 _1591_ _1597_ VPWR VGND sg13g2_nor3_2
XFILLER_22_832 VPWR VGND sg13g2_decap_8
Xoutput25 net25 uo_out[0] VPWR VGND sg13g2_buf_1
Xoutput14 net14 uio_oe[5] VPWR VGND sg13g2_buf_1
XFILLER_1_703 VPWR VGND sg13g2_decap_8
XFILLER_49_729 VPWR VGND sg13g2_decap_8
XFILLER_48_206 VPWR VGND sg13g2_fill_1
XFILLER_48_239 VPWR VGND sg13g2_fill_2
XFILLER_45_935 VPWR VGND sg13g2_decap_8
XFILLER_44_456 VPWR VGND sg13g2_decap_8
XFILLER_17_648 VPWR VGND sg13g2_decap_8
XFILLER_32_629 VPWR VGND sg13g2_decap_8
XFILLER_13_865 VPWR VGND sg13g2_decap_8
XFILLER_40_695 VPWR VGND sg13g2_decap_8
XFILLER_9_847 VPWR VGND sg13g2_decap_8
Xclkbuf_5_26__f_sap_3_inst.alu.clk_regs clknet_4_13_0_sap_3_inst.alu.clk_regs clknet_5_26__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_4_585 VPWR VGND sg13g2_decap_8
X_3080_ _0607_ VPWR _0608_ VGND _1588_ _1748_ sg13g2_o21ai_1
XFILLER_0_780 VPWR VGND sg13g2_decap_8
X_2100_ net778 _1515_ net763 _1520_ VPWR VGND sg13g2_nor3_2
XFILLER_39_239 VPWR VGND sg13g2_fill_2
XFILLER_48_773 VPWR VGND sg13g2_decap_8
X_2031_ VPWR _1453_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_36_913 VPWR VGND sg13g2_decap_8
X_3982_ net709 net801 _1397_ VPWR VGND sg13g2_nor2b_1
X_2933_ _0489_ _0459_ _0487_ VPWR VGND sg13g2_nand2_1
XFILLER_22_139 VPWR VGND sg13g2_fill_1
XFILLER_31_640 VPWR VGND sg13g2_decap_8
X_2864_ sap_3_inst.alu.tmp\[3\] net799 _0422_ VPWR VGND sg13g2_xor2_1
X_2795_ _0355_ net803 sap_3_inst.alu.tmp\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_30_194 VPWR VGND sg13g2_fill_1
XFILLER_8_880 VPWR VGND sg13g2_decap_8
Xfanout804 sap_3_inst.alu.acc\[1\] net804 VPWR VGND sg13g2_buf_1
X_3416_ net586 _0938_ _0940_ _0941_ VPWR VGND sg13g2_nor3_1
Xfanout815 sap_3_inst.reg_file.array_serializer_inst.word_index\[3\] net815 VPWR VGND
+ sg13g2_buf_8
Xfanout826 net827 net826 VPWR VGND sg13g2_buf_8
Xfanout848 net849 net848 VPWR VGND sg13g2_buf_1
Xfanout837 net840 net837 VPWR VGND sg13g2_buf_8
X_3347_ _0066_ _0871_ _0830_ net587 _1468_ VPWR VGND sg13g2_a22oi_1
X_3278_ _0722_ _0805_ _0806_ VPWR VGND sg13g2_nor2_1
XFILLER_39_740 VPWR VGND sg13g2_decap_8
X_2229_ _1649_ net732 _1648_ VPWR VGND sg13g2_nand2_1
XFILLER_26_401 VPWR VGND sg13g2_decap_8
XFILLER_27_924 VPWR VGND sg13g2_decap_8
XFILLER_42_905 VPWR VGND sg13g2_decap_8
XFILLER_14_618 VPWR VGND sg13g2_decap_8
XFILLER_26_478 VPWR VGND sg13g2_decap_8
XFILLER_41_448 VPWR VGND sg13g2_decap_8
XFILLER_13_117 VPWR VGND sg13g2_fill_1
XFILLER_35_990 VPWR VGND sg13g2_decap_8
XFILLER_10_802 VPWR VGND sg13g2_decap_8
XFILLER_21_172 VPWR VGND sg13g2_fill_1
XFILLER_6_817 VPWR VGND sg13g2_decap_8
XFILLER_10_879 VPWR VGND sg13g2_decap_8
XFILLER_1_500 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_1_577 VPWR VGND sg13g2_decap_8
XFILLER_27_1022 VPWR VGND sg13g2_decap_8
XFILLER_49_526 VPWR VGND sg13g2_decap_8
XFILLER_18_924 VPWR VGND sg13g2_decap_8
XFILLER_45_732 VPWR VGND sg13g2_decap_8
XFILLER_44_231 VPWR VGND sg13g2_fill_2
XFILLER_17_445 VPWR VGND sg13g2_fill_1
XFILLER_33_938 VPWR VGND sg13g2_decap_8
XFILLER_13_662 VPWR VGND sg13g2_decap_8
XFILLER_34_1004 VPWR VGND sg13g2_decap_8
XFILLER_9_644 VPWR VGND sg13g2_decap_8
XFILLER_40_492 VPWR VGND sg13g2_decap_8
X_2580_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] net649
+ net644 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] _1990_ net723 sg13g2_a221oi_1
XFILLER_5_861 VPWR VGND sg13g2_decap_8
X_4181_ net829 VGND VPWR _0145_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\]
+ clknet_5_26__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3201_ _0726_ VPWR _0729_ VGND _1486_ net612 sg13g2_o21ai_1
XFILLER_41_1008 VPWR VGND sg13g2_decap_8
X_3132_ net706 net690 _0660_ VPWR VGND sg13g2_and2_1
XFILLER_48_570 VPWR VGND sg13g2_decap_8
X_3063_ _0598_ net782 net739 VPWR VGND sg13g2_nand2_1
XFILLER_36_710 VPWR VGND sg13g2_decap_8
XFILLER_24_916 VPWR VGND sg13g2_decap_8
XFILLER_36_787 VPWR VGND sg13g2_decap_8
X_3965_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] _1189_ net657 _0173_
+ VPWR VGND sg13g2_mux2_1
X_2916_ VGND VPWR net575 _0458_ _0473_ net707 sg13g2_a21oi_1
X_3896_ _1328_ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] _1306_
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_32_993 VPWR VGND sg13g2_decap_8
X_2847_ _0403_ _0404_ _0392_ _0406_ VPWR VGND _0405_ sg13g2_nand4_1
X_2778_ _1957_ net683 net762 _0339_ VPWR VGND sg13g2_nand3_1
Xfanout612 net615 net612 VPWR VGND sg13g2_buf_1
Xfanout601 net604 net601 VPWR VGND sg13g2_buf_8
Xfanout623 net624 net623 VPWR VGND sg13g2_buf_8
Xfanout656 net659 net656 VPWR VGND sg13g2_buf_8
Xfanout645 _1803_ net645 VPWR VGND sg13g2_buf_8
Xfanout634 net635 net634 VPWR VGND sg13g2_buf_8
Xfanout667 net668 net667 VPWR VGND sg13g2_buf_8
Xfanout678 _0663_ net678 VPWR VGND sg13g2_buf_8
Xfanout689 _0687_ net689 VPWR VGND sg13g2_buf_8
XFILLER_27_721 VPWR VGND sg13g2_decap_8
XFILLER_42_702 VPWR VGND sg13g2_decap_8
XFILLER_15_938 VPWR VGND sg13g2_decap_8
XFILLER_27_798 VPWR VGND sg13g2_decap_8
XFILLER_42_779 VPWR VGND sg13g2_decap_8
XFILLER_23_960 VPWR VGND sg13g2_decap_8
XFILLER_30_919 VPWR VGND sg13g2_decap_8
XFILLER_6_614 VPWR VGND sg13g2_decap_8
XFILLER_10_676 VPWR VGND sg13g2_decap_8
XFILLER_2_875 VPWR VGND sg13g2_decap_8
XFILLER_49_323 VPWR VGND sg13g2_decap_8
XFILLER_18_721 VPWR VGND sg13g2_decap_8
XFILLER_17_275 VPWR VGND sg13g2_fill_2
XFILLER_18_798 VPWR VGND sg13g2_decap_8
XFILLER_33_735 VPWR VGND sg13g2_decap_8
X_3750_ _0129_ _1214_ _1069_ net594 _1496_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_982 VPWR VGND sg13g2_decap_8
X_2701_ _1764_ _0283_ _0284_ VPWR VGND sg13g2_nor2_2
X_3681_ net652 _1169_ _1170_ VPWR VGND sg13g2_nor2_1
X_2632_ _0221_ _0219_ _0220_ VPWR VGND sg13g2_nand2_1
X_2563_ _1975_ net633 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] net723
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2494_ _1905_ _1909_ _1904_ _1910_ VPWR VGND sg13g2_nand3_1
XFILLER_4_83 VPWR VGND sg13g2_fill_1
X_4164_ net826 VGND VPWR _0128_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\]
+ clknet_5_13__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4095_ net818 VGND VPWR _0059_ sap_3_inst.controller.opcode\[1\] clknet_5_5__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3115_ _0642_ _1516_ _0641_ _0643_ VPWR VGND sg13g2_a21o_1
XFILLER_28_518 VPWR VGND sg13g2_decap_8
XFILLER_49_890 VPWR VGND sg13g2_decap_8
X_3046_ _0591_ sap_3_inst.alu.carry _0589_ VPWR VGND sg13g2_nand2b_1
XFILLER_24_713 VPWR VGND sg13g2_decap_8
XFILLER_36_584 VPWR VGND sg13g2_decap_8
XFILLER_23_37 VPWR VGND sg13g2_fill_1
XFILLER_20_941 VPWR VGND sg13g2_decap_8
XFILLER_32_790 VPWR VGND sg13g2_decap_8
X_3948_ _1374_ _1314_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] net809
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3879_ VGND VPWR net815 net816 _1312_ _1311_ sg13g2_a21oi_1
XFILLER_3_617 VPWR VGND sg13g2_decap_8
XFILLER_2_149 VPWR VGND sg13g2_fill_1
XFILLER_24_1014 VPWR VGND sg13g2_decap_8
XFILLER_47_816 VPWR VGND sg13g2_decap_8
XFILLER_19_507 VPWR VGND sg13g2_decap_8
XFILLER_46_359 VPWR VGND sg13g2_decap_8
XFILLER_14_201 VPWR VGND sg13g2_fill_2
XFILLER_15_735 VPWR VGND sg13g2_decap_8
XFILLER_27_595 VPWR VGND sg13g2_decap_8
XFILLER_42_576 VPWR VGND sg13g2_decap_8
XFILLER_30_716 VPWR VGND sg13g2_decap_8
XFILLER_7_901 VPWR VGND sg13g2_decap_8
XFILLER_11_930 VPWR VGND sg13g2_decap_8
XFILLER_31_1018 VPWR VGND sg13g2_decap_8
XFILLER_7_978 VPWR VGND sg13g2_decap_8
XFILLER_9_1008 VPWR VGND sg13g2_decap_8
XFILLER_2_672 VPWR VGND sg13g2_decap_8
XFILLER_38_849 VPWR VGND sg13g2_decap_8
XFILLER_18_595 VPWR VGND sg13g2_decap_8
XFILLER_33_532 VPWR VGND sg13g2_decap_8
X_3802_ _0756_ _0836_ _1254_ VPWR VGND sg13g2_nor2_1
X_3733_ _0120_ _1110_ _1206_ net617 _1489_ VPWR VGND sg13g2_a22oi_1
X_3664_ VGND VPWR _1102_ _1155_ _1156_ net624 sg13g2_a21oi_1
X_2615_ _0204_ _1946_ _0203_ VPWR VGND sg13g2_nand2_1
X_3595_ _1103_ _1102_ _1101_ VPWR VGND sg13g2_nand2b_1
X_2546_ _1958_ _1956_ _1957_ VPWR VGND sg13g2_nand2_2
X_2477_ _1893_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] net647
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4216_ net832 VGND VPWR _0179_ sap_3_inst.alu.act\[2\] clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
Xclkbuf_5_0__f_sap_3_inst.alu.clk_regs clknet_4_0_0_sap_3_inst.alu.clk_regs clknet_5_0__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_4147_ net824 VGND VPWR _0111_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\]
+ clknet_5_11__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4078_ net831 VGND VPWR _0042_ sap_3_inst.out\[1\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3029_ _0574_ _0202_ _0333_ VPWR VGND sg13g2_nand2_1
XFILLER_24_510 VPWR VGND sg13g2_decap_8
XFILLER_24_587 VPWR VGND sg13g2_decap_8
XFILLER_12_749 VPWR VGND sg13g2_decap_8
Xclkload2 clknet_3_2__leaf_clk clkload2/X VPWR VGND sg13g2_buf_1
XFILLER_47_613 VPWR VGND sg13g2_decap_8
XFILLER_35_808 VPWR VGND sg13g2_decap_8
XFILLER_28_882 VPWR VGND sg13g2_decap_8
XFILLER_15_532 VPWR VGND sg13g2_decap_8
XFILLER_43_896 VPWR VGND sg13g2_decap_8
XFILLER_30_513 VPWR VGND sg13g2_decap_8
XFILLER_7_775 VPWR VGND sg13g2_decap_8
X_2400_ _1723_ _1819_ _1820_ VPWR VGND sg13g2_nor2b_1
X_3380_ _0901_ _0905_ net622 _0906_ VPWR VGND sg13g2_nand3_1
X_2331_ VPWR VGND net752 _1659_ _1655_ _1611_ _1751_ _1644_ sg13g2_a221oi_1
XFILLER_3_981 VPWR VGND sg13g2_decap_8
X_2262_ VGND VPWR _1603_ net748 _1682_ net727 sg13g2_a21oi_1
X_4001_ _1411_ VPWR _0183_ VGND net583 _1410_ sg13g2_o21ai_1
X_2193_ net780 _1512_ _1563_ _1613_ VPWR VGND sg13g2_nor3_2
XFILLER_38_646 VPWR VGND sg13g2_decap_8
XFILLER_19_871 VPWR VGND sg13g2_decap_8
XFILLER_34_885 VPWR VGND sg13g2_decap_8
XFILLER_14_1024 VPWR VGND sg13g2_decap_4
XFILLER_21_557 VPWR VGND sg13g2_decap_8
X_3716_ _1197_ net603 _1042_ VPWR VGND sg13g2_nand2_1
X_3647_ _1135_ VPWR _0098_ VGND _1136_ _1142_ sg13g2_o21ai_1
X_3578_ net668 VPWR _1089_ VGND _1087_ _1088_ sg13g2_o21ai_1
X_2529_ _1940_ VPWR _1941_ VGND _1550_ net727 sg13g2_o21ai_1
Xhold14 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[3\] VPWR VGND net63
+ sg13g2_dlygate4sd3_1
Xhold25 sap_3_inst.reg_file.array_serializer_inst.word_index\[0\] VPWR VGND net74
+ sg13g2_dlygate4sd3_1
XFILLER_21_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_657 VPWR VGND sg13g2_decap_8
XFILLER_44_638 VPWR VGND sg13g2_decap_8
XFILLER_16_329 VPWR VGND sg13g2_fill_1
XFILLER_25_841 VPWR VGND sg13g2_decap_8
XFILLER_40_800 VPWR VGND sg13g2_decap_8
XFILLER_12_546 VPWR VGND sg13g2_decap_8
XFILLER_24_384 VPWR VGND sg13g2_decap_8
XFILLER_40_877 VPWR VGND sg13g2_decap_8
XFILLER_4_767 VPWR VGND sg13g2_decap_8
XFILLER_3_266 VPWR VGND sg13g2_fill_1
XFILLER_0_962 VPWR VGND sg13g2_decap_8
XFILLER_48_955 VPWR VGND sg13g2_decap_8
XFILLER_47_410 VPWR VGND sg13g2_decap_8
XFILLER_35_605 VPWR VGND sg13g2_decap_8
XFILLER_47_487 VPWR VGND sg13g2_decap_8
XFILLER_16_885 VPWR VGND sg13g2_decap_8
XFILLER_37_1024 VPWR VGND sg13g2_decap_4
XFILLER_43_693 VPWR VGND sg13g2_decap_8
X_2880_ _0431_ _0437_ _0429_ _0438_ VPWR VGND sg13g2_nand3_1
XFILLER_31_822 VPWR VGND sg13g2_decap_8
XFILLER_30_376 VPWR VGND sg13g2_fill_1
XFILLER_31_899 VPWR VGND sg13g2_decap_8
XFILLER_7_572 VPWR VGND sg13g2_decap_8
X_3501_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] net672
+ net666 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] _1022_ net677 sg13g2_a221oi_1
X_3432_ _0908_ _0930_ net590 _0956_ VPWR VGND _0953_ sg13g2_nand4_1
X_3363_ VGND VPWR _0710_ _0846_ _0890_ _0883_ sg13g2_a21oi_1
X_3294_ _1654_ net742 _0809_ _0822_ VPWR VGND sg13g2_a21o_1
X_2314_ _1732_ net765 _1660_ _1734_ VPWR VGND sg13g2_a21o_1
X_2245_ _1658_ _1663_ _1665_ VPWR VGND sg13g2_nor2_1
XFILLER_39_922 VPWR VGND sg13g2_decap_8
X_2176_ _1590_ _1593_ _1511_ _1596_ VPWR VGND sg13g2_nand3_1
XFILLER_39_999 VPWR VGND sg13g2_decap_8
XFILLER_22_811 VPWR VGND sg13g2_decap_8
XFILLER_34_682 VPWR VGND sg13g2_decap_8
XFILLER_22_888 VPWR VGND sg13g2_decap_8
Xoutput15 net15 uio_oe[6] VPWR VGND sg13g2_buf_1
Xoutput26 net26 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_759 VPWR VGND sg13g2_decap_8
XFILLER_49_708 VPWR VGND sg13g2_decap_8
XFILLER_5_1022 VPWR VGND sg13g2_decap_8
XFILLER_45_914 VPWR VGND sg13g2_decap_8
XFILLER_17_627 VPWR VGND sg13g2_decap_8
XFILLER_44_435 VPWR VGND sg13g2_decap_8
XFILLER_32_608 VPWR VGND sg13g2_decap_8
XFILLER_12_321 VPWR VGND sg13g2_fill_2
XFILLER_13_844 VPWR VGND sg13g2_decap_8
XFILLER_9_826 VPWR VGND sg13g2_decap_8
XFILLER_40_674 VPWR VGND sg13g2_decap_8
XFILLER_4_564 VPWR VGND sg13g2_decap_8
XFILLER_48_752 VPWR VGND sg13g2_decap_8
X_2030_ VPWR _1452_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_36_969 VPWR VGND sg13g2_decap_8
X_3981_ _1396_ VPWR _0178_ VGND net582 _1395_ sg13g2_o21ai_1
X_2932_ VPWR _0488_ _0487_ VGND sg13g2_inv_1
XFILLER_16_682 VPWR VGND sg13g2_decap_8
XFILLER_43_490 VPWR VGND sg13g2_decap_8
X_2863_ net798 sap_3_inst.alu.tmp\[3\] _0421_ VPWR VGND sg13g2_nor2_1
XFILLER_31_696 VPWR VGND sg13g2_decap_8
X_2794_ VGND VPWR _1459_ net580 _0033_ _0354_ sg13g2_a21oi_1
XFILLER_7_61 VPWR VGND sg13g2_fill_2
Xfanout805 net806 net805 VPWR VGND sg13g2_buf_8
X_3415_ VGND VPWR net572 net595 _0940_ _0939_ sg13g2_a21oi_1
Xfanout816 sap_3_inst.reg_file.array_serializer_inst.word_index\[2\] net816 VPWR VGND
+ sg13g2_buf_8
Xfanout827 net830 net827 VPWR VGND sg13g2_buf_8
Xfanout849 rst_n net849 VPWR VGND sg13g2_buf_8
Xfanout838 net840 net838 VPWR VGND sg13g2_buf_8
X_3346_ net598 VPWR _0874_ VGND net592 net654 sg13g2_o21ai_1
XFILLER_27_903 VPWR VGND sg13g2_decap_8
X_3277_ _0741_ _0755_ _0732_ _0805_ VPWR VGND _0802_ sg13g2_nand4_1
X_2228_ _1648_ _1642_ net755 net746 _1534_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_796 VPWR VGND sg13g2_decap_8
X_2159_ VGND VPWR _1569_ _1574_ _1579_ _1578_ sg13g2_a21oi_1
XFILLER_26_48 VPWR VGND sg13g2_fill_1
XFILLER_26_457 VPWR VGND sg13g2_decap_8
XFILLER_41_427 VPWR VGND sg13g2_decap_8
XFILLER_42_36 VPWR VGND sg13g2_fill_1
XFILLER_22_685 VPWR VGND sg13g2_decap_8
XFILLER_10_858 VPWR VGND sg13g2_decap_8
XFILLER_27_1001 VPWR VGND sg13g2_decap_8
XFILLER_49_505 VPWR VGND sg13g2_decap_8
XFILLER_1_556 VPWR VGND sg13g2_decap_8
XFILLER_18_903 VPWR VGND sg13g2_decap_8
XFILLER_45_711 VPWR VGND sg13g2_decap_8
XFILLER_45_788 VPWR VGND sg13g2_decap_8
XFILLER_33_917 VPWR VGND sg13g2_decap_8
XFILLER_32_438 VPWR VGND sg13g2_fill_2
XFILLER_13_641 VPWR VGND sg13g2_decap_8
XFILLER_41_994 VPWR VGND sg13g2_decap_8
XFILLER_9_623 VPWR VGND sg13g2_decap_8
XFILLER_40_471 VPWR VGND sg13g2_decap_8
XFILLER_8_122 VPWR VGND sg13g2_fill_1
XFILLER_5_840 VPWR VGND sg13g2_decap_8
X_4180_ net826 VGND VPWR _0144_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3200_ _0728_ net655 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] net664
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] VPWR VGND sg13g2_a22oi_1
X_3131_ VPWR VGND _0656_ _0643_ _0654_ net757 _0659_ _0640_ sg13g2_a221oi_1
X_3062_ net31 net785 net738 _0058_ VPWR VGND sg13g2_mux2_1
XFILLER_36_766 VPWR VGND sg13g2_decap_8
XFILLER_17_991 VPWR VGND sg13g2_decap_8
XFILLER_35_298 VPWR VGND sg13g2_decap_4
X_3964_ _1385_ VPWR _0172_ VGND net608 _1186_ sg13g2_o21ai_1
XFILLER_23_449 VPWR VGND sg13g2_decap_8
X_2915_ _0471_ VPWR _0472_ VGND _0448_ _0449_ sg13g2_o21ai_1
X_3895_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] _1308_
+ _1327_ net807 sg13g2_a21oi_1
XFILLER_32_972 VPWR VGND sg13g2_decap_8
X_2846_ _0405_ _0401_ _0329_ _0383_ _0342_ VPWR VGND sg13g2_a22oi_1
XFILLER_31_493 VPWR VGND sg13g2_decap_8
X_2777_ _1956_ _0199_ _0338_ VPWR VGND sg13g2_nor2_1
Xfanout613 net615 net613 VPWR VGND sg13g2_buf_8
Xfanout602 net603 net602 VPWR VGND sg13g2_buf_8
Xfanout624 _0664_ net624 VPWR VGND sg13g2_buf_8
Xfanout657 net659 net657 VPWR VGND sg13g2_buf_8
Xfanout646 _1802_ net646 VPWR VGND sg13g2_buf_8
Xfanout635 _1809_ net635 VPWR VGND sg13g2_buf_8
X_3329_ _1847_ _0852_ _0853_ _0857_ VPWR VGND sg13g2_nor3_1
Xfanout679 _0663_ net679 VPWR VGND sg13g2_buf_8
Xfanout668 _0695_ net668 VPWR VGND sg13g2_buf_8
XFILLER_27_700 VPWR VGND sg13g2_decap_8
XFILLER_37_36 VPWR VGND sg13g2_fill_1
XFILLER_39_593 VPWR VGND sg13g2_decap_8
XFILLER_15_917 VPWR VGND sg13g2_decap_8
XFILLER_27_777 VPWR VGND sg13g2_decap_8
XFILLER_42_758 VPWR VGND sg13g2_decap_8
XFILLER_22_482 VPWR VGND sg13g2_decap_8
XFILLER_10_655 VPWR VGND sg13g2_decap_8
XFILLER_5_125 VPWR VGND sg13g2_fill_1
XFILLER_2_854 VPWR VGND sg13g2_decap_8
XFILLER_49_302 VPWR VGND sg13g2_decap_8
XFILLER_49_379 VPWR VGND sg13g2_decap_8
XFILLER_18_700 VPWR VGND sg13g2_decap_8
XFILLER_18_777 VPWR VGND sg13g2_decap_8
XFILLER_45_585 VPWR VGND sg13g2_decap_8
XFILLER_33_714 VPWR VGND sg13g2_decap_8
XFILLER_14_961 VPWR VGND sg13g2_decap_8
XFILLER_41_791 VPWR VGND sg13g2_decap_8
X_2700_ VPWR VGND _0279_ _1531_ _0282_ net728 _0283_ _0280_ sg13g2_a221oi_1
X_3680_ VGND VPWR net34 _1138_ _1169_ _1168_ sg13g2_a21oi_1
XFILLER_9_497 VPWR VGND sg13g2_decap_8
X_2631_ _0220_ net630 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] net644
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2562_ _1974_ net646 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] net649
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2493_ _1909_ _1906_ _1907_ _1908_ VPWR VGND sg13g2_and3_1
X_4232_ net835 VGND VPWR net62 u_ser.bit_pos\[2\] clknet_3_1__leaf_clk sg13g2_dfrbpq_1
X_4163_ net826 VGND VPWR _0127_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\]
+ clknet_5_9__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4094_ net818 VGND VPWR _0058_ sap_3_inst.controller.opcode\[0\] clknet_5_4__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3114_ net729 _1716_ sap_3_inst.controller.opcode\[4\] _0642_ VPWR VGND sg13g2_nand3_1
X_3045_ _0589_ VPWR _0590_ VGND _0574_ _0575_ sg13g2_o21ai_1
XFILLER_36_563 VPWR VGND sg13g2_decap_8
XFILLER_24_769 VPWR VGND sg13g2_decap_8
X_3947_ net811 net53 _1373_ _0167_ VPWR VGND sg13g2_a21o_1
XFILLER_20_920 VPWR VGND sg13g2_decap_8
X_3878_ sap_3_inst.reg_file.array_serializer_inst.word_index\[1\] sap_3_inst.reg_file.array_serializer_inst.word_index\[0\]
+ net815 net816 _1311_ VPWR VGND sg13g2_nor4_1
X_2829_ _0386_ _0384_ _0388_ VPWR VGND sg13g2_xor2_1
XFILLER_20_997 VPWR VGND sg13g2_decap_8
XFILLER_15_714 VPWR VGND sg13g2_decap_8
XFILLER_27_574 VPWR VGND sg13g2_decap_8
XFILLER_42_555 VPWR VGND sg13g2_decap_8
XFILLER_11_986 VPWR VGND sg13g2_decap_8
XFILLER_7_957 VPWR VGND sg13g2_decap_8
XFILLER_2_651 VPWR VGND sg13g2_decap_8
XFILLER_38_828 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_18_574 VPWR VGND sg13g2_decap_8
X_4046__11 VPWR net47 clknet_leaf_1_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_33_511 VPWR VGND sg13g2_decap_8
XFILLER_45_382 VPWR VGND sg13g2_decap_8
X_3801_ VGND VPWR net662 _1186_ _0141_ _1253_ sg13g2_a21oi_1
XFILLER_33_588 VPWR VGND sg13g2_decap_8
XFILLER_21_739 VPWR VGND sg13g2_decap_8
X_3732_ net665 _1064_ _1206_ VPWR VGND sg13g2_and2_1
X_2082__2 VPWR net38 clknet_leaf_0_sap_3_inst.alu.clk VGND sg13g2_inv_1
X_3663_ _1155_ _1149_ net13 VPWR VGND sg13g2_nand2b_1
X_2614_ _0199_ _0201_ _1959_ _0203_ VPWR VGND _0202_ sg13g2_nand4_1
X_3594_ _1102_ net685 net21 VPWR VGND sg13g2_nand2b_1
XFILLER_47_1026 VPWR VGND sg13g2_fill_2
X_2545_ _1442_ _1948_ _1957_ VPWR VGND sg13g2_nor2_2
X_2476_ _1892_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] net645
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4215_ net832 VGND VPWR _0178_ sap_3_inst.alu.act\[1\] clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_4146_ net841 VGND VPWR _0110_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\]
+ clknet_5_31__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_839 VPWR VGND sg13g2_decap_8
X_4077_ net831 VGND VPWR _0041_ sap_3_inst.out\[0\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3028_ net788 sap_3_inst.out\[7\] net718 _0048_ VPWR VGND sg13g2_mux2_1
XFILLER_12_728 VPWR VGND sg13g2_decap_8
XFILLER_24_566 VPWR VGND sg13g2_decap_8
XFILLER_11_238 VPWR VGND sg13g2_fill_2
Xclkload3 VPWR clkload3/Y clknet_3_3__leaf_clk VGND sg13g2_inv_1
XFILLER_20_794 VPWR VGND sg13g2_decap_8
XFILLER_4_949 VPWR VGND sg13g2_decap_8
XFILLER_8_1020 VPWR VGND sg13g2_decap_8
XFILLER_47_669 VPWR VGND sg13g2_decap_8
XFILLER_28_861 VPWR VGND sg13g2_decap_8
XFILLER_15_511 VPWR VGND sg13g2_decap_8
XFILLER_43_875 VPWR VGND sg13g2_decap_8
XFILLER_15_588 VPWR VGND sg13g2_decap_8
XFILLER_42_385 VPWR VGND sg13g2_decap_4
XFILLER_42_374 VPWR VGND sg13g2_fill_1
XFILLER_30_569 VPWR VGND sg13g2_decap_8
XFILLER_11_783 VPWR VGND sg13g2_decap_8
XFILLER_7_754 VPWR VGND sg13g2_decap_8
XFILLER_3_960 VPWR VGND sg13g2_decap_8
X_2330_ net730 _1749_ _1750_ VPWR VGND sg13g2_nor2_1
X_2261_ VGND VPWR _1582_ _1598_ _1681_ _1634_ sg13g2_a21oi_1
X_4000_ _1411_ sap_3_inst.alu.act\[6\] net583 VPWR VGND sg13g2_nand2_1
X_2192_ net780 net786 _1563_ _1612_ VPWR VGND sg13g2_nor3_1
XFILLER_38_625 VPWR VGND sg13g2_decap_8
XFILLER_19_850 VPWR VGND sg13g2_decap_8
XFILLER_34_864 VPWR VGND sg13g2_decap_8
XFILLER_21_536 VPWR VGND sg13g2_decap_8
XFILLER_14_1003 VPWR VGND sg13g2_decap_8
X_3715_ net603 _1071_ _1196_ VPWR VGND sg13g2_nor2_1
X_3646_ VGND VPWR _1140_ _1141_ _1142_ _0874_ sg13g2_a21oi_1
X_3577_ net605 VPWR _1088_ VGND net10 _1076_ sg13g2_o21ai_1
X_2528_ net724 _1939_ _1940_ VPWR VGND sg13g2_nor2_1
Xhold15 u_ser.shadow_reg\[2\] VPWR VGND net64 sg13g2_dlygate4sd3_1
Xhold26 sap_3_inst.reg_file.array_serializer_inst.state\[1\] VPWR VGND net75 sg13g2_dlygate4sd3_1
X_2459_ _1877_ _1876_ _1723_ VPWR VGND sg13g2_nand2b_1
XFILLER_29_636 VPWR VGND sg13g2_decap_8
XFILLER_17_809 VPWR VGND sg13g2_decap_8
X_4129_ net829 VGND VPWR _0093_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\]
+ clknet_5_3__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_44_617 VPWR VGND sg13g2_decap_8
XFILLER_16_308 VPWR VGND sg13g2_fill_2
XFILLER_25_820 VPWR VGND sg13g2_decap_8
XFILLER_36_190 VPWR VGND sg13g2_fill_1
XFILLER_12_525 VPWR VGND sg13g2_decap_8
XFILLER_25_897 VPWR VGND sg13g2_decap_8
XFILLER_40_856 VPWR VGND sg13g2_decap_8
XFILLER_20_591 VPWR VGND sg13g2_decap_8
XFILLER_4_746 VPWR VGND sg13g2_decap_8
XFILLER_0_941 VPWR VGND sg13g2_decap_8
XFILLER_48_934 VPWR VGND sg13g2_decap_8
XFILLER_47_466 VPWR VGND sg13g2_decap_8
XFILLER_34_138 VPWR VGND sg13g2_fill_2
XFILLER_43_672 VPWR VGND sg13g2_decap_8
XFILLER_16_864 VPWR VGND sg13g2_decap_8
XFILLER_31_801 VPWR VGND sg13g2_decap_8
XFILLER_37_1003 VPWR VGND sg13g2_decap_8
XFILLER_15_385 VPWR VGND sg13g2_fill_2
XFILLER_31_878 VPWR VGND sg13g2_decap_8
X_3500_ _1021_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] net664 VPWR
+ VGND sg13g2_nand2_1
XFILLER_7_551 VPWR VGND sg13g2_decap_8
XFILLER_11_580 VPWR VGND sg13g2_decap_8
X_3431_ _0930_ _0953_ _0908_ _0955_ VPWR VGND sg13g2_nand3_1
X_3362_ net591 _0888_ _0889_ VPWR VGND sg13g2_nor2_1
X_2313_ _1574_ VPWR _1733_ VGND net752 _1727_ sg13g2_o21ai_1
X_3293_ VGND VPWR _0821_ _0819_ _0818_ sg13g2_or2_1
XFILLER_39_901 VPWR VGND sg13g2_decap_8
X_2244_ VGND VPWR _1573_ net730 _1664_ _1598_ sg13g2_a21oi_1
X_2175_ _1512_ _1591_ _1594_ _1595_ VPWR VGND sg13g2_nor3_2
XFILLER_39_978 VPWR VGND sg13g2_decap_8
XFILLER_26_639 VPWR VGND sg13g2_decap_8
XFILLER_25_149 VPWR VGND sg13g2_fill_1
XFILLER_38_499 VPWR VGND sg13g2_decap_8
XFILLER_41_609 VPWR VGND sg13g2_decap_8
XFILLER_15_28 VPWR VGND sg13g2_fill_1
XFILLER_34_661 VPWR VGND sg13g2_decap_8
XFILLER_22_867 VPWR VGND sg13g2_decap_8
X_3629_ _1054_ _1055_ _1121_ _1130_ VPWR VGND sg13g2_nor3_1
Xoutput27 net27 uo_out[2] VPWR VGND sg13g2_buf_1
Xoutput16 net16 uio_oe[7] VPWR VGND sg13g2_buf_1
XFILLER_1_738 VPWR VGND sg13g2_decap_8
XFILLER_5_1001 VPWR VGND sg13g2_decap_8
XFILLER_44_414 VPWR VGND sg13g2_decap_8
XFILLER_17_606 VPWR VGND sg13g2_decap_8
XFILLER_13_823 VPWR VGND sg13g2_decap_8
XFILLER_25_694 VPWR VGND sg13g2_decap_8
XFILLER_40_653 VPWR VGND sg13g2_decap_8
XFILLER_9_805 VPWR VGND sg13g2_decap_8
XFILLER_8_337 VPWR VGND sg13g2_fill_1
XFILLER_4_543 VPWR VGND sg13g2_decap_8
XFILLER_39_219 VPWR VGND sg13g2_fill_2
XFILLER_48_731 VPWR VGND sg13g2_decap_8
XFILLER_36_948 VPWR VGND sg13g2_decap_8
X_3980_ _1396_ sap_3_inst.alu.act\[1\] net582 VPWR VGND sg13g2_nand2_1
XFILLER_16_661 VPWR VGND sg13g2_decap_8
XFILLER_44_981 VPWR VGND sg13g2_decap_8
X_2931_ _0487_ _0485_ _0486_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_2862_ _0419_ VPWR _0420_ VGND net799 _0324_ sg13g2_o21ai_1
XFILLER_31_675 VPWR VGND sg13g2_decap_8
X_2793_ VPWR VGND _0353_ net580 _0352_ net31 _0354_ net626 sg13g2_a221oi_1
XFILLER_7_40 VPWR VGND sg13g2_fill_2
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_392 VPWR VGND sg13g2_fill_1
X_3414_ _0287_ _0869_ _0939_ VPWR VGND sg13g2_and2_1
Xfanout806 sap_3_inst.alu.acc\[0\] net806 VPWR VGND sg13g2_buf_8
Xfanout828 net829 net828 VPWR VGND sg13g2_buf_8
Xfanout839 net840 net839 VPWR VGND sg13g2_buf_1
X_3345_ _0873_ net652 _0827_ VPWR VGND sg13g2_nand2_2
Xfanout817 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[0\] net817 VPWR VGND
+ sg13g2_buf_2
X_3276_ _0804_ _0741_ _0803_ VPWR VGND sg13g2_nand2_1
X_2227_ _1647_ _1534_ net747 VPWR VGND sg13g2_nand2_1
Xclkbuf_4_0_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_0_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_39_775 VPWR VGND sg13g2_decap_8
X_2158_ _1575_ net731 _1578_ VPWR VGND sg13g2_nor2_1
XFILLER_26_436 VPWR VGND sg13g2_decap_8
XFILLER_27_959 VPWR VGND sg13g2_decap_8
XFILLER_38_274 VPWR VGND sg13g2_fill_2
X_2089_ _1506_ _1508_ _1509_ VPWR VGND sg13g2_nor2_1
XFILLER_22_664 VPWR VGND sg13g2_decap_8
XFILLER_10_837 VPWR VGND sg13g2_decap_8
XFILLER_1_535 VPWR VGND sg13g2_decap_8
XFILLER_18_959 VPWR VGND sg13g2_decap_8
XFILLER_29_285 VPWR VGND sg13g2_fill_1
XFILLER_45_767 VPWR VGND sg13g2_decap_8
XFILLER_9_602 VPWR VGND sg13g2_decap_8
XFILLER_13_620 VPWR VGND sg13g2_decap_8
XFILLER_25_491 VPWR VGND sg13g2_decap_8
XFILLER_41_973 VPWR VGND sg13g2_decap_8
XFILLER_12_141 VPWR VGND sg13g2_fill_1
XFILLER_8_145 VPWR VGND sg13g2_fill_2
XFILLER_12_196 VPWR VGND sg13g2_fill_2
XFILLER_13_697 VPWR VGND sg13g2_decap_8
XFILLER_9_679 VPWR VGND sg13g2_decap_8
XFILLER_32_81 VPWR VGND sg13g2_fill_1
XFILLER_5_896 VPWR VGND sg13g2_decap_8
X_3130_ _0658_ _0654_ _0656_ VPWR VGND sg13g2_nand2_2
X_3061_ sap_3_inst.alu.tmp\[7\] net24 net716 _0057_ VPWR VGND sg13g2_mux2_1
XFILLER_36_745 VPWR VGND sg13g2_decap_8
XFILLER_17_970 VPWR VGND sg13g2_decap_8
XFILLER_23_428 VPWR VGND sg13g2_decap_8
X_3963_ _1385_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] net608 VPWR
+ VGND sg13g2_nand2_1
XFILLER_32_951 VPWR VGND sg13g2_decap_8
X_2914_ net574 _0454_ _0456_ _0470_ _0471_ VPWR VGND sg13g2_nor4_1
X_3894_ _1326_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] net810
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2845_ VPWR VGND net800 _0397_ net682 net804 _0404_ net683 sg13g2_a221oi_1
X_2776_ net625 net574 _0335_ _0337_ VPWR VGND sg13g2_or3_1
Xfanout614 net615 net614 VPWR VGND sg13g2_buf_1
Xfanout603 net604 net603 VPWR VGND sg13g2_buf_8
Xfanout658 net659 net658 VPWR VGND sg13g2_buf_1
X_3328_ _1753_ VPWR _0856_ VGND _1576_ _1638_ sg13g2_o21ai_1
Xfanout625 _0332_ net625 VPWR VGND sg13g2_buf_8
Xfanout636 _1808_ net636 VPWR VGND sg13g2_buf_8
Xfanout647 _1802_ net647 VPWR VGND sg13g2_buf_8
Xfanout669 net670 net669 VPWR VGND sg13g2_buf_8
X_3259_ _0780_ _0781_ _0779_ _0787_ VPWR VGND _0783_ sg13g2_nand4_1
XFILLER_2_1015 VPWR VGND sg13g2_decap_8
XFILLER_39_572 VPWR VGND sg13g2_decap_8
XFILLER_27_756 VPWR VGND sg13g2_decap_8
XFILLER_42_737 VPWR VGND sg13g2_decap_8
XFILLER_41_247 VPWR VGND sg13g2_fill_2
XFILLER_22_461 VPWR VGND sg13g2_decap_8
XFILLER_10_634 VPWR VGND sg13g2_decap_8
XFILLER_23_995 VPWR VGND sg13g2_decap_8
XFILLER_6_649 VPWR VGND sg13g2_decap_8
XFILLER_2_833 VPWR VGND sg13g2_decap_8
XFILLER_49_358 VPWR VGND sg13g2_decap_8
XFILLER_40_1010 VPWR VGND sg13g2_decap_8
XFILLER_45_564 VPWR VGND sg13g2_decap_8
XFILLER_18_756 VPWR VGND sg13g2_decap_8
XFILLER_14_940 VPWR VGND sg13g2_decap_8
XFILLER_41_770 VPWR VGND sg13g2_decap_8
XFILLER_13_483 VPWR VGND sg13g2_fill_1
XFILLER_13_494 VPWR VGND sg13g2_decap_8
X_2630_ _0219_ net633 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] net635
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2561_ _1972_ VPWR _1973_ VGND _1445_ net629 sg13g2_o21ai_1
X_2492_ _1908_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] net637
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_693 VPWR VGND sg13g2_decap_8
X_4231_ net836 VGND VPWR _0194_ u_ser.bit_pos\[1\] clknet_3_2__leaf_clk sg13g2_dfrbpq_2
X_4162_ net845 VGND VPWR _0126_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\]
+ clknet_5_25__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3113_ _1530_ VPWR _0641_ VGND sap_3_inst.controller.stage\[1\] _1506_ sg13g2_o21ai_1
X_4093_ net839 VGND VPWR _0057_ sap_3_inst.alu.tmp\[7\] clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3044_ _1945_ _0203_ _0589_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_542 VPWR VGND sg13g2_decap_8
XFILLER_23_203 VPWR VGND sg13g2_fill_1
XFILLER_24_748 VPWR VGND sg13g2_decap_8
XFILLER_17_1012 VPWR VGND sg13g2_decap_8
X_3946_ VPWR VGND _1372_ net812 _1368_ _1484_ _1373_ net807 sg13g2_a221oi_1
X_3877_ sap_3_inst.reg_file.array_serializer_inst.word_index\[3\] sap_3_inst.reg_file.array_serializer_inst.word_index\[2\]
+ _1302_ _1310_ VPWR VGND sg13g2_nor3_1
XFILLER_20_976 VPWR VGND sg13g2_decap_8
X_2828_ _0384_ _0386_ _0387_ VPWR VGND sg13g2_nor2_1
X_2759_ VGND VPWR _0317_ _0319_ _0320_ _0316_ sg13g2_a21oi_1
XFILLER_27_553 VPWR VGND sg13g2_decap_8
XFILLER_14_203 VPWR VGND sg13g2_fill_1
XFILLER_42_534 VPWR VGND sg13g2_decap_8
XFILLER_14_214 VPWR VGND sg13g2_fill_1
XFILLER_23_792 VPWR VGND sg13g2_decap_8
XFILLER_11_965 VPWR VGND sg13g2_decap_8
XFILLER_7_936 VPWR VGND sg13g2_decap_8
XFILLER_2_630 VPWR VGND sg13g2_decap_8
XFILLER_38_807 VPWR VGND sg13g2_decap_8
XFILLER_18_553 VPWR VGND sg13g2_decap_8
XFILLER_46_884 VPWR VGND sg13g2_decap_8
XFILLER_45_361 VPWR VGND sg13g2_decap_8
XFILLER_21_718 VPWR VGND sg13g2_decap_8
X_3800_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\] net661 _1253_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_33_567 VPWR VGND sg13g2_decap_8
X_3731_ _1204_ VPWR _0119_ VGND _1159_ _1205_ sg13g2_o21ai_1
Xclkload10 VPWR clkload10/Y clknet_5_3__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_3662_ _1099_ _1100_ _1154_ VPWR VGND sg13g2_and2_1
X_2613_ _0202_ net775 _1947_ VPWR VGND sg13g2_nand2_1
X_3593_ net713 VPWR _1101_ VGND net13 _1076_ sg13g2_o21ai_1
X_2544_ _1952_ net721 _1954_ _1956_ VPWR VGND sg13g2_or3_1
XFILLER_47_1005 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_5_490 VPWR VGND sg13g2_decap_8
X_2475_ _1891_ net640 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] net643
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4214_ net832 VGND VPWR _0177_ sap_3_inst.alu.act\[0\] clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_4145_ net833 VGND VPWR _0109_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\]
+ clknet_5_18__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_818 VPWR VGND sg13g2_decap_8
X_4076_ net839 VGND VPWR _0040_ sap_3_inst.alu.acc\[7\] clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3027_ net790 sap_3_inst.out\[6\] net718 _0047_ VPWR VGND sg13g2_mux2_1
XFILLER_37_884 VPWR VGND sg13g2_decap_8
XFILLER_24_545 VPWR VGND sg13g2_decap_8
XFILLER_12_707 VPWR VGND sg13g2_decap_8
X_4044__9 VPWR net45 clknet_leaf_2_sap_3_inst.alu.clk VGND sg13g2_inv_1
Xclkload4 VPWR clkload4/Y clknet_3_5__leaf_clk VGND sg13g2_inv_1
X_3929_ net811 net50 _1357_ _0165_ VPWR VGND sg13g2_a21o_1
XFILLER_20_773 VPWR VGND sg13g2_decap_8
XFILLER_4_928 VPWR VGND sg13g2_decap_8
XFILLER_3_438 VPWR VGND sg13g2_fill_1
XFILLER_47_648 VPWR VGND sg13g2_decap_8
XFILLER_28_840 VPWR VGND sg13g2_decap_8
XFILLER_43_854 VPWR VGND sg13g2_decap_8
XFILLER_15_567 VPWR VGND sg13g2_decap_8
XFILLER_30_548 VPWR VGND sg13g2_decap_8
XFILLER_7_733 VPWR VGND sg13g2_decap_8
XFILLER_11_762 VPWR VGND sg13g2_decap_8
X_2260_ VGND VPWR net732 _1639_ _1680_ _1581_ sg13g2_a21oi_1
XFILLER_38_604 VPWR VGND sg13g2_decap_8
X_2191_ _1611_ _1600_ _1609_ VPWR VGND sg13g2_nand2_1
XFILLER_46_681 VPWR VGND sg13g2_decap_8
XFILLER_34_843 VPWR VGND sg13g2_decap_8
XFILLER_21_515 VPWR VGND sg13g2_decap_8
Xclkbuf_5_5__f_sap_3_inst.alu.clk_regs clknet_4_2_0_sap_3_inst.alu.clk_regs clknet_5_5__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3714_ _1195_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] net579 VPWR
+ VGND sg13g2_nand2_1
X_3645_ _1080_ VPWR _1141_ VGND _0663_ _0789_ sg13g2_o21ai_1
X_3576_ net18 net684 _1087_ VPWR VGND sg13g2_nor2b_1
X_2527_ net741 _1550_ _1716_ _1939_ VPWR VGND sg13g2_nor3_1
X_2458_ _1876_ _1874_ _1875_ net650 _1484_ VPWR VGND sg13g2_a22oi_1
Xhold16 u_ser.shadow_reg\[6\] VPWR VGND net65 sg13g2_dlygate4sd3_1
Xhold27 _0159_ VPWR VGND net76 sg13g2_dlygate4sd3_1
X_2389_ _1739_ _1783_ _1798_ _1809_ VPWR VGND sg13g2_nor3_2
XFILLER_29_615 VPWR VGND sg13g2_decap_8
XFILLER_21_1019 VPWR VGND sg13g2_decap_8
X_4128_ net841 VGND VPWR _0092_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\]
+ clknet_5_29__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4059_ net822 VGND VPWR _0027_ sap_3_inst.alu.flags\[2\] net40 sg13g2_dfrbpq_1
XFILLER_37_681 VPWR VGND sg13g2_decap_8
XFILLER_25_876 VPWR VGND sg13g2_decap_8
XFILLER_40_835 VPWR VGND sg13g2_decap_8
XFILLER_12_504 VPWR VGND sg13g2_decap_8
XFILLER_20_570 VPWR VGND sg13g2_decap_8
XFILLER_4_725 VPWR VGND sg13g2_decap_8
XFILLER_10_51 VPWR VGND sg13g2_fill_1
XFILLER_3_246 VPWR VGND sg13g2_fill_2
XFILLER_0_920 VPWR VGND sg13g2_decap_8
XFILLER_48_913 VPWR VGND sg13g2_decap_8
XFILLER_0_997 VPWR VGND sg13g2_decap_8
XFILLER_47_445 VPWR VGND sg13g2_decap_8
XFILLER_16_843 VPWR VGND sg13g2_decap_8
XFILLER_43_651 VPWR VGND sg13g2_decap_8
XFILLER_30_301 VPWR VGND sg13g2_fill_2
Xclkbuf_5_12__f_sap_3_inst.alu.clk_regs clknet_4_6_0_sap_3_inst.alu.clk_regs clknet_5_12__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_31_857 VPWR VGND sg13g2_decap_8
XFILLER_7_530 VPWR VGND sg13g2_decap_8
X_3430_ VPWR _0954_ _0953_ VGND sg13g2_inv_1
X_3361_ _0841_ _0883_ _0710_ _0888_ VPWR VGND sg13g2_nand3_1
X_2312_ VGND VPWR _1639_ net727 _1732_ net748 sg13g2_a21oi_1
X_3292_ _0818_ _0819_ _0820_ VPWR VGND sg13g2_nor2_2
X_2243_ VGND VPWR _1573_ _1654_ _1663_ net751 sg13g2_a21oi_1
X_2174_ _1594_ net773 VPWR VGND net774 sg13g2_nand2b_2
XFILLER_39_957 VPWR VGND sg13g2_decap_8
XFILLER_26_618 VPWR VGND sg13g2_decap_8
XFILLER_38_478 VPWR VGND sg13g2_decap_8
XFILLER_34_640 VPWR VGND sg13g2_decap_8
XFILLER_22_846 VPWR VGND sg13g2_decap_8
X_3628_ VGND VPWR _1122_ _1129_ _0092_ _1128_ sg13g2_a21oi_1
Xoutput17 net31 uio_out[0] VPWR VGND sg13g2_buf_1
Xoutput28 net28 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_717 VPWR VGND sg13g2_decap_8
X_3559_ net598 _1042_ _1072_ VPWR VGND sg13g2_nor2_1
XFILLER_29_489 VPWR VGND sg13g2_decap_8
XFILLER_45_949 VPWR VGND sg13g2_decap_8
XFILLER_13_802 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_sap_3_inst.alu.clk clknet_0_sap_3_inst.alu.clk clknet_1_1__leaf_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_12_301 VPWR VGND sg13g2_fill_1
XFILLER_25_673 VPWR VGND sg13g2_decap_8
XFILLER_40_632 VPWR VGND sg13g2_decap_8
XFILLER_12_323 VPWR VGND sg13g2_fill_1
XFILLER_12_356 VPWR VGND sg13g2_fill_2
XFILLER_13_879 VPWR VGND sg13g2_decap_8
XFILLER_4_522 VPWR VGND sg13g2_decap_8
XFILLER_4_599 VPWR VGND sg13g2_decap_8
XFILLER_48_710 VPWR VGND sg13g2_decap_8
XFILLER_0_794 VPWR VGND sg13g2_decap_8
XFILLER_48_787 VPWR VGND sg13g2_decap_8
XFILLER_36_927 VPWR VGND sg13g2_decap_8
XFILLER_47_297 VPWR VGND sg13g2_decap_8
XFILLER_44_960 VPWR VGND sg13g2_decap_8
XFILLER_16_640 VPWR VGND sg13g2_decap_8
X_2930_ VGND VPWR _0452_ _0457_ _0486_ _0450_ sg13g2_a21oi_1
XFILLER_31_654 VPWR VGND sg13g2_decap_8
X_2861_ sap_3_inst.alu.tmp\[3\] _0344_ net798 _0419_ VPWR VGND sg13g2_nand3_1
X_2792_ net626 _0351_ _0353_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1007 VPWR VGND sg13g2_decap_8
XFILLER_8_894 VPWR VGND sg13g2_decap_8
X_3413_ net606 _0937_ _0938_ VPWR VGND sg13g2_and2_1
Xfanout807 net808 net807 VPWR VGND sg13g2_buf_8
Xfanout829 net830 net829 VPWR VGND sg13g2_buf_8
Xfanout818 net820 net818 VPWR VGND sg13g2_buf_8
X_3344_ net653 net712 _0872_ VPWR VGND sg13g2_nor2_2
XFILLER_30_0 VPWR VGND sg13g2_fill_2
X_3275_ _0755_ _0802_ _0803_ VPWR VGND sg13g2_and2_1
X_2226_ net761 _1645_ _1646_ VPWR VGND sg13g2_nor2_1
XFILLER_39_754 VPWR VGND sg13g2_decap_8
X_2157_ _1577_ _1536_ net754 VPWR VGND sg13g2_nand2_2
XFILLER_26_415 VPWR VGND sg13g2_decap_8
XFILLER_27_938 VPWR VGND sg13g2_decap_8
XFILLER_42_919 VPWR VGND sg13g2_decap_8
X_2088_ _1508_ sap_3_inst.controller.stage\[1\] net761 VPWR VGND sg13g2_nand2_2
XFILLER_22_643 VPWR VGND sg13g2_decap_8
XFILLER_10_816 VPWR VGND sg13g2_decap_8
XFILLER_1_514 VPWR VGND sg13g2_decap_8
XFILLER_45_746 VPWR VGND sg13g2_decap_8
XFILLER_18_938 VPWR VGND sg13g2_decap_8
XFILLER_44_256 VPWR VGND sg13g2_fill_2
XFILLER_44_267 VPWR VGND sg13g2_fill_1
XFILLER_25_470 VPWR VGND sg13g2_decap_8
XFILLER_26_982 VPWR VGND sg13g2_decap_8
XFILLER_41_952 VPWR VGND sg13g2_decap_8
XFILLER_13_676 VPWR VGND sg13g2_decap_8
XFILLER_34_1018 VPWR VGND sg13g2_decap_8
XFILLER_9_658 VPWR VGND sg13g2_decap_8
XFILLER_8_157 VPWR VGND sg13g2_fill_2
XFILLER_5_875 VPWR VGND sg13g2_decap_8
XFILLER_0_591 VPWR VGND sg13g2_decap_8
X_3060_ sap_3_inst.alu.tmp\[6\] net23 net715 _0056_ VPWR VGND sg13g2_mux2_1
XFILLER_48_584 VPWR VGND sg13g2_decap_8
XFILLER_36_724 VPWR VGND sg13g2_decap_8
XFILLER_23_407 VPWR VGND sg13g2_decap_8
X_3962_ VGND VPWR net657 _1129_ _0171_ _1384_ sg13g2_a21oi_1
XFILLER_32_930 VPWR VGND sg13g2_decap_8
X_2913_ _0469_ VPWR _0470_ VGND _0328_ _0460_ sg13g2_o21ai_1
X_3893_ _1325_ _1301_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] _1300_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_31_440 VPWR VGND sg13g2_decap_4
X_2844_ _0403_ _0390_ _0326_ _0384_ _0335_ VPWR VGND sg13g2_a22oi_1
XFILLER_8_691 VPWR VGND sg13g2_decap_8
X_2775_ VGND VPWR _0336_ _0319_ _1951_ sg13g2_or2_1
Xfanout615 _0703_ net615 VPWR VGND sg13g2_buf_8
Xfanout604 _0833_ net604 VPWR VGND sg13g2_buf_2
Xfanout626 net627 net626 VPWR VGND sg13g2_buf_8
X_3327_ _0855_ _1551_ _0611_ VPWR VGND sg13g2_nand2_1
Xfanout648 _1801_ net648 VPWR VGND sg13g2_buf_8
Xfanout637 _1808_ net637 VPWR VGND sg13g2_buf_8
Xfanout659 _0704_ net659 VPWR VGND sg13g2_buf_8
X_3258_ _0782_ _0784_ _0778_ _0786_ VPWR VGND sg13g2_nand3_1
XFILLER_39_551 VPWR VGND sg13g2_decap_8
X_3189_ _0714_ VPWR _0717_ VGND _1499_ net620 sg13g2_o21ai_1
X_2209_ _1629_ net778 _1628_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_735 VPWR VGND sg13g2_decap_8
XFILLER_42_716 VPWR VGND sg13g2_decap_8
XFILLER_41_215 VPWR VGND sg13g2_fill_1
XFILLER_23_974 VPWR VGND sg13g2_decap_8
XFILLER_10_613 VPWR VGND sg13g2_decap_8
XFILLER_6_628 VPWR VGND sg13g2_decap_8
XFILLER_2_812 VPWR VGND sg13g2_decap_8
XFILLER_1_300 VPWR VGND sg13g2_fill_1
XFILLER_2_889 VPWR VGND sg13g2_decap_8
XFILLER_49_337 VPWR VGND sg13g2_decap_8
XFILLER_18_735 VPWR VGND sg13g2_decap_8
XFILLER_45_543 VPWR VGND sg13g2_decap_8
XFILLER_33_749 VPWR VGND sg13g2_decap_8
XFILLER_13_451 VPWR VGND sg13g2_fill_2
XFILLER_43_81 VPWR VGND sg13g2_fill_1
XFILLER_14_996 VPWR VGND sg13g2_decap_8
X_2560_ _1972_ _1858_ net4 _1839_ sap_3_inst.alu.flags\[3\] VPWR VGND sg13g2_a22oi_1
X_2491_ _1907_ net640 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] net647
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_672 VPWR VGND sg13g2_decap_8
X_4230_ net836 VGND VPWR _0193_ u_ser.bit_pos\[0\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
X_4161_ net822 VGND VPWR _0125_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\]
+ clknet_5_7__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3112_ _0639_ VPWR _0640_ VGND _0624_ _0634_ sg13g2_o21ai_1
X_4092_ net839 VGND VPWR _0056_ sap_3_inst.alu.tmp\[6\] clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3043_ _0578_ _0579_ _0587_ _0588_ VPWR VGND sg13g2_nor3_1
XFILLER_36_521 VPWR VGND sg13g2_decap_8
XFILLER_48_381 VPWR VGND sg13g2_decap_8
XFILLER_24_727 VPWR VGND sg13g2_decap_8
XFILLER_36_598 VPWR VGND sg13g2_decap_8
X_3945_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] _1371_
+ net809 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] _1372_ _1308_ sg13g2_a221oi_1
X_3876_ _1299_ _1303_ _1309_ VPWR VGND sg13g2_nor2_2
XFILLER_20_955 VPWR VGND sg13g2_decap_8
X_2827_ VGND VPWR _0357_ _0358_ _0386_ _0385_ sg13g2_a21oi_1
X_2758_ VGND VPWR _0319_ _1957_ _1955_ sg13g2_or2_1
X_2689_ VPWR VGND _1638_ _0271_ _0270_ net750 _0272_ _1644_ sg13g2_a221oi_1
XFILLER_48_15 VPWR VGND sg13g2_decap_8
XFILLER_48_26 VPWR VGND sg13g2_fill_2
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_532 VPWR VGND sg13g2_decap_8
XFILLER_42_513 VPWR VGND sg13g2_decap_8
XFILLER_15_749 VPWR VGND sg13g2_decap_8
XFILLER_23_771 VPWR VGND sg13g2_decap_8
XFILLER_7_915 VPWR VGND sg13g2_decap_8
XFILLER_11_944 VPWR VGND sg13g2_decap_8
XFILLER_10_487 VPWR VGND sg13g2_decap_8
XFILLER_2_686 VPWR VGND sg13g2_decap_8
XFILLER_18_532 VPWR VGND sg13g2_decap_8
XFILLER_46_863 VPWR VGND sg13g2_decap_8
XFILLER_33_546 VPWR VGND sg13g2_decap_8
X_3730_ _1205_ net665 _1191_ VPWR VGND sg13g2_nand2_1
XFILLER_14_793 VPWR VGND sg13g2_decap_8
X_3661_ _0101_ _0935_ _1153_ net623 _1450_ VPWR VGND sg13g2_a22oi_1
X_2612_ VGND VPWR _0201_ _1950_ net714 sg13g2_or2_1
Xclkload11 VPWR clkload11/Y clknet_5_5__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_3592_ _1100_ net607 _0962_ VPWR VGND sg13g2_nand2_1
X_2543_ _1952_ net721 _1954_ _1955_ VPWR VGND sg13g2_nor3_2
XFILLER_47_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_992 VPWR VGND sg13g2_decap_8
X_2474_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[5\] _1801_ _1890_ VPWR
+ VGND sg13g2_nor2_1
X_4213_ net831 VGND VPWR net37 clk_div_out clknet_3_0__leaf_clk sg13g2_dfrbpq_1
X_4144_ net842 VGND VPWR _0108_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\]
+ clknet_5_29__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_307 VPWR VGND sg13g2_fill_2
X_4075_ net839 VGND VPWR _0039_ sap_3_inst.alu.acc\[6\] clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3026_ net793 sap_3_inst.out\[5\] net718 _0046_ VPWR VGND sg13g2_mux2_1
XFILLER_37_863 VPWR VGND sg13g2_decap_8
XFILLER_24_524 VPWR VGND sg13g2_decap_8
XFILLER_20_752 VPWR VGND sg13g2_decap_8
Xclkload5 VPWR clkload5/Y clknet_3_6__leaf_clk VGND sg13g2_inv_1
X_3928_ VPWR VGND _1356_ net811 _1352_ _1474_ _1357_ net808 sg13g2_a221oi_1
XFILLER_30_1010 VPWR VGND sg13g2_decap_8
X_3859_ _1292_ VPWR _1293_ VGND sap_3_inst.reg_file.array_serializer_inst.bit_pos\[0\]
+ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[5\] sg13g2_o21ai_1
XFILLER_4_907 VPWR VGND sg13g2_decap_8
XFILLER_47_627 VPWR VGND sg13g2_decap_8
XFILLER_43_833 VPWR VGND sg13g2_decap_8
XFILLER_28_896 VPWR VGND sg13g2_decap_8
XFILLER_15_546 VPWR VGND sg13g2_decap_8
XFILLER_30_527 VPWR VGND sg13g2_decap_8
XFILLER_11_741 VPWR VGND sg13g2_decap_8
XFILLER_7_712 VPWR VGND sg13g2_decap_8
XFILLER_7_789 VPWR VGND sg13g2_decap_8
XFILLER_3_995 VPWR VGND sg13g2_decap_8
XFILLER_2_483 VPWR VGND sg13g2_decap_8
X_2190_ net750 _1608_ _1610_ VPWR VGND sg13g2_nor2_2
XFILLER_46_660 VPWR VGND sg13g2_decap_8
XFILLER_19_885 VPWR VGND sg13g2_decap_8
XFILLER_34_822 VPWR VGND sg13g2_decap_8
XFILLER_34_899 VPWR VGND sg13g2_decap_8
XFILLER_14_590 VPWR VGND sg13g2_decap_8
X_3713_ _0112_ _1194_ _1065_ net578 _1490_ VPWR VGND sg13g2_a22oi_1
X_3644_ _1138_ net17 _1139_ _1140_ VPWR VGND sg13g2_a21o_1
X_3575_ net605 _0886_ _1086_ VPWR VGND sg13g2_nor2_1
X_2526_ net724 _1935_ _1937_ _1938_ VPWR VGND sg13g2_nor3_1
XFILLER_0_409 VPWR VGND sg13g2_fill_1
X_2457_ net648 _1869_ _1870_ _1871_ _1875_ VPWR VGND sg13g2_and4_1
Xhold17 u_ser.shadow_reg\[5\] VPWR VGND net66 sg13g2_dlygate4sd3_1
XFILLER_29_28 VPWR VGND sg13g2_fill_1
XFILLER_29_39 VPWR VGND sg13g2_fill_1
Xhold28 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\] VPWR VGND net77 sg13g2_dlygate4sd3_1
X_2388_ _1766_ _1783_ _1799_ _1808_ VPWR VGND sg13g2_nor3_2
X_4127_ net820 VGND VPWR _0091_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\]
+ clknet_5_1__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4058_ net834 VGND VPWR _0026_ sap_3_inst.alu.flags\[1\] net39 sg13g2_dfrbpq_2
XFILLER_37_660 VPWR VGND sg13g2_decap_8
X_3009_ _0562_ _0526_ _0563_ VPWR VGND sg13g2_xor2_1
XFILLER_25_855 VPWR VGND sg13g2_decap_8
XFILLER_40_814 VPWR VGND sg13g2_decap_8
XFILLER_8_509 VPWR VGND sg13g2_decap_8
XFILLER_24_398 VPWR VGND sg13g2_decap_8
XFILLER_4_704 VPWR VGND sg13g2_decap_8
XFILLER_3_214 VPWR VGND sg13g2_fill_1
XFILLER_10_74 VPWR VGND sg13g2_fill_2
XFILLER_0_976 VPWR VGND sg13g2_decap_8
XFILLER_48_969 VPWR VGND sg13g2_decap_8
XFILLER_47_424 VPWR VGND sg13g2_decap_8
XFILLER_19_148 VPWR VGND sg13g2_fill_2
XFILLER_35_619 VPWR VGND sg13g2_decap_8
XFILLER_16_822 VPWR VGND sg13g2_decap_8
XFILLER_27_170 VPWR VGND sg13g2_fill_1
XFILLER_28_693 VPWR VGND sg13g2_decap_8
XFILLER_43_630 VPWR VGND sg13g2_decap_8
XFILLER_16_899 VPWR VGND sg13g2_decap_8
XFILLER_31_836 VPWR VGND sg13g2_decap_8
XFILLER_7_586 VPWR VGND sg13g2_decap_8
X_3360_ net606 _0886_ _0887_ VPWR VGND sg13g2_and2_1
XFILLER_44_1009 VPWR VGND sg13g2_decap_8
X_2311_ VGND VPWR _1657_ _1729_ _1731_ _1610_ sg13g2_a21oi_1
XFILLER_3_792 VPWR VGND sg13g2_decap_8
X_3291_ _1535_ VPWR _0819_ VGND net776 _0636_ sg13g2_o21ai_1
X_2242_ VGND VPWR net732 _1648_ _1662_ net749 sg13g2_a21oi_1
XFILLER_39_936 VPWR VGND sg13g2_decap_8
X_2173_ net774 net772 _1593_ VPWR VGND sg13g2_nor2b_2
XFILLER_38_468 VPWR VGND sg13g2_fill_1
XFILLER_47_991 VPWR VGND sg13g2_decap_8
XFILLER_18_170 VPWR VGND sg13g2_fill_2
XFILLER_19_682 VPWR VGND sg13g2_decap_8
XFILLER_22_825 VPWR VGND sg13g2_decap_8
XFILLER_34_696 VPWR VGND sg13g2_decap_8
XFILLER_30_891 VPWR VGND sg13g2_decap_8
X_3627_ VPWR VGND _0835_ _1052_ _0918_ net601 _1129_ _0911_ sg13g2_a221oi_1
X_3558_ _1071_ _1069_ _1070_ VPWR VGND sg13g2_nand2b_1
Xoutput18 net18 uio_out[1] VPWR VGND sg13g2_buf_1
Xoutput29 net29 uo_out[4] VPWR VGND sg13g2_buf_1
X_2509_ _1923_ net628 _1922_ VPWR VGND sg13g2_nand2_1
X_3489_ VGND VPWR net669 _1008_ _1011_ _1010_ sg13g2_a21oi_1
XFILLER_45_928 VPWR VGND sg13g2_decap_8
XFILLER_44_449 VPWR VGND sg13g2_decap_8
XFILLER_25_652 VPWR VGND sg13g2_decap_8
XFILLER_40_611 VPWR VGND sg13g2_decap_8
XFILLER_13_858 VPWR VGND sg13g2_decap_8
XFILLER_40_688 VPWR VGND sg13g2_decap_8
XFILLER_4_501 VPWR VGND sg13g2_decap_8
XFILLER_4_578 VPWR VGND sg13g2_decap_8
XFILLER_0_773 VPWR VGND sg13g2_decap_8
XFILLER_48_766 VPWR VGND sg13g2_decap_8
XFILLER_36_906 VPWR VGND sg13g2_decap_8
XFILLER_28_490 VPWR VGND sg13g2_decap_8
X_2860_ _0418_ net798 sap_3_inst.alu.tmp\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_16_696 VPWR VGND sg13g2_decap_8
XFILLER_31_633 VPWR VGND sg13g2_decap_8
X_2791_ _0352_ net708 sap_3_inst.alu.act\[0\] VPWR VGND sg13g2_nand2b_1
XFILLER_8_873 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_fill_1
X_3412_ _0937_ _0913_ _0930_ VPWR VGND sg13g2_xnor2_1
Xfanout819 net820 net819 VPWR VGND sg13g2_buf_8
X_3343_ _0848_ net587 _0870_ _0871_ VPWR VGND sg13g2_nor3_1
Xfanout808 _1313_ net808 VPWR VGND sg13g2_buf_8
X_3274_ _0766_ _0775_ net591 net588 _0802_ VPWR VGND sg13g2_and4_1
X_2225_ _1645_ net760 net747 VPWR VGND sg13g2_nand2_1
XFILLER_39_733 VPWR VGND sg13g2_decap_8
XFILLER_27_917 VPWR VGND sg13g2_decap_8
X_2156_ _1536_ _1557_ _1576_ VPWR VGND sg13g2_and2_1
X_2087_ net760 net761 _1507_ VPWR VGND sg13g2_and2_1
XFILLER_35_983 VPWR VGND sg13g2_decap_8
XFILLER_22_622 VPWR VGND sg13g2_decap_8
XFILLER_34_493 VPWR VGND sg13g2_decap_8
X_2989_ _0543_ net788 net721 VPWR VGND sg13g2_xnor2_1
XFILLER_22_699 VPWR VGND sg13g2_decap_8
XFILLER_27_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_519 VPWR VGND sg13g2_decap_8
XFILLER_18_917 VPWR VGND sg13g2_decap_8
XFILLER_45_725 VPWR VGND sg13g2_decap_8
XFILLER_44_213 VPWR VGND sg13g2_fill_2
XFILLER_26_961 VPWR VGND sg13g2_decap_8
XFILLER_41_931 VPWR VGND sg13g2_decap_8
XFILLER_13_655 VPWR VGND sg13g2_decap_8
XFILLER_9_637 VPWR VGND sg13g2_decap_8
XFILLER_40_485 VPWR VGND sg13g2_decap_8
XFILLER_5_854 VPWR VGND sg13g2_decap_8
XFILLER_0_570 VPWR VGND sg13g2_decap_8
XFILLER_48_563 VPWR VGND sg13g2_decap_8
XFILLER_36_703 VPWR VGND sg13g2_decap_8
XFILLER_24_909 VPWR VGND sg13g2_decap_8
X_3961_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] net657 _1384_ VPWR
+ VGND sg13g2_nor2_1
X_2912_ VGND VPWR _0326_ _0465_ _0469_ _0468_ sg13g2_a21oi_1
XFILLER_16_493 VPWR VGND sg13g2_decap_8
XFILLER_32_986 VPWR VGND sg13g2_decap_8
X_3892_ net811 net54 _1324_ _0161_ VPWR VGND sg13g2_a21o_1
X_2843_ _0391_ VPWR _0402_ VGND net802 _0324_ sg13g2_o21ai_1
X_2774_ _1951_ _0319_ _0335_ VPWR VGND sg13g2_nor2_2
XFILLER_8_670 VPWR VGND sg13g2_decap_8
Xfanout605 _0829_ net605 VPWR VGND sg13g2_buf_8
Xfanout616 net617 net616 VPWR VGND sg13g2_buf_8
X_3326_ _0629_ VPWR _0854_ VGND net765 _1850_ sg13g2_o21ai_1
Xfanout627 _0311_ net627 VPWR VGND sg13g2_buf_8
Xfanout649 _1800_ net649 VPWR VGND sg13g2_buf_8
Xfanout638 net639 net638 VPWR VGND sg13g2_buf_8
X_3257_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] net676 _0785_ VPWR
+ VGND sg13g2_and2_1
XFILLER_39_530 VPWR VGND sg13g2_decap_8
X_2208_ net775 sap_3_inst.alu.flags\[0\] net762 sap_3_inst.alu.flags\[2\] sap_3_inst.alu.flags\[3\]
+ net773 _1628_ VPWR VGND sg13g2_mux4_1
XFILLER_27_714 VPWR VGND sg13g2_decap_8
X_3188_ _0716_ net666 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] net672
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2139_ net755 net754 _1559_ VPWR VGND sg13g2_and2_1
XFILLER_35_780 VPWR VGND sg13g2_decap_8
XFILLER_23_953 VPWR VGND sg13g2_decap_8
XFILLER_6_607 VPWR VGND sg13g2_decap_8
XFILLER_10_669 VPWR VGND sg13g2_decap_8
XFILLER_22_496 VPWR VGND sg13g2_decap_8
XFILLER_5_139 VPWR VGND sg13g2_fill_1
XFILLER_2_868 VPWR VGND sg13g2_decap_8
XFILLER_49_316 VPWR VGND sg13g2_decap_8
XFILLER_18_714 VPWR VGND sg13g2_decap_8
XFILLER_45_522 VPWR VGND sg13g2_decap_8
XFILLER_17_235 VPWR VGND sg13g2_fill_1
XFILLER_33_728 VPWR VGND sg13g2_decap_8
XFILLER_45_599 VPWR VGND sg13g2_decap_8
XFILLER_14_975 VPWR VGND sg13g2_decap_8
XFILLER_43_93 VPWR VGND sg13g2_fill_2
X_2490_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] net643
+ net638 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] _1906_ net722 sg13g2_a221oi_1
XFILLER_5_651 VPWR VGND sg13g2_decap_8
X_4160_ net841 VGND VPWR _0124_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\]
+ clknet_5_29__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3111_ VGND VPWR net725 _0638_ _0639_ _1520_ sg13g2_a21oi_1
X_4091_ net838 VGND VPWR _0055_ sap_3_inst.alu.tmp\[5\] clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_49_883 VPWR VGND sg13g2_decap_8
XFILLER_48_360 VPWR VGND sg13g2_decap_8
X_3042_ _0586_ VPWR _0587_ VGND _0582_ _0583_ sg13g2_o21ai_1
XFILLER_36_500 VPWR VGND sg13g2_decap_8
XFILLER_24_706 VPWR VGND sg13g2_decap_8
XFILLER_36_577 VPWR VGND sg13g2_decap_8
X_3944_ _1367_ _1369_ _1366_ _1371_ VPWR VGND _1370_ sg13g2_nand4_1
X_3875_ sap_3_inst.reg_file.array_serializer_inst.word_index\[1\] sap_3_inst.reg_file.array_serializer_inst.word_index\[0\]
+ _1303_ _1308_ VPWR VGND sg13g2_nor3_2
XFILLER_20_934 VPWR VGND sg13g2_decap_8
XFILLER_32_783 VPWR VGND sg13g2_decap_8
X_2826_ sap_3_inst.alu.tmp\[1\] net804 _0385_ VPWR VGND sg13g2_nor2b_1
X_2757_ _1955_ _1957_ _0318_ VPWR VGND sg13g2_nor2_1
X_2688_ _1792_ VPWR _0271_ VGND net734 _1617_ sg13g2_o21ai_1
XFILLER_24_1007 VPWR VGND sg13g2_decap_8
XFILLER_47_809 VPWR VGND sg13g2_decap_8
X_3309_ _0755_ _0766_ _0775_ _0837_ VGND VPWR net589 sg13g2_nor4_2
XFILLER_27_511 VPWR VGND sg13g2_decap_8
XFILLER_15_728 VPWR VGND sg13g2_decap_8
XFILLER_27_588 VPWR VGND sg13g2_decap_8
XFILLER_42_569 VPWR VGND sg13g2_decap_8
XFILLER_23_750 VPWR VGND sg13g2_decap_8
XFILLER_30_709 VPWR VGND sg13g2_decap_8
Xfanout31 net17 net31 VPWR VGND sg13g2_buf_2
XFILLER_11_923 VPWR VGND sg13g2_decap_8
XFILLER_2_665 VPWR VGND sg13g2_decap_8
XFILLER_49_157 VPWR VGND sg13g2_fill_1
XFILLER_18_511 VPWR VGND sg13g2_decap_8
XFILLER_46_842 VPWR VGND sg13g2_decap_8
XFILLER_45_396 VPWR VGND sg13g2_decap_8
XFILLER_18_588 VPWR VGND sg13g2_decap_8
XFILLER_33_525 VPWR VGND sg13g2_decap_8
XFILLER_14_772 VPWR VGND sg13g2_decap_8
XFILLER_13_293 VPWR VGND sg13g2_fill_2
XFILLER_9_275 VPWR VGND sg13g2_fill_1
X_3660_ net623 _0938_ _1152_ _1153_ VPWR VGND sg13g2_nor3_1
X_2611_ _0200_ _1959_ _0199_ VPWR VGND sg13g2_nand2_1
X_3591_ _1099_ net601 _0957_ VPWR VGND sg13g2_nand2_2
Xclkload12 VPWR clkload12/Y clknet_5_9__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_2542_ net748 _1633_ _1954_ VPWR VGND sg13g2_nor2_1
XFILLER_6_971 VPWR VGND sg13g2_decap_8
X_4212_ net828 VGND VPWR _0176_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\]
+ clknet_5_15__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2473_ sap_3_inst.alu.flags\[6\] net33 _1867_ _0031_ VPWR VGND sg13g2_mux2_1
X_4143_ net820 VGND VPWR _0107_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\]
+ clknet_5_6__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4074_ net838 VGND VPWR _0038_ sap_3_inst.alu.acc\[5\] clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_49_680 VPWR VGND sg13g2_decap_8
X_3025_ _0573_ VPWR _0045_ VGND _1460_ net718 sg13g2_o21ai_1
XFILLER_37_842 VPWR VGND sg13g2_decap_8
XFILLER_24_503 VPWR VGND sg13g2_decap_8
XFILLER_20_731 VPWR VGND sg13g2_decap_8
XFILLER_32_580 VPWR VGND sg13g2_decap_8
X_3927_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] _1355_
+ _1308_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\] _1356_ _1301_ sg13g2_a221oi_1
X_3858_ _1292_ net817 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[6\] VPWR
+ VGND sg13g2_nand2b_1
Xclkload6 VPWR clkload6/Y clknet_3_7__leaf_clk VGND sg13g2_inv_1
X_2809_ _0342_ VPWR _0369_ VGND net803 sap_3_inst.alu.tmp\[1\] sg13g2_o21ai_1
X_3789_ _1027_ _1012_ _1246_ VPWR VGND sg13g2_xor2_1
Xclkbuf_5_20__f_sap_3_inst.alu.clk_regs clknet_4_10_0_sap_3_inst.alu.clk_regs clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_47_606 VPWR VGND sg13g2_decap_8
XFILLER_43_812 VPWR VGND sg13g2_decap_8
XFILLER_28_875 VPWR VGND sg13g2_decap_8
XFILLER_15_525 VPWR VGND sg13g2_decap_8
XFILLER_27_385 VPWR VGND sg13g2_decap_4
XFILLER_27_396 VPWR VGND sg13g2_decap_4
XFILLER_43_889 VPWR VGND sg13g2_decap_8
XFILLER_30_506 VPWR VGND sg13g2_decap_8
XFILLER_11_720 VPWR VGND sg13g2_decap_8
XFILLER_7_768 VPWR VGND sg13g2_decap_8
XFILLER_11_797 VPWR VGND sg13g2_decap_8
XFILLER_3_974 VPWR VGND sg13g2_decap_8
XFILLER_38_639 VPWR VGND sg13g2_decap_8
XFILLER_19_864 VPWR VGND sg13g2_decap_8
XFILLER_34_801 VPWR VGND sg13g2_decap_8
XFILLER_33_300 VPWR VGND sg13g2_fill_2
XFILLER_34_878 VPWR VGND sg13g2_decap_8
X_3712_ _1132_ net578 _1194_ VPWR VGND sg13g2_nor2_1
XFILLER_14_1017 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
X_3643_ VGND VPWR _0829_ _1138_ _1139_ _1077_ sg13g2_a21oi_1
X_3574_ _1085_ net600 _0891_ VPWR VGND sg13g2_nand2_1
X_2525_ _1937_ _1936_ net748 _1633_ net734 VPWR VGND sg13g2_a22oi_1
X_2456_ _1872_ _1873_ _1874_ VPWR VGND sg13g2_and2_1
Xhold18 u_ser.shadow_reg\[4\] VPWR VGND net67 sg13g2_dlygate4sd3_1
Xhold29 sap_3_outputReg_serial VPWR VGND net78 sg13g2_dlygate4sd3_1
X_4126_ net843 VGND VPWR _0090_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\]
+ clknet_5_26__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2387_ _1766_ _1784_ _1798_ _1807_ VPWR VGND sg13g2_nor3_2
X_4057_ net833 VGND VPWR _0025_ sap_3_inst.alu.flags\[0\] net38 sg13g2_dfrbpq_1
X_3008_ _0562_ _0549_ _0561_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_834 VPWR VGND sg13g2_decap_8
XFILLER_24_377 VPWR VGND sg13g2_decap_8
XFILLER_12_539 VPWR VGND sg13g2_decap_8
XFILLER_0_955 VPWR VGND sg13g2_decap_8
XFILLER_47_403 VPWR VGND sg13g2_decap_8
XFILLER_48_948 VPWR VGND sg13g2_decap_8
XFILLER_16_801 VPWR VGND sg13g2_decap_8
XFILLER_28_672 VPWR VGND sg13g2_decap_8
XFILLER_43_686 VPWR VGND sg13g2_decap_8
XFILLER_16_878 VPWR VGND sg13g2_decap_8
XFILLER_31_815 VPWR VGND sg13g2_decap_8
XFILLER_37_1017 VPWR VGND sg13g2_decap_8
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_594 VPWR VGND sg13g2_decap_8
XFILLER_7_565 VPWR VGND sg13g2_decap_8
X_3290_ VGND VPWR _0811_ _0817_ _0818_ _0275_ sg13g2_a21oi_1
XFILLER_3_771 VPWR VGND sg13g2_decap_8
X_2310_ _1610_ _1657_ _1730_ VPWR VGND sg13g2_nor2_2
X_2241_ VGND VPWR _1661_ _1660_ _1659_ sg13g2_or2_1
XFILLER_39_915 VPWR VGND sg13g2_decap_8
X_2172_ _1512_ _1591_ _1592_ VPWR VGND sg13g2_nor2_1
XFILLER_47_970 VPWR VGND sg13g2_decap_8
XFILLER_19_661 VPWR VGND sg13g2_decap_8
XFILLER_22_804 VPWR VGND sg13g2_decap_8
XFILLER_34_675 VPWR VGND sg13g2_decap_8
XFILLER_30_870 VPWR VGND sg13g2_decap_8
X_3626_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] _1122_ _1128_ VPWR
+ VGND sg13g2_nor2_1
Xoutput19 net19 uio_out[2] VPWR VGND sg13g2_buf_1
X_3557_ _0872_ _1034_ _1070_ VPWR VGND sg13g2_and2_1
X_2508_ _1922_ sap_3_inst.alu.flags\[4\] _1839_ VPWR VGND sg13g2_nand2_1
X_3488_ net606 VPWR _1010_ VGND net669 _1009_ sg13g2_o21ai_1
X_2439_ net8 _1858_ _1859_ VPWR VGND sg13g2_and2_1
XFILLER_5_1015 VPWR VGND sg13g2_decap_8
XFILLER_45_907 VPWR VGND sg13g2_decap_8
X_4109_ net824 VGND VPWR _0073_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[7\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
XFILLER_44_428 VPWR VGND sg13g2_decap_8
XFILLER_25_631 VPWR VGND sg13g2_decap_8
XFILLER_13_837 VPWR VGND sg13g2_decap_8
XFILLER_40_667 VPWR VGND sg13g2_decap_8
XFILLER_9_819 VPWR VGND sg13g2_decap_8
XFILLER_21_30 VPWR VGND sg13g2_fill_2
XFILLER_4_557 VPWR VGND sg13g2_decap_8
Xclkbuf_5_17__f_sap_3_inst.alu.clk_regs clknet_4_8_0_sap_3_inst.alu.clk_regs clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_0_752 VPWR VGND sg13g2_decap_8
XFILLER_48_745 VPWR VGND sg13g2_decap_8
XFILLER_44_995 VPWR VGND sg13g2_decap_8
XFILLER_16_675 VPWR VGND sg13g2_decap_8
XFILLER_43_483 VPWR VGND sg13g2_decap_8
XFILLER_31_612 VPWR VGND sg13g2_decap_8
X_2790_ VPWR VGND _0330_ _0350_ _0349_ _0323_ _0351_ _0337_ sg13g2_a221oi_1
XFILLER_31_689 VPWR VGND sg13g2_decap_8
XFILLER_8_852 VPWR VGND sg13g2_decap_8
X_3411_ _0907_ _0931_ _0885_ _0936_ VPWR VGND sg13g2_nand3_1
X_3342_ net9 net31 net596 _0870_ VPWR VGND sg13g2_mux2_1
Xfanout809 _1310_ net809 VPWR VGND sg13g2_buf_8
X_3273_ _0801_ _0775_ net588 VPWR VGND sg13g2_nand2_1
X_2224_ _1507_ _1642_ _1644_ VPWR VGND sg13g2_and2_1
XFILLER_39_712 VPWR VGND sg13g2_decap_8
X_2155_ _1575_ _1568_ VPWR VGND _1564_ sg13g2_nand2b_2
XFILLER_16_0 VPWR VGND sg13g2_fill_2
XFILLER_39_789 VPWR VGND sg13g2_decap_8
X_2086_ VGND VPWR _1506_ net759 sap_3_inst.controller.stage\[3\] sg13g2_or2_1
XFILLER_38_299 VPWR VGND sg13g2_fill_1
XFILLER_22_601 VPWR VGND sg13g2_decap_8
XFILLER_35_962 VPWR VGND sg13g2_decap_8
XFILLER_42_29 VPWR VGND sg13g2_fill_2
XFILLER_22_678 VPWR VGND sg13g2_decap_8
X_2988_ _0542_ _0529_ _0534_ VPWR VGND sg13g2_nand2_1
X_3609_ net619 _1111_ _1114_ _1115_ VPWR VGND sg13g2_nor3_1
XFILLER_1_549 VPWR VGND sg13g2_decap_8
XFILLER_45_704 VPWR VGND sg13g2_decap_8
XFILLER_29_233 VPWR VGND sg13g2_decap_4
XFILLER_17_417 VPWR VGND sg13g2_fill_2
XFILLER_26_940 VPWR VGND sg13g2_decap_8
XFILLER_44_258 VPWR VGND sg13g2_fill_1
XFILLER_41_910 VPWR VGND sg13g2_decap_8
XFILLER_16_30 VPWR VGND sg13g2_fill_1
XFILLER_13_634 VPWR VGND sg13g2_decap_8
XFILLER_16_85 VPWR VGND sg13g2_fill_1
XFILLER_16_96 VPWR VGND sg13g2_fill_2
XFILLER_9_616 VPWR VGND sg13g2_decap_8
XFILLER_41_987 VPWR VGND sg13g2_decap_8
XFILLER_40_464 VPWR VGND sg13g2_decap_8
XFILLER_5_833 VPWR VGND sg13g2_decap_8
XFILLER_48_542 VPWR VGND sg13g2_decap_8
XFILLER_35_225 VPWR VGND sg13g2_fill_1
XFILLER_36_759 VPWR VGND sg13g2_decap_8
XFILLER_17_984 VPWR VGND sg13g2_decap_8
X_3960_ _1383_ VPWR _0170_ VGND _1462_ net655 sg13g2_o21ai_1
XFILLER_44_792 VPWR VGND sg13g2_decap_8
X_2911_ _0468_ _0466_ _0467_ VPWR VGND sg13g2_nand2_1
XFILLER_31_431 VPWR VGND sg13g2_fill_1
XFILLER_32_965 VPWR VGND sg13g2_decap_8
X_3891_ VPWR VGND _1323_ net812 _1319_ _1468_ _1324_ net808 sg13g2_a221oi_1
X_2842_ _0401_ _0370_ _0399_ VPWR VGND sg13g2_xnor2_1
X_2773_ _0325_ _0333_ _0334_ VPWR VGND sg13g2_and2_1
Xfanout606 net607 net606 VPWR VGND sg13g2_buf_8
X_3325_ VGND VPWR _1643_ net727 _0853_ _1610_ sg13g2_a21oi_1
Xfanout628 net629 net628 VPWR VGND sg13g2_buf_2
Xfanout639 _1807_ net639 VPWR VGND sg13g2_buf_8
Xfanout617 _0698_ net617 VPWR VGND sg13g2_buf_8
X_3256_ net699 net691 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] _0784_
+ VPWR VGND net686 sg13g2_nand4_1
X_2207_ _1442_ net772 _1627_ VPWR VGND sg13g2_nor2_1
X_3187_ _0712_ VPWR _0715_ VGND _1497_ _0666_ sg13g2_o21ai_1
XFILLER_39_586 VPWR VGND sg13g2_decap_8
X_2138_ _1558_ net759 VPWR VGND sap_3_inst.controller.stage\[3\] sg13g2_nand2b_2
X_2069_ VPWR _1491_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_23_932 VPWR VGND sg13g2_decap_8
XFILLER_22_475 VPWR VGND sg13g2_decap_8
XFILLER_10_648 VPWR VGND sg13g2_decap_8
XFILLER_2_847 VPWR VGND sg13g2_decap_8
XFILLER_45_501 VPWR VGND sg13g2_decap_8
XFILLER_40_1024 VPWR VGND sg13g2_decap_4
XFILLER_45_578 VPWR VGND sg13g2_decap_8
XFILLER_33_707 VPWR VGND sg13g2_decap_8
XFILLER_14_954 VPWR VGND sg13g2_decap_8
XFILLER_43_61 VPWR VGND sg13g2_fill_1
XFILLER_41_784 VPWR VGND sg13g2_decap_8
XFILLER_5_630 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_fill_2
XFILLER_4_195 VPWR VGND sg13g2_fill_2
XFILLER_4_55 VPWR VGND sg13g2_fill_2
X_3110_ net774 VPWR _0638_ VGND _0635_ _0637_ sg13g2_o21ai_1
X_4090_ net838 VGND VPWR _0054_ sap_3_inst.alu.tmp\[4\] clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_49_862 VPWR VGND sg13g2_decap_8
X_3041_ VPWR VGND net805 _0585_ net682 net789 _0586_ net683 sg13g2_a221oi_1
XFILLER_36_556 VPWR VGND sg13g2_decap_8
XFILLER_17_781 VPWR VGND sg13g2_decap_8
X_3943_ _1370_ _1314_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] _1300_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_17_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_913 VPWR VGND sg13g2_decap_8
XFILLER_32_762 VPWR VGND sg13g2_decap_8
X_3874_ net815 net816 _1305_ _1307_ VPWR VGND sg13g2_nor3_2
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
X_2825_ _0382_ _0383_ _0384_ VPWR VGND sg13g2_nor2b_2
XFILLER_9_980 VPWR VGND sg13g2_decap_8
X_2756_ _1947_ _1949_ _0317_ VPWR VGND sg13g2_and2_1
X_2687_ _0270_ _1570_ _1587_ VPWR VGND sg13g2_nand2_1
X_3308_ _0766_ _0835_ _0836_ VPWR VGND sg13g2_nor2_1
X_3239_ net697 net692 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] _0767_
+ VPWR VGND net688 sg13g2_nand4_1
XFILLER_15_707 VPWR VGND sg13g2_decap_8
XFILLER_27_567 VPWR VGND sg13g2_decap_8
XFILLER_42_548 VPWR VGND sg13g2_decap_8
XFILLER_11_902 VPWR VGND sg13g2_decap_8
Xfanout32 net21 net32 VPWR VGND sg13g2_buf_2
XFILLER_22_294 VPWR VGND sg13g2_fill_1
XFILLER_11_979 VPWR VGND sg13g2_decap_8
XFILLER_13_64 VPWR VGND sg13g2_fill_2
XFILLER_2_644 VPWR VGND sg13g2_decap_8
XFILLER_46_821 VPWR VGND sg13g2_decap_8
XFILLER_18_567 VPWR VGND sg13g2_decap_8
XFILLER_33_504 VPWR VGND sg13g2_decap_8
XFILLER_46_898 VPWR VGND sg13g2_decap_8
XFILLER_45_375 VPWR VGND sg13g2_decap_8
XFILLER_14_751 VPWR VGND sg13g2_decap_8
XFILLER_41_581 VPWR VGND sg13g2_decap_8
Xclkload13 VPWR clkload13/Y clknet_5_13__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_2610_ _0199_ _1947_ VPWR VGND _1949_ sg13g2_nand2b_2
X_3590_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] net667 _1098_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_6_950 VPWR VGND sg13g2_decap_8
X_2541_ _1550_ _1796_ _1953_ VPWR VGND sg13g2_nor2_1
XFILLER_47_1019 VPWR VGND sg13g2_decap_8
X_2472_ _1881_ _1889_ _1877_ net23 VPWR VGND sg13g2_nand3_1
X_4211_ net826 VGND VPWR _0175_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\]
+ clknet_5_13__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4142_ net844 VGND VPWR _0106_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4073_ net838 VGND VPWR _0037_ sap_3_inst.alu.acc\[4\] clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3024_ _0573_ sap_3_inst.out\[4\] net717 VPWR VGND sg13g2_nand2_1
XFILLER_37_821 VPWR VGND sg13g2_decap_8
XFILLER_37_898 VPWR VGND sg13g2_decap_8
XFILLER_24_559 VPWR VGND sg13g2_decap_8
XFILLER_20_710 VPWR VGND sg13g2_decap_8
X_3926_ _1351_ _1353_ _1350_ _1355_ VPWR VGND _1354_ sg13g2_nand4_1
Xclkload7 clknet_1_1__leaf_clk_div_out clkload7/X VPWR VGND sg13g2_buf_1
X_3857_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[3\] sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\]
+ _1290_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[4\] _1291_ _1279_ sg13g2_a221oi_1
X_3788_ _1245_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] net614 VPWR
+ VGND sg13g2_nand2_1
X_2808_ VPWR VGND net801 _0367_ net682 net806 _0368_ net683 sg13g2_a221oi_1
XFILLER_20_787 VPWR VGND sg13g2_decap_8
X_2739_ net729 _1715_ _1516_ _0300_ VPWR VGND sg13g2_nand3_1
XFILLER_8_1013 VPWR VGND sg13g2_decap_8
XFILLER_28_854 VPWR VGND sg13g2_decap_8
XFILLER_15_504 VPWR VGND sg13g2_decap_8
XFILLER_43_868 VPWR VGND sg13g2_decap_8
XFILLER_42_378 VPWR VGND sg13g2_decap_8
XFILLER_42_356 VPWR VGND sg13g2_decap_4
XFILLER_24_41 VPWR VGND sg13g2_fill_2
XFILLER_24_85 VPWR VGND sg13g2_fill_1
XFILLER_11_776 VPWR VGND sg13g2_decap_8
XFILLER_24_96 VPWR VGND sg13g2_fill_1
XFILLER_7_747 VPWR VGND sg13g2_decap_8
XFILLER_6_213 VPWR VGND sg13g2_fill_2
XFILLER_6_279 VPWR VGND sg13g2_fill_2
XFILLER_3_953 VPWR VGND sg13g2_decap_8
XFILLER_1_23 VPWR VGND sg13g2_fill_2
XFILLER_38_618 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_fill_2
XFILLER_19_843 VPWR VGND sg13g2_decap_8
XFILLER_46_695 VPWR VGND sg13g2_decap_8
XFILLER_34_857 VPWR VGND sg13g2_decap_8
XFILLER_21_529 VPWR VGND sg13g2_decap_8
X_3711_ _1193_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] net578 _0111_
+ VPWR VGND sg13g2_mux2_1
X_3642_ _1138_ net678 VPWR VGND net685 sg13g2_nand2b_2
X_3573_ _1074_ VPWR _0082_ VGND _1082_ _1084_ sg13g2_o21ai_1
XFILLER_46_0 VPWR VGND sg13g2_fill_1
X_2524_ _1936_ net735 _1565_ VPWR VGND sg13g2_nand2_1
X_2455_ _1873_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] net638
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] VPWR VGND sg13g2_a22oi_1
Xhold19 u_ser.shadow_reg\[7\] VPWR VGND net68 sg13g2_dlygate4sd3_1
X_2386_ _1766_ _1783_ _1798_ _1806_ VPWR VGND sg13g2_nor3_2
X_4125_ net826 VGND VPWR _0089_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_629 VPWR VGND sg13g2_decap_8
X_4056_ net836 VGND VPWR _0024_ u_ser.shadow_reg\[7\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
X_3007_ VGND VPWR _0510_ _0524_ _0561_ _0509_ sg13g2_a21oi_1
XFILLER_25_813 VPWR VGND sg13g2_decap_8
XFILLER_37_695 VPWR VGND sg13g2_decap_8
XFILLER_12_518 VPWR VGND sg13g2_decap_8
XFILLER_40_849 VPWR VGND sg13g2_decap_8
X_3909_ _0154_ VPWR _1340_ VGND sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[2\]
+ _1312_ sg13g2_o21ai_1
XFILLER_20_584 VPWR VGND sg13g2_decap_8
XFILLER_10_10 VPWR VGND sg13g2_fill_1
XFILLER_4_739 VPWR VGND sg13g2_decap_8
XFILLER_10_76 VPWR VGND sg13g2_fill_1
XFILLER_0_934 VPWR VGND sg13g2_decap_8
XFILLER_48_927 VPWR VGND sg13g2_decap_8
XFILLER_19_41 VPWR VGND sg13g2_fill_1
XFILLER_47_459 VPWR VGND sg13g2_decap_8
XFILLER_28_651 VPWR VGND sg13g2_decap_8
XFILLER_16_857 VPWR VGND sg13g2_decap_8
XFILLER_43_665 VPWR VGND sg13g2_decap_8
XFILLER_11_573 VPWR VGND sg13g2_decap_8
XFILLER_7_544 VPWR VGND sg13g2_decap_8
XFILLER_3_750 VPWR VGND sg13g2_decap_8
X_2240_ net742 _1617_ _1660_ VPWR VGND sg13g2_nor2_1
X_2171_ net768 net780 net770 _1591_ VPWR VGND sg13g2_or3_1
XFILLER_19_640 VPWR VGND sg13g2_decap_8
XFILLER_20_1011 VPWR VGND sg13g2_decap_8
XFILLER_38_459 VPWR VGND sg13g2_fill_1
XFILLER_25_109 VPWR VGND sg13g2_fill_1
XFILLER_46_492 VPWR VGND sg13g2_decap_8
XFILLER_34_654 VPWR VGND sg13g2_decap_8
X_3625_ _1127_ VPWR _0091_ VGND _1465_ _1122_ sg13g2_o21ai_1
X_3556_ net34 _1068_ _1069_ VPWR VGND sg13g2_nor2_2
X_2507_ _1921_ net5 _1858_ VPWR VGND sg13g2_nand2_1
X_3487_ _1009_ _0733_ _0804_ VPWR VGND sg13g2_xnor2_1
X_2438_ _1533_ VPWR _1858_ VGND _1842_ _1857_ sg13g2_o21ai_1
X_2369_ net743 _1676_ net786 _1789_ VPWR VGND _1788_ sg13g2_nand4_1
XFILLER_29_415 VPWR VGND sg13g2_fill_2
X_4108_ net824 VGND VPWR _0072_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[6\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
XFILLER_44_407 VPWR VGND sg13g2_decap_8
XFILLER_25_610 VPWR VGND sg13g2_decap_8
XFILLER_38_982 VPWR VGND sg13g2_decap_8
XFILLER_37_492 VPWR VGND sg13g2_decap_8
XFILLER_13_816 VPWR VGND sg13g2_decap_8
XFILLER_25_687 VPWR VGND sg13g2_decap_8
XFILLER_40_646 VPWR VGND sg13g2_decap_8
XFILLER_12_348 VPWR VGND sg13g2_fill_2
XFILLER_21_893 VPWR VGND sg13g2_decap_8
XFILLER_4_536 VPWR VGND sg13g2_decap_8
XFILLER_0_731 VPWR VGND sg13g2_decap_8
XFILLER_43_1022 VPWR VGND sg13g2_decap_8
XFILLER_48_724 VPWR VGND sg13g2_decap_8
XFILLER_29_993 VPWR VGND sg13g2_decap_8
XFILLER_44_974 VPWR VGND sg13g2_decap_8
XFILLER_43_462 VPWR VGND sg13g2_decap_8
XFILLER_16_654 VPWR VGND sg13g2_decap_8
XFILLER_31_668 VPWR VGND sg13g2_decap_8
XFILLER_8_831 VPWR VGND sg13g2_decap_8
XFILLER_12_882 VPWR VGND sg13g2_decap_8
X_3410_ VGND VPWR _0935_ _0934_ net598 sg13g2_or2_1
Xclkbuf_4_11_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_11_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3341_ _0869_ net597 net595 VPWR VGND sg13g2_nand2_2
X_3272_ _0775_ net588 _0800_ VPWR VGND sg13g2_and2_1
X_2223_ _1643_ net759 _1507_ VPWR VGND sg13g2_nand2_1
X_2154_ _1574_ net742 net732 VPWR VGND sg13g2_nand2_1
XFILLER_39_768 VPWR VGND sg13g2_decap_8
XFILLER_26_429 VPWR VGND sg13g2_decap_8
XFILLER_38_256 VPWR VGND sg13g2_fill_2
X_2085_ sap_3_inst.controller.stage\[3\] net759 _1505_ VPWR VGND sg13g2_nor2_2
XFILLER_35_941 VPWR VGND sg13g2_decap_8
XFILLER_22_657 VPWR VGND sg13g2_decap_8
X_2987_ _0541_ _0311_ net34 VPWR VGND sg13g2_nand2b_1
X_3608_ net605 _1008_ _1114_ VPWR VGND sg13g2_nor2_1
XFILLER_1_528 VPWR VGND sg13g2_decap_8
X_3539_ net584 _1054_ _1055_ _1056_ VPWR VGND sg13g2_nor3_1
XFILLER_44_204 VPWR VGND sg13g2_fill_2
XFILLER_44_215 VPWR VGND sg13g2_fill_1
XFILLER_13_613 VPWR VGND sg13g2_decap_8
XFILLER_25_484 VPWR VGND sg13g2_decap_8
XFILLER_26_996 VPWR VGND sg13g2_decap_8
XFILLER_41_966 VPWR VGND sg13g2_decap_8
XFILLER_12_178 VPWR VGND sg13g2_fill_2
XFILLER_21_690 VPWR VGND sg13g2_decap_8
XFILLER_5_812 VPWR VGND sg13g2_decap_8
XFILLER_5_889 VPWR VGND sg13g2_decap_8
XFILLER_48_521 VPWR VGND sg13g2_decap_8
XFILLER_48_598 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_3_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_29_790 VPWR VGND sg13g2_decap_8
XFILLER_36_738 VPWR VGND sg13g2_decap_8
XFILLER_17_963 VPWR VGND sg13g2_decap_8
XFILLER_44_771 VPWR VGND sg13g2_decap_8
X_2910_ _0467_ net682 net793 net683 net798 VPWR VGND sg13g2_a22oi_1
XFILLER_43_292 VPWR VGND sg13g2_fill_1
XFILLER_32_944 VPWR VGND sg13g2_decap_8
X_3890_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] _1322_
+ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] _1323_ _1308_ sg13g2_a221oi_1
X_2841_ _0370_ _0399_ _0400_ VPWR VGND sg13g2_nor2b_2
X_2772_ _0200_ _0330_ net625 _0333_ VPWR VGND sg13g2_nor3_1
X_3324_ VGND VPWR _1577_ net730 _0852_ _1620_ sg13g2_a21oi_1
Xfanout629 _1837_ net629 VPWR VGND sg13g2_buf_8
Xfanout618 net620 net618 VPWR VGND sg13g2_buf_8
Xfanout607 _0828_ net607 VPWR VGND sg13g2_buf_8
X_3255_ net704 net698 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] _0783_
+ VPWR VGND net695 sg13g2_nand4_1
X_2206_ _1626_ _1579_ _1623_ VPWR VGND sg13g2_nand2_1
X_3186_ _0714_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] net663 VPWR
+ VGND sg13g2_nand2_1
XFILLER_2_1008 VPWR VGND sg13g2_decap_8
XFILLER_39_565 VPWR VGND sg13g2_decap_8
X_2137_ sap_3_inst.controller.stage\[3\] net759 _1557_ VPWR VGND sg13g2_nor2b_2
XFILLER_27_749 VPWR VGND sg13g2_decap_8
X_2068_ VPWR _1490_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_41_207 VPWR VGND sg13g2_fill_2
XFILLER_23_911 VPWR VGND sg13g2_decap_8
XFILLER_10_627 VPWR VGND sg13g2_decap_8
XFILLER_22_454 VPWR VGND sg13g2_decap_8
XFILLER_23_988 VPWR VGND sg13g2_decap_8
XFILLER_5_108 VPWR VGND sg13g2_fill_1
XFILLER_2_826 VPWR VGND sg13g2_decap_8
XFILLER_40_1003 VPWR VGND sg13g2_decap_8
XFILLER_18_749 VPWR VGND sg13g2_decap_8
XFILLER_45_557 VPWR VGND sg13g2_decap_8
XFILLER_14_933 VPWR VGND sg13g2_decap_8
XFILLER_26_793 VPWR VGND sg13g2_decap_8
XFILLER_41_763 VPWR VGND sg13g2_decap_8
XFILLER_9_458 VPWR VGND sg13g2_fill_2
XFILLER_5_686 VPWR VGND sg13g2_decap_8
XFILLER_4_152 VPWR VGND sg13g2_fill_1
XFILLER_4_34 VPWR VGND sg13g2_decap_4
XFILLER_49_841 VPWR VGND sg13g2_decap_8
XFILLER_1_892 VPWR VGND sg13g2_decap_8
X_3040_ VGND VPWR sap_3_inst.alu.flags\[1\] _1956_ _0585_ _0584_ sg13g2_a21oi_1
XFILLER_48_395 VPWR VGND sg13g2_decap_8
XFILLER_36_535 VPWR VGND sg13g2_decap_8
XFILLER_17_760 VPWR VGND sg13g2_decap_8
X_3942_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\] net810
+ _1369_ net807 sg13g2_a21oi_1
XFILLER_17_1005 VPWR VGND sg13g2_decap_8
XFILLER_32_741 VPWR VGND sg13g2_decap_8
X_3873_ _1298_ _1305_ _1306_ VPWR VGND sg13g2_nor2_2
X_2824_ VGND VPWR _0383_ sap_3_inst.alu.tmp\[2\] net802 sg13g2_or2_1
XFILLER_20_969 VPWR VGND sg13g2_decap_8
X_2755_ _1951_ _1958_ _0316_ VPWR VGND sg13g2_nor2_1
X_2686_ VGND VPWR net749 _0268_ _0269_ _0266_ sg13g2_a21oi_1
X_3307_ VGND VPWR _0835_ net589 _0775_ sg13g2_or2_1
X_3238_ _0761_ _0762_ _0764_ _0765_ _0766_ VPWR VGND sg13g2_and4_1
X_3169_ _0697_ net703 net701 net692 VPWR VGND sg13g2_and3_2
XFILLER_27_546 VPWR VGND sg13g2_decap_8
XFILLER_42_527 VPWR VGND sg13g2_decap_8
XFILLER_23_785 VPWR VGND sg13g2_decap_8
Xfanout33 net23 net33 VPWR VGND sg13g2_buf_2
XFILLER_11_958 VPWR VGND sg13g2_decap_8
XFILLER_7_929 VPWR VGND sg13g2_decap_8
XFILLER_13_43 VPWR VGND sg13g2_fill_1
XFILLER_2_623 VPWR VGND sg13g2_decap_8
XFILLER_49_104 VPWR VGND sg13g2_fill_1
XFILLER_46_800 VPWR VGND sg13g2_decap_8
XFILLER_46_877 VPWR VGND sg13g2_decap_8
XFILLER_45_354 VPWR VGND sg13g2_decap_8
XFILLER_18_546 VPWR VGND sg13g2_decap_8
XFILLER_14_730 VPWR VGND sg13g2_decap_8
XFILLER_26_590 VPWR VGND sg13g2_decap_8
XFILLER_41_560 VPWR VGND sg13g2_decap_8
XFILLER_13_295 VPWR VGND sg13g2_fill_1
Xclkload14 VPWR clkload14/Y clknet_5_17__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
XFILLER_10_991 VPWR VGND sg13g2_decap_8
X_2540_ _1441_ _1948_ _1952_ VPWR VGND sg13g2_nor2_1
XFILLER_5_483 VPWR VGND sg13g2_decap_8
X_2471_ net576 VPWR _1889_ VGND _1884_ _1888_ sg13g2_o21ai_1
X_4210_ net828 VGND VPWR _0174_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\]
+ clknet_5_14__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4141_ net826 VGND VPWR _0105_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\]
+ clknet_5_11__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4072_ net838 VGND VPWR _0036_ sap_3_inst.alu.acc\[3\] clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_37_800 VPWR VGND sg13g2_decap_8
X_3023_ _0572_ VPWR _0044_ VGND _1445_ net717 sg13g2_o21ai_1
XFILLER_37_877 VPWR VGND sg13g2_decap_8
XFILLER_24_538 VPWR VGND sg13g2_decap_8
X_3925_ _1354_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] _1310_
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] VPWR VGND sg13g2_a22oi_1
Xclkload8 clknet_1_1__leaf_sap_3_inst.alu.clk clkload8/X VPWR VGND sg13g2_buf_8
XFILLER_20_766 VPWR VGND sg13g2_decap_8
X_3856_ net817 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\] _1290_ VPWR
+ VGND sg13g2_nor2b_1
X_3787_ _0136_ _1110_ _1244_ net612 _1487_ VPWR VGND sg13g2_a22oi_1
X_2807_ VGND VPWR net805 _0365_ _0367_ _0366_ sg13g2_a21oi_1
XFILLER_30_1024 VPWR VGND sg13g2_decap_4
X_2738_ net68 sap_3_inst.out\[7\] _0185_ _0024_ VPWR VGND sg13g2_mux2_1
X_2669_ sap_3_inst.alu.act\[5\] sap_3_inst.alu.act\[4\] sap_3_inst.alu.act\[7\] sap_3_inst.alu.act\[6\]
+ _0255_ VPWR VGND sg13g2_nor4_1
XFILLER_28_833 VPWR VGND sg13g2_decap_8
XFILLER_27_321 VPWR VGND sg13g2_fill_1
XFILLER_39_192 VPWR VGND sg13g2_fill_1
XFILLER_43_847 VPWR VGND sg13g2_decap_8
XFILLER_23_582 VPWR VGND sg13g2_decap_8
XFILLER_11_755 VPWR VGND sg13g2_decap_8
XFILLER_7_726 VPWR VGND sg13g2_decap_8
XFILLER_3_932 VPWR VGND sg13g2_decap_8
XFILLER_2_497 VPWR VGND sg13g2_decap_8
Xfanout790 net792 net790 VPWR VGND sg13g2_buf_8
XFILLER_19_822 VPWR VGND sg13g2_decap_8
XFILLER_46_674 VPWR VGND sg13g2_decap_8
XFILLER_19_899 VPWR VGND sg13g2_decap_8
XFILLER_33_302 VPWR VGND sg13g2_fill_1
XFILLER_34_836 VPWR VGND sg13g2_decap_8
XFILLER_21_508 VPWR VGND sg13g2_decap_8
XFILLER_42_891 VPWR VGND sg13g2_decap_8
X_3710_ VGND VPWR net711 _0990_ _1193_ _1192_ sg13g2_a21oi_1
X_3641_ net623 net684 _1137_ VPWR VGND sg13g2_nor2_2
X_3572_ _1084_ _0695_ _1083_ VPWR VGND sg13g2_nand2b_1
X_2523_ net771 _1934_ _1935_ VPWR VGND sg13g2_nor2_2
X_2454_ _1872_ net637 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] net647
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2385_ VPWR _1805_ net642 VGND sg13g2_inv_1
X_4124_ net825 VGND VPWR _0088_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_608 VPWR VGND sg13g2_decap_8
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
X_4055_ net836 VGND VPWR _0023_ u_ser.shadow_reg\[6\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
X_3006_ net575 _0554_ _0558_ _0559_ _0560_ VPWR VGND sg13g2_nor4_1
XFILLER_37_674 VPWR VGND sg13g2_decap_8
XFILLER_25_869 VPWR VGND sg13g2_decap_8
Xclkbuf_5_25__f_sap_3_inst.alu.clk_regs clknet_4_12_0_sap_3_inst.alu.clk_regs clknet_5_25__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_40_828 VPWR VGND sg13g2_decap_8
X_3908_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] _1338_
+ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] _1339_ _1308_ sg13g2_a221oi_1
XFILLER_20_563 VPWR VGND sg13g2_decap_8
X_3839_ sap_3_inst.reg_file.array_serializer_inst.state\[0\] sap_3_inst.reg_file.array_serializer_inst.state\[1\]
+ _1278_ VPWR VGND sg13g2_nor2b_2
XFILLER_4_718 VPWR VGND sg13g2_decap_8
XFILLER_10_66 VPWR VGND sg13g2_fill_1
XFILLER_0_913 VPWR VGND sg13g2_decap_8
XFILLER_48_906 VPWR VGND sg13g2_decap_8
XFILLER_47_438 VPWR VGND sg13g2_decap_8
XFILLER_19_118 VPWR VGND sg13g2_fill_2
XFILLER_28_630 VPWR VGND sg13g2_decap_8
XFILLER_43_644 VPWR VGND sg13g2_decap_8
XFILLER_16_836 VPWR VGND sg13g2_decap_8
XFILLER_7_523 VPWR VGND sg13g2_decap_8
XFILLER_11_552 VPWR VGND sg13g2_decap_8
X_2170_ net768 sap_3_inst.controller.opcode\[2\] net771 _1590_ VPWR VGND sg13g2_nor3_2
XFILLER_46_471 VPWR VGND sg13g2_decap_8
XFILLER_19_696 VPWR VGND sg13g2_decap_8
XFILLER_34_633 VPWR VGND sg13g2_decap_8
XFILLER_21_305 VPWR VGND sg13g2_fill_2
XFILLER_22_839 VPWR VGND sg13g2_decap_8
X_3624_ _1125_ _1126_ _1122_ _1127_ VPWR VGND sg13g2_nand3_1
X_3555_ _0829_ _1032_ _1068_ VPWR VGND sg13g2_nor2_1
X_2506_ _1920_ _1919_ _1723_ VPWR VGND sg13g2_nand2b_1
X_3486_ _1007_ _0992_ _1008_ VPWR VGND sg13g2_xor2_1
X_2437_ _1516_ _1855_ _1856_ _1857_ VPWR VGND sg13g2_nor3_1
X_2368_ _1788_ _1515_ _1787_ VPWR VGND sg13g2_nand2_1
X_2299_ _1719_ _1710_ _1713_ _1718_ VPWR VGND sg13g2_and3_1
X_4107_ net823 VGND VPWR _0071_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[5\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_38_961 VPWR VGND sg13g2_decap_8
XFILLER_24_110 VPWR VGND sg13g2_fill_1
XFILLER_25_666 VPWR VGND sg13g2_decap_8
XFILLER_40_625 VPWR VGND sg13g2_decap_8
XFILLER_21_872 VPWR VGND sg13g2_decap_8
XFILLER_4_515 VPWR VGND sg13g2_decap_8
XFILLER_0_710 VPWR VGND sg13g2_decap_8
XFILLER_48_703 VPWR VGND sg13g2_decap_8
XFILLER_43_1001 VPWR VGND sg13g2_decap_8
XFILLER_0_787 VPWR VGND sg13g2_decap_8
XFILLER_29_972 VPWR VGND sg13g2_decap_8
XFILLER_16_633 VPWR VGND sg13g2_decap_8
XFILLER_44_953 VPWR VGND sg13g2_decap_8
XFILLER_43_441 VPWR VGND sg13g2_decap_8
XFILLER_31_647 VPWR VGND sg13g2_decap_8
XFILLER_8_810 VPWR VGND sg13g2_decap_8
XFILLER_12_861 VPWR VGND sg13g2_decap_8
XFILLER_8_887 VPWR VGND sg13g2_decap_8
X_3340_ _0868_ net673 net684 VPWR VGND sg13g2_nand2b_1
X_3271_ _0791_ _0796_ _0797_ _0798_ _0799_ VPWR VGND sg13g2_and4_1
X_2222_ sap_3_inst.controller.stage\[3\] net759 _1642_ VPWR VGND sg13g2_and2_1
X_2153_ _1573_ _1534_ net754 _1507_ _1505_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_747 VPWR VGND sg13g2_decap_8
XFILLER_26_408 VPWR VGND sg13g2_decap_8
X_2084_ VGND VPWR _1504_ net761 net760 sg13g2_or2_1
XFILLER_35_920 VPWR VGND sg13g2_decap_8
XFILLER_35_997 VPWR VGND sg13g2_decap_8
XFILLER_10_809 VPWR VGND sg13g2_decap_8
XFILLER_22_636 VPWR VGND sg13g2_decap_8
X_2986_ _0540_ net788 net581 VPWR VGND sg13g2_nand2_1
X_3607_ _1113_ _0840_ _1112_ VPWR VGND sg13g2_nand2_1
XFILLER_1_507 VPWR VGND sg13g2_decap_8
X_3538_ net598 _0946_ _1055_ VPWR VGND sg13g2_nor2_1
X_3469_ _0885_ _0907_ _0931_ _0991_ _0992_ VPWR VGND sg13g2_and4_1
XFILLER_45_739 VPWR VGND sg13g2_decap_8
XFILLER_44_238 VPWR VGND sg13g2_fill_2
XFILLER_26_975 VPWR VGND sg13g2_decap_8
XFILLER_37_290 VPWR VGND sg13g2_fill_2
XFILLER_25_463 VPWR VGND sg13g2_decap_8
XFILLER_41_945 VPWR VGND sg13g2_decap_8
XFILLER_13_669 VPWR VGND sg13g2_decap_8
XFILLER_40_499 VPWR VGND sg13g2_decap_8
XFILLER_5_868 VPWR VGND sg13g2_decap_8
XFILLER_48_500 VPWR VGND sg13g2_decap_8
XFILLER_0_584 VPWR VGND sg13g2_decap_8
XFILLER_48_577 VPWR VGND sg13g2_decap_8
XFILLER_36_717 VPWR VGND sg13g2_decap_8
XFILLER_44_750 VPWR VGND sg13g2_decap_8
XFILLER_17_942 VPWR VGND sg13g2_decap_8
XFILLER_31_411 VPWR VGND sg13g2_decap_4
XFILLER_32_923 VPWR VGND sg13g2_decap_8
X_2840_ _0398_ _0384_ _0399_ VPWR VGND sg13g2_xor2_1
X_2771_ _0201_ _0331_ _0332_ VPWR VGND sg13g2_nor2_2
XFILLER_8_684 VPWR VGND sg13g2_decap_8
Xfanout619 net620 net619 VPWR VGND sg13g2_buf_2
X_3323_ net729 _1716_ _1516_ _0851_ VPWR VGND sg13g2_nand3_1
Xfanout608 _0705_ net608 VPWR VGND sg13g2_buf_8
XFILLER_21_0 VPWR VGND sg13g2_fill_2
X_3254_ net698 net695 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] _0782_
+ VPWR VGND net686 sg13g2_nand4_1
X_2205_ _1625_ _1579_ _1607_ _1622_ VPWR VGND sg13g2_and3_1
XFILLER_39_544 VPWR VGND sg13g2_decap_8
X_3185_ _0713_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] net675 VPWR
+ VGND sg13g2_nand2_1
X_2136_ _1551_ _1555_ _1556_ VPWR VGND sg13g2_nor2_2
XFILLER_26_227 VPWR VGND sg13g2_fill_2
XFILLER_27_728 VPWR VGND sg13g2_decap_8
X_2067_ VPWR _1489_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_42_709 VPWR VGND sg13g2_decap_8
XFILLER_23_967 VPWR VGND sg13g2_decap_8
XFILLER_35_794 VPWR VGND sg13g2_decap_8
XFILLER_10_606 VPWR VGND sg13g2_decap_8
X_2969_ _0482_ VPWR _0524_ VGND _0483_ _0486_ sg13g2_o21ai_1
XFILLER_33_1022 VPWR VGND sg13g2_decap_8
XFILLER_2_805 VPWR VGND sg13g2_decap_8
XFILLER_45_536 VPWR VGND sg13g2_decap_8
XFILLER_18_728 VPWR VGND sg13g2_decap_8
XFILLER_14_912 VPWR VGND sg13g2_decap_8
XFILLER_25_260 VPWR VGND sg13g2_decap_4
XFILLER_26_772 VPWR VGND sg13g2_decap_8
XFILLER_32_208 VPWR VGND sg13g2_fill_2
XFILLER_41_742 VPWR VGND sg13g2_decap_8
XFILLER_13_466 VPWR VGND sg13g2_fill_2
XFILLER_13_477 VPWR VGND sg13g2_fill_1
XFILLER_14_989 VPWR VGND sg13g2_decap_8
XFILLER_40_274 VPWR VGND sg13g2_fill_2
XFILLER_5_665 VPWR VGND sg13g2_decap_8
XFILLER_4_175 VPWR VGND sg13g2_fill_2
XFILLER_4_57 VPWR VGND sg13g2_fill_1
XFILLER_1_871 VPWR VGND sg13g2_decap_8
XFILLER_49_820 VPWR VGND sg13g2_decap_8
XFILLER_0_381 VPWR VGND sg13g2_fill_1
XFILLER_49_897 VPWR VGND sg13g2_decap_8
XFILLER_48_374 VPWR VGND sg13g2_decap_8
XFILLER_36_514 VPWR VGND sg13g2_decap_8
X_3941_ _1368_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] _1307_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_32_720 VPWR VGND sg13g2_decap_8
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
X_3872_ _1305_ sap_3_inst.reg_file.array_serializer_inst.word_index\[1\] VPWR VGND
+ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\] sg13g2_nand2b_2
X_2823_ net802 sap_3_inst.alu.tmp\[2\] _0382_ VPWR VGND sg13g2_and2_1
XFILLER_20_948 VPWR VGND sg13g2_decap_8
XFILLER_32_797 VPWR VGND sg13g2_decap_8
X_2754_ _0315_ _1945_ net708 VPWR VGND sg13g2_nand2b_1
XFILLER_8_481 VPWR VGND sg13g2_decap_8
X_2685_ _0268_ net719 _1704_ VPWR VGND sg13g2_nand2b_1
X_3306_ _0834_ net651 net712 VPWR VGND sg13g2_nand2_2
X_3237_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] _0759_
+ net657 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\] _0765_ net661 sg13g2_a221oi_1
X_3168_ _0696_ net687 _0694_ VPWR VGND sg13g2_nand2_1
XFILLER_27_525 VPWR VGND sg13g2_decap_8
X_2119_ _1539_ net740 _1520_ VPWR VGND sg13g2_nand2_1
XFILLER_42_506 VPWR VGND sg13g2_decap_8
X_3099_ _0627_ _1577_ _1654_ VPWR VGND sg13g2_nand2_1
XFILLER_35_591 VPWR VGND sg13g2_decap_8
Xfanout34 net24 net34 VPWR VGND sg13g2_buf_2
XFILLER_23_764 VPWR VGND sg13g2_decap_8
XFILLER_7_908 VPWR VGND sg13g2_decap_8
XFILLER_11_937 VPWR VGND sg13g2_decap_8
XFILLER_2_602 VPWR VGND sg13g2_decap_8
XFILLER_2_679 VPWR VGND sg13g2_decap_8
XFILLER_18_525 VPWR VGND sg13g2_decap_8
XFILLER_46_856 VPWR VGND sg13g2_decap_8
XFILLER_33_539 VPWR VGND sg13g2_decap_8
XFILLER_14_786 VPWR VGND sg13g2_decap_8
XFILLER_10_970 VPWR VGND sg13g2_decap_8
Xclkload15 clknet_5_19__leaf_sap_3_inst.alu.clk_regs clkload15/X VPWR VGND sg13g2_buf_1
X_2470_ _1886_ _1887_ _1885_ _1888_ VPWR VGND sg13g2_nand3_1
XFILLER_6_985 VPWR VGND sg13g2_decap_8
X_4140_ net825 VGND VPWR _0104_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\]
+ clknet_5_10__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4071_ net833 VGND VPWR _0035_ sap_3_inst.alu.acc\[2\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_49_694 VPWR VGND sg13g2_decap_8
X_3022_ _0572_ sap_3_inst.out\[3\] net717 VPWR VGND sg13g2_nand2_1
XFILLER_37_856 VPWR VGND sg13g2_decap_8
XFILLER_24_517 VPWR VGND sg13g2_decap_8
X_3924_ _1353_ _1314_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] _1300_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_32_594 VPWR VGND sg13g2_decap_8
XFILLER_20_745 VPWR VGND sg13g2_decap_8
Xclkload9 VPWR clkload9/Y clknet_5_1__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_3855_ _1288_ VPWR _1289_ VGND net817 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[1\]
+ sg13g2_o21ai_1
X_3786_ net15 net611 _1243_ _1244_ VPWR VGND sg13g2_nor3_1
X_2806_ net714 VPWR _0366_ VGND net805 _0365_ sg13g2_o21ai_1
XFILLER_30_1003 VPWR VGND sg13g2_decap_8
X_2737_ net65 sap_3_inst.out\[6\] _0185_ _0023_ VPWR VGND sg13g2_mux2_1
X_2668_ sap_3_inst.alu.act\[1\] sap_3_inst.alu.act\[0\] sap_3_inst.alu.act\[3\] sap_3_inst.alu.act\[2\]
+ _0254_ VPWR VGND sg13g2_nor4_1
X_2599_ VPWR _2008_ net19 VGND sg13g2_inv_1
XFILLER_27_300 VPWR VGND sg13g2_fill_2
XFILLER_28_812 VPWR VGND sg13g2_decap_8
XFILLER_43_826 VPWR VGND sg13g2_decap_8
XFILLER_28_889 VPWR VGND sg13g2_decap_8
XFILLER_15_539 VPWR VGND sg13g2_decap_8
XFILLER_11_734 VPWR VGND sg13g2_decap_8
XFILLER_23_561 VPWR VGND sg13g2_decap_8
XFILLER_7_705 VPWR VGND sg13g2_decap_8
XFILLER_10_255 VPWR VGND sg13g2_fill_1
XFILLER_3_911 VPWR VGND sg13g2_decap_8
XFILLER_46_1010 VPWR VGND sg13g2_decap_8
XFILLER_3_988 VPWR VGND sg13g2_decap_8
XFILLER_2_476 VPWR VGND sg13g2_decap_8
Xfanout780 net781 net780 VPWR VGND sg13g2_buf_8
Xfanout791 net792 net791 VPWR VGND sg13g2_buf_1
XFILLER_19_801 VPWR VGND sg13g2_decap_8
XFILLER_46_653 VPWR VGND sg13g2_decap_8
XFILLER_1_69 VPWR VGND sg13g2_fill_1
XFILLER_19_878 VPWR VGND sg13g2_decap_8
XFILLER_34_815 VPWR VGND sg13g2_decap_8
XFILLER_42_870 VPWR VGND sg13g2_decap_8
XFILLER_14_583 VPWR VGND sg13g2_decap_8
XFILLER_41_391 VPWR VGND sg13g2_fill_2
XFILLER_41_380 VPWR VGND sg13g2_fill_1
X_3640_ _1136_ net678 _1083_ VPWR VGND sg13g2_nand2b_1
X_3571_ net603 _0847_ _1083_ VPWR VGND sg13g2_and2_1
XFILLER_6_782 VPWR VGND sg13g2_decap_8
X_2522_ _1934_ net729 net769 _1675_ net745 VPWR VGND sg13g2_a22oi_1
X_2453_ _1871_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] net722
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2384_ _1739_ _1784_ _1799_ _1804_ VPWR VGND sg13g2_nor3_2
X_4123_ net824 VGND VPWR _0087_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\]
+ clknet_5_10__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4054_ net836 VGND VPWR _0022_ u_ser.shadow_reg\[5\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
XFILLER_49_491 VPWR VGND sg13g2_decap_8
X_3005_ _0556_ VPWR _0559_ VGND _0336_ _0549_ sg13g2_o21ai_1
XFILLER_37_653 VPWR VGND sg13g2_decap_8
XFILLER_25_848 VPWR VGND sg13g2_decap_8
XFILLER_40_807 VPWR VGND sg13g2_decap_8
XFILLER_20_542 VPWR VGND sg13g2_decap_8
X_3907_ _1335_ _1336_ _1334_ _1338_ VPWR VGND _1337_ sg13g2_nand4_1
X_3838_ _0154_ net811 VPWR VGND sg13g2_inv_2
X_3769_ _1224_ VPWR _0132_ VGND _1225_ _1230_ sg13g2_o21ai_1
XFILLER_0_969 VPWR VGND sg13g2_decap_8
XFILLER_47_417 VPWR VGND sg13g2_decap_8
XFILLER_16_815 VPWR VGND sg13g2_decap_8
XFILLER_43_623 VPWR VGND sg13g2_decap_8
XFILLER_28_686 VPWR VGND sg13g2_decap_8
XFILLER_35_42 VPWR VGND sg13g2_fill_2
XFILLER_27_196 VPWR VGND sg13g2_fill_1
XFILLER_24_881 VPWR VGND sg13g2_decap_8
XFILLER_31_829 VPWR VGND sg13g2_decap_8
XFILLER_11_531 VPWR VGND sg13g2_decap_8
XFILLER_7_502 VPWR VGND sg13g2_decap_8
XFILLER_7_579 VPWR VGND sg13g2_decap_8
XFILLER_3_785 VPWR VGND sg13g2_decap_8
XFILLER_2_273 VPWR VGND sg13g2_fill_1
XFILLER_39_929 VPWR VGND sg13g2_decap_8
XFILLER_47_984 VPWR VGND sg13g2_decap_8
XFILLER_46_450 VPWR VGND sg13g2_decap_8
XFILLER_19_675 VPWR VGND sg13g2_decap_8
XFILLER_33_100 VPWR VGND sg13g2_fill_1
XFILLER_34_612 VPWR VGND sg13g2_decap_8
XFILLER_18_196 VPWR VGND sg13g2_fill_1
XFILLER_22_818 VPWR VGND sg13g2_decap_8
XFILLER_34_689 VPWR VGND sg13g2_decap_8
XFILLER_30_884 VPWR VGND sg13g2_decap_8
X_3623_ _1126_ net600 _0898_ VPWR VGND sg13g2_nand2b_1
X_3554_ _0080_ _1064_ _1067_ net584 _1493_ VPWR VGND sg13g2_a22oi_1
X_3485_ _1006_ VPWR _1007_ VGND _1001_ _1005_ sg13g2_o21ai_1
X_2505_ _1919_ _1915_ _1918_ net649 _1474_ VPWR VGND sg13g2_a22oi_1
X_2436_ _1541_ _1678_ _1856_ VPWR VGND sg13g2_nor2_1
X_2367_ _1546_ _1565_ _1566_ _1787_ VGND VPWR _1786_ sg13g2_nor4_2
X_2298_ _1718_ _1556_ _1717_ VPWR VGND sg13g2_nand2b_1
X_4106_ net823 VGND VPWR _0070_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[4\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
XFILLER_38_940 VPWR VGND sg13g2_decap_8
X_4037_ _0195_ _1439_ _1436_ net61 _1437_ VPWR VGND sg13g2_a22oi_1
XFILLER_37_450 VPWR VGND sg13g2_fill_1
XFILLER_25_645 VPWR VGND sg13g2_decap_8
XFILLER_40_604 VPWR VGND sg13g2_decap_8
XFILLER_21_851 VPWR VGND sg13g2_decap_8
XFILLER_0_766 VPWR VGND sg13g2_decap_8
XFILLER_48_759 VPWR VGND sg13g2_decap_8
XFILLER_47_247 VPWR VGND sg13g2_fill_2
XFILLER_29_951 VPWR VGND sg13g2_decap_8
XFILLER_44_932 VPWR VGND sg13g2_decap_8
XFILLER_16_612 VPWR VGND sg13g2_decap_8
XFILLER_28_483 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_decap_8
XFILLER_15_122 VPWR VGND sg13g2_fill_1
XFILLER_16_689 VPWR VGND sg13g2_decap_8
XFILLER_31_626 VPWR VGND sg13g2_decap_8
XFILLER_43_497 VPWR VGND sg13g2_decap_8
XFILLER_12_840 VPWR VGND sg13g2_decap_8
XFILLER_30_136 VPWR VGND sg13g2_fill_2
XFILLER_8_866 VPWR VGND sg13g2_decap_8
XFILLER_3_582 VPWR VGND sg13g2_decap_8
X_3270_ _0792_ _0793_ _0794_ _0795_ _0798_ VPWR VGND sg13g2_and4_1
X_2221_ _1613_ VPWR _1641_ VGND _1638_ _1640_ sg13g2_o21ai_1
XFILLER_39_726 VPWR VGND sg13g2_decap_8
X_2152_ _1572_ _1534_ net754 VPWR VGND sg13g2_nand2_1
X_2083_ net760 net761 _1503_ VPWR VGND sg13g2_nor2_2
XFILLER_47_781 VPWR VGND sg13g2_decap_8
XFILLER_35_976 VPWR VGND sg13g2_decap_8
XFILLER_22_615 VPWR VGND sg13g2_decap_8
XFILLER_34_486 VPWR VGND sg13g2_decap_8
X_2985_ net581 net791 _0539_ _0039_ VPWR VGND sg13g2_a21o_1
XFILLER_30_681 VPWR VGND sg13g2_decap_8
X_3606_ VGND VPWR _0732_ _0839_ _1112_ _0873_ sg13g2_a21oi_1
X_3537_ _0943_ _0828_ net20 _1054_ VPWR VGND sg13g2_a21o_1
XFILLER_27_1008 VPWR VGND sg13g2_decap_8
X_3468_ _0953_ _0977_ _0991_ VPWR VGND sg13g2_nor2_1
X_2419_ net763 _1575_ _1639_ _1839_ VPWR VGND sg13g2_nor3_2
X_3399_ _0924_ net666 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] net676
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_45_718 VPWR VGND sg13g2_decap_8
XFILLER_44_206 VPWR VGND sg13g2_fill_1
XFILLER_25_442 VPWR VGND sg13g2_decap_8
XFILLER_26_954 VPWR VGND sg13g2_decap_8
XFILLER_41_924 VPWR VGND sg13g2_decap_8
XFILLER_13_648 VPWR VGND sg13g2_decap_8
XFILLER_40_478 VPWR VGND sg13g2_decap_8
XFILLER_5_847 VPWR VGND sg13g2_decap_8
XFILLER_10_1012 VPWR VGND sg13g2_decap_8
XFILLER_0_563 VPWR VGND sg13g2_decap_8
XFILLER_48_556 VPWR VGND sg13g2_decap_8
XFILLER_17_921 VPWR VGND sg13g2_decap_8
XFILLER_16_420 VPWR VGND sg13g2_fill_1
XFILLER_17_998 VPWR VGND sg13g2_decap_8
XFILLER_32_902 VPWR VGND sg13g2_decap_8
XFILLER_16_486 VPWR VGND sg13g2_decap_8
XFILLER_32_979 VPWR VGND sg13g2_decap_8
X_2770_ _0331_ _1955_ _1957_ VPWR VGND sg13g2_nand2_2
XFILLER_8_663 VPWR VGND sg13g2_decap_8
XFILLER_7_195 VPWR VGND sg13g2_fill_1
X_3322_ _0850_ net653 net712 VPWR VGND sg13g2_nand2_2
Xfanout609 _0705_ net609 VPWR VGND sg13g2_buf_1
X_3253_ net702 net695 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] _0781_
+ VPWR VGND net689 sg13g2_nand4_1
X_3184_ _0712_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] net678 VPWR
+ VGND sg13g2_nand2_1
X_2204_ _1624_ _1607_ _1622_ VPWR VGND sg13g2_nand2_1
XFILLER_39_523 VPWR VGND sg13g2_decap_8
X_2135_ net767 _1554_ _1555_ VPWR VGND sg13g2_nor2_1
XFILLER_27_707 VPWR VGND sg13g2_decap_8
X_2066_ VPWR _1488_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_35_773 VPWR VGND sg13g2_decap_8
XFILLER_22_423 VPWR VGND sg13g2_decap_8
XFILLER_23_946 VPWR VGND sg13g2_decap_8
XFILLER_33_1001 VPWR VGND sg13g2_decap_8
X_2968_ _0518_ _0519_ _0520_ _0522_ _0523_ VPWR VGND sg13g2_and4_1
XFILLER_22_489 VPWR VGND sg13g2_decap_8
XFILLER_31_990 VPWR VGND sg13g2_decap_8
X_2899_ _0455_ VPWR _0456_ VGND net796 _0324_ sg13g2_o21ai_1
XFILLER_49_309 VPWR VGND sg13g2_decap_8
XFILLER_18_707 VPWR VGND sg13g2_decap_8
XFILLER_45_515 VPWR VGND sg13g2_decap_8
XFILLER_26_751 VPWR VGND sg13g2_decap_8
XFILLER_41_721 VPWR VGND sg13g2_decap_8
XFILLER_14_968 VPWR VGND sg13g2_decap_8
XFILLER_41_798 VPWR VGND sg13g2_decap_8
XFILLER_5_644 VPWR VGND sg13g2_decap_8
XFILLER_4_110 VPWR VGND sg13g2_fill_2
XFILLER_1_850 VPWR VGND sg13g2_decap_8
XFILLER_49_876 VPWR VGND sg13g2_decap_8
XFILLER_48_353 VPWR VGND sg13g2_decap_8
X_3940_ _1367_ _1309_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] _1301_
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_17_795 VPWR VGND sg13g2_decap_8
XFILLER_32_776 VPWR VGND sg13g2_decap_8
X_3871_ _1302_ _1303_ _1304_ VPWR VGND sg13g2_nor2_1
X_2822_ net580 net803 _0381_ _0034_ VPWR VGND sg13g2_a21o_1
XFILLER_20_927 VPWR VGND sg13g2_decap_8
X_2753_ _0313_ VPWR _0314_ VGND _1543_ net732 sg13g2_o21ai_1
XFILLER_9_994 VPWR VGND sg13g2_decap_8
X_2684_ _1528_ _1585_ net743 _0267_ VPWR VGND _1627_ sg13g2_nand4_1
X_3305_ net653 net711 _0833_ VPWR VGND sg13g2_nor2_1
X_3236_ _0757_ _0758_ _0760_ _0763_ _0764_ VPWR VGND sg13g2_and4_1
XFILLER_27_504 VPWR VGND sg13g2_decap_8
X_3167_ net705 net699 _0658_ _0695_ VGND VPWR net689 sg13g2_nor4_2
XFILLER_39_386 VPWR VGND sg13g2_fill_2
X_3098_ _0626_ _1702_ net731 _1619_ _1582_ VPWR VGND sg13g2_a22oi_1
X_2118_ VGND VPWR net740 _1516_ _1538_ _1537_ sg13g2_a21oi_1
X_2049_ VPWR _1471_ sap_3_inst.alu.tmp\[2\] VGND sg13g2_inv_1
XFILLER_35_570 VPWR VGND sg13g2_decap_8
XFILLER_11_916 VPWR VGND sg13g2_decap_8
XFILLER_23_743 VPWR VGND sg13g2_decap_8
XFILLER_2_658 VPWR VGND sg13g2_decap_8
XFILLER_1_179 VPWR VGND sg13g2_fill_1
XFILLER_46_835 VPWR VGND sg13g2_decap_8
XFILLER_18_504 VPWR VGND sg13g2_decap_8
XFILLER_33_518 VPWR VGND sg13g2_decap_8
XFILLER_45_389 VPWR VGND sg13g2_decap_8
XFILLER_14_765 VPWR VGND sg13g2_decap_8
XFILLER_41_595 VPWR VGND sg13g2_decap_8
Xclkload16 VPWR clkload16/Y clknet_5_21__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
XFILLER_6_964 VPWR VGND sg13g2_decap_8
X_4070_ net833 VGND VPWR _0034_ sap_3_inst.alu.acc\[1\] clknet_5_18__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_49_673 VPWR VGND sg13g2_decap_8
X_3021_ net801 sap_3_inst.out\[2\] net717 _0043_ VPWR VGND sg13g2_mux2_1
XFILLER_37_835 VPWR VGND sg13g2_decap_8
XFILLER_17_592 VPWR VGND sg13g2_decap_8
X_3923_ _1352_ _1307_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] _1306_
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_724 VPWR VGND sg13g2_decap_8
XFILLER_32_573 VPWR VGND sg13g2_decap_8
X_3854_ VGND VPWR net817 _1502_ _1288_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\]
+ sg13g2_a21oi_1
X_2805_ _0363_ _0364_ _0365_ VPWR VGND sg13g2_nor2b_1
X_3785_ VGND VPWR _0978_ _1007_ _1243_ _1242_ sg13g2_a21oi_1
X_2736_ net66 sap_3_inst.out\[5\] net813 _0022_ VPWR VGND sg13g2_mux2_1
XFILLER_9_791 VPWR VGND sg13g2_decap_8
X_2667_ _0251_ _0252_ _1960_ _0253_ VPWR VGND sg13g2_nand3_1
X_2598_ _1999_ _2007_ _1995_ net19 VPWR VGND sg13g2_nand3_1
XFILLER_8_1027 VPWR VGND sg13g2_fill_2
X_3219_ net698 net694 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] _0747_
+ VPWR VGND net686 sg13g2_nand4_1
X_4199_ net846 VGND VPWR _0163_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[2\]
+ clknet_3_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_28_868 VPWR VGND sg13g2_decap_8
XFILLER_43_805 VPWR VGND sg13g2_decap_8
XFILLER_15_518 VPWR VGND sg13g2_decap_8
XFILLER_23_540 VPWR VGND sg13g2_decap_8
XFILLER_24_33 VPWR VGND sg13g2_fill_2
XFILLER_11_713 VPWR VGND sg13g2_decap_8
XFILLER_3_967 VPWR VGND sg13g2_decap_8
XFILLER_49_52 VPWR VGND sg13g2_fill_1
Xfanout781 sap_3_inst.controller.opcode\[2\] net781 VPWR VGND sg13g2_buf_8
Xfanout770 sap_3_inst.controller.opcode\[6\] net770 VPWR VGND sg13g2_buf_8
Xfanout792 sap_3_inst.alu.acc\[6\] net792 VPWR VGND sg13g2_buf_8
XFILLER_46_632 VPWR VGND sg13g2_decap_8
XFILLER_19_857 VPWR VGND sg13g2_decap_8
XFILLER_14_562 VPWR VGND sg13g2_decap_8
X_3570_ VGND VPWR _1079_ _1081_ _1082_ _0874_ sg13g2_a21oi_1
X_2521_ net724 VPWR _1933_ VGND _1543_ net734 sg13g2_o21ai_1
XFILLER_6_761 VPWR VGND sg13g2_decap_8
X_2452_ _1870_ net640 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] net643
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2383_ _1738_ _1765_ _1784_ _1803_ VGND VPWR _1799_ sg13g2_nor4_2
X_4122_ net842 VGND VPWR _0086_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\]
+ clknet_5_30__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4053_ net836 VGND VPWR _0021_ u_ser.shadow_reg\[4\] clknet_3_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_49_470 VPWR VGND sg13g2_decap_8
X_3004_ _0557_ VPWR _0558_ VGND net787 _0324_ sg13g2_o21ai_1
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_37_632 VPWR VGND sg13g2_decap_8
XFILLER_36_131 VPWR VGND sg13g2_fill_1
XFILLER_25_827 VPWR VGND sg13g2_decap_8
X_3906_ _1337_ net809 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] _1300_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_882 VPWR VGND sg13g2_decap_8
XFILLER_20_521 VPWR VGND sg13g2_decap_8
X_3837_ VGND VPWR _1277_ sap_3_inst.reg_file.array_serializer_inst.state\[0\] sap_3_inst.reg_file.array_serializer_inst.state\[1\]
+ sg13g2_or2_1
XFILLER_20_598 VPWR VGND sg13g2_decap_8
X_3768_ VGND VPWR net606 _0921_ _1230_ _1229_ sg13g2_a21oi_1
X_2719_ _1589_ VPWR _0290_ VGND _1697_ _1725_ sg13g2_o21ai_1
X_3699_ _1183_ VPWR _1184_ VGND net654 _1182_ sg13g2_o21ai_1
XFILLER_10_57 VPWR VGND sg13g2_fill_2
XFILLER_0_948 VPWR VGND sg13g2_decap_8
XFILLER_43_602 VPWR VGND sg13g2_decap_8
XFILLER_28_665 VPWR VGND sg13g2_decap_8
XFILLER_42_112 VPWR VGND sg13g2_fill_2
XFILLER_31_808 VPWR VGND sg13g2_decap_8
XFILLER_35_54 VPWR VGND sg13g2_fill_2
XFILLER_43_679 VPWR VGND sg13g2_decap_8
XFILLER_24_860 VPWR VGND sg13g2_decap_8
XFILLER_11_510 VPWR VGND sg13g2_decap_8
XFILLER_30_329 VPWR VGND sg13g2_decap_4
XFILLER_7_558 VPWR VGND sg13g2_decap_8
XFILLER_11_587 VPWR VGND sg13g2_decap_8
XFILLER_3_764 VPWR VGND sg13g2_decap_8
XFILLER_39_908 VPWR VGND sg13g2_decap_8
XFILLER_47_963 VPWR VGND sg13g2_decap_8
XFILLER_19_654 VPWR VGND sg13g2_decap_8
XFILLER_20_1025 VPWR VGND sg13g2_decap_4
XFILLER_18_186 VPWR VGND sg13g2_fill_1
XFILLER_34_668 VPWR VGND sg13g2_decap_8
XFILLER_15_882 VPWR VGND sg13g2_decap_8
XFILLER_30_863 VPWR VGND sg13g2_decap_8
X_3622_ _1125_ _1051_ _1124_ VPWR VGND sg13g2_nand2_1
X_3553_ net584 _1066_ _1067_ VPWR VGND sg13g2_nor2_1
X_2504_ net648 _1913_ _1916_ _1917_ _1918_ VPWR VGND sg13g2_and4_1
X_3484_ _1006_ _1484_ net670 VPWR VGND sg13g2_nand2_1
X_2435_ VPWR VGND _1854_ net724 _1845_ net737 _1855_ _1780_ sg13g2_a221oi_1
XFILLER_5_1008 VPWR VGND sg13g2_decap_8
X_2366_ _1524_ _1676_ _1786_ VPWR VGND sg13g2_nor2_2
X_4105_ net823 VGND VPWR _0069_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[3\]
+ clknet_5_0__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
X_2297_ net741 _1715_ _1717_ VPWR VGND sg13g2_nor2_1
X_4036_ net814 _1415_ u_ser.bit_pos\[1\] _1436_ VPWR VGND sg13g2_nand3_1
XFILLER_25_624 VPWR VGND sg13g2_decap_8
XFILLER_38_996 VPWR VGND sg13g2_decap_8
XFILLER_21_830 VPWR VGND sg13g2_decap_8
XFILLER_0_745 VPWR VGND sg13g2_decap_8
XFILLER_48_738 VPWR VGND sg13g2_decap_8
XFILLER_29_930 VPWR VGND sg13g2_decap_8
XFILLER_44_911 VPWR VGND sg13g2_decap_8
XFILLER_28_462 VPWR VGND sg13g2_decap_8
XFILLER_16_668 VPWR VGND sg13g2_decap_8
XFILLER_44_988 VPWR VGND sg13g2_decap_8
XFILLER_43_476 VPWR VGND sg13g2_decap_8
XFILLER_31_605 VPWR VGND sg13g2_decap_8
XFILLER_8_845 VPWR VGND sg13g2_decap_8
XFILLER_12_896 VPWR VGND sg13g2_decap_8
XFILLER_3_561 VPWR VGND sg13g2_decap_8
X_2220_ _1640_ net732 _1630_ VPWR VGND sg13g2_nand2_1
XFILLER_39_705 VPWR VGND sg13g2_decap_8
X_2151_ _1534_ net754 _1571_ VPWR VGND sg13g2_and2_1
XFILLER_47_760 VPWR VGND sg13g2_decap_8
XFILLER_35_955 VPWR VGND sg13g2_decap_8
X_2984_ net581 _0507_ _0538_ _0539_ VPWR VGND sg13g2_nor3_1
XFILLER_30_660 VPWR VGND sg13g2_decap_8
X_3605_ net33 net15 _1075_ _1111_ VPWR VGND sg13g2_mux2_1
X_3536_ VGND VPWR _1457_ net585 _0076_ _1053_ sg13g2_a21oi_1
X_3467_ _0990_ _0988_ _0989_ _0987_ net653 VPWR VGND sg13g2_a22oi_1
X_2418_ net789 net628 _1838_ VPWR VGND sg13g2_nor2_1
X_3398_ _0923_ net661 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] net663
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2349_ VGND VPWR net740 net727 _1769_ _1603_ sg13g2_a21oi_1
XFILLER_29_226 VPWR VGND sg13g2_fill_1
XFILLER_29_237 VPWR VGND sg13g2_fill_1
X_4019_ _1423_ _1425_ _0186_ _1427_ VPWR VGND _1426_ sg13g2_nand4_1
XFILLER_26_933 VPWR VGND sg13g2_decap_8
XFILLER_38_793 VPWR VGND sg13g2_decap_8
XFILLER_25_421 VPWR VGND sg13g2_decap_8
XFILLER_37_281 VPWR VGND sg13g2_fill_1
XFILLER_41_903 VPWR VGND sg13g2_decap_8
XFILLER_13_627 VPWR VGND sg13g2_decap_8
XFILLER_25_498 VPWR VGND sg13g2_decap_8
XFILLER_9_609 VPWR VGND sg13g2_decap_8
XFILLER_40_457 VPWR VGND sg13g2_decap_8
XFILLER_5_826 VPWR VGND sg13g2_decap_8
XFILLER_4_358 VPWR VGND sg13g2_fill_1
XFILLER_0_542 VPWR VGND sg13g2_decap_8
XFILLER_48_535 VPWR VGND sg13g2_decap_8
XFILLER_17_900 VPWR VGND sg13g2_decap_8
XFILLER_44_785 VPWR VGND sg13g2_decap_8
XFILLER_17_977 VPWR VGND sg13g2_decap_8
XFILLER_32_958 VPWR VGND sg13g2_decap_8
XFILLER_8_642 VPWR VGND sg13g2_decap_8
XFILLER_12_693 VPWR VGND sg13g2_decap_8
XFILLER_7_152 VPWR VGND sg13g2_fill_2
X_3321_ net651 net711 _0849_ VPWR VGND sg13g2_nor2_2
X_3252_ net698 net694 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] _0780_
+ VPWR VGND net689 sg13g2_nand4_1
XFILLER_39_502 VPWR VGND sg13g2_decap_8
X_2203_ _1607_ _1622_ _1623_ VPWR VGND sg13g2_and2_1
X_3183_ _0711_ _0710_ VPWR VGND sg13g2_inv_2
X_2134_ _1554_ net745 _1546_ VPWR VGND sg13g2_nand2_1
XFILLER_39_579 VPWR VGND sg13g2_decap_8
X_2065_ VPWR _1487_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_26_229 VPWR VGND sg13g2_fill_1
XFILLER_23_925 VPWR VGND sg13g2_decap_8
XFILLER_35_752 VPWR VGND sg13g2_decap_8
XFILLER_22_468 VPWR VGND sg13g2_decap_8
X_2967_ _0522_ _0515_ _0521_ VPWR VGND sg13g2_nand2b_1
X_2898_ _0342_ VPWR _0455_ VGND net796 sap_3_inst.alu.tmp\[4\] sg13g2_o21ai_1
X_3519_ _1027_ _1013_ _1040_ VPWR VGND sg13g2_xor2_1
XFILLER_40_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_1017 VPWR VGND sg13g2_decap_8
XFILLER_26_730 VPWR VGND sg13g2_decap_8
XFILLER_38_590 VPWR VGND sg13g2_decap_8
XFILLER_41_700 VPWR VGND sg13g2_decap_8
XFILLER_14_947 VPWR VGND sg13g2_decap_8
XFILLER_41_777 VPWR VGND sg13g2_decap_8
XFILLER_13_435 VPWR VGND sg13g2_fill_2
XFILLER_13_468 VPWR VGND sg13g2_fill_1
XFILLER_5_623 VPWR VGND sg13g2_decap_8
XFILLER_49_855 VPWR VGND sg13g2_decap_8
XFILLER_48_332 VPWR VGND sg13g2_decap_8
XFILLER_1_1011 VPWR VGND sg13g2_decap_8
XFILLER_36_549 VPWR VGND sg13g2_decap_8
XFILLER_17_774 VPWR VGND sg13g2_decap_8
XFILLER_44_582 VPWR VGND sg13g2_decap_8
XFILLER_17_1019 VPWR VGND sg13g2_decap_8
XFILLER_20_906 VPWR VGND sg13g2_decap_8
XFILLER_32_755 VPWR VGND sg13g2_decap_8
X_3870_ _1303_ net816 VPWR VGND net815 sg13g2_nand2b_2
X_2821_ VPWR VGND _0380_ net580 _0379_ _0227_ _0381_ net626 sg13g2_a221oi_1
X_2752_ _0312_ VPWR _0313_ VGND net736 _1827_ sg13g2_o21ai_1
XFILLER_12_490 VPWR VGND sg13g2_decap_8
XFILLER_13_991 VPWR VGND sg13g2_decap_8
XFILLER_9_973 VPWR VGND sg13g2_decap_8
X_2683_ _0266_ _1787_ _1658_ VPWR VGND sg13g2_nand2b_1
X_3304_ _0822_ _0824_ _0816_ _0832_ VPWR VGND _0831_ sg13g2_nand4_1
X_3235_ net697 net691 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] _0763_
+ VPWR VGND net687 sg13g2_nand4_1
X_3166_ net700 net691 _0694_ VPWR VGND sg13g2_nor2_1
X_3097_ net731 _1598_ _0625_ VPWR VGND sg13g2_nor2_1
X_2117_ _1533_ _1535_ _1530_ _1537_ VPWR VGND sg13g2_nand3_1
X_2048_ VPWR _1470_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] VGND
+ sg13g2_inv_1
XFILLER_23_722 VPWR VGND sg13g2_decap_8
X_3999_ _1409_ VPWR _1410_ VGND net790 net710 sg13g2_o21ai_1
XFILLER_23_799 VPWR VGND sg13g2_decap_8
XFILLER_2_637 VPWR VGND sg13g2_decap_8
Xclkbuf_5_4__f_sap_3_inst.alu.clk_regs clknet_4_2_0_sap_3_inst.alu.clk_regs clknet_5_4__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_46_814 VPWR VGND sg13g2_decap_8
XFILLER_45_368 VPWR VGND sg13g2_decap_8
XFILLER_13_232 VPWR VGND sg13g2_fill_2
XFILLER_14_744 VPWR VGND sg13g2_decap_8
XFILLER_41_574 VPWR VGND sg13g2_decap_8
Xclkload17 clknet_5_23__leaf_sap_3_inst.alu.clk_regs clkload17/X VPWR VGND sg13g2_buf_1
XFILLER_6_943 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_4
XFILLER_5_497 VPWR VGND sg13g2_decap_8
XFILLER_49_652 VPWR VGND sg13g2_decap_8
XFILLER_23_1023 VPWR VGND sg13g2_decap_4
X_3020_ _0571_ VPWR _0042_ VGND _1458_ net717 sg13g2_o21ai_1
XFILLER_37_814 VPWR VGND sg13g2_decap_8
XFILLER_17_571 VPWR VGND sg13g2_decap_8
X_3922_ _1351_ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] _1304_
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_703 VPWR VGND sg13g2_decap_8
XFILLER_32_552 VPWR VGND sg13g2_decap_8
X_3853_ net71 _0155_ _1287_ VPWR VGND sg13g2_nor2_1
X_2804_ _1458_ VPWR _0364_ VGND _1550_ _1796_ sg13g2_o21ai_1
XFILLER_9_770 VPWR VGND sg13g2_decap_8
X_3784_ _0872_ VPWR _1242_ VGND _0978_ _1007_ sg13g2_o21ai_1
X_2735_ net67 sap_3_inst.out\[4\] net813 _0021_ VPWR VGND sg13g2_mux2_1
X_2666_ net800 net802 net803 net805 _0252_ VPWR VGND sg13g2_nor4_1
XFILLER_8_1006 VPWR VGND sg13g2_decap_8
X_2597_ net577 VPWR _2007_ VGND _2004_ _2006_ sg13g2_o21ai_1
Xclkbuf_5_11__f_sap_3_inst.alu.clk_regs clknet_4_5_0_sap_3_inst.alu.clk_regs clknet_5_11__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_27_302 VPWR VGND sg13g2_fill_1
X_4198_ net846 VGND VPWR _0162_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[1\]
+ clknet_3_3__leaf_clk sg13g2_dfrbpq_1
X_3218_ net704 net701 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] _0746_
+ VPWR VGND net694 sg13g2_nand4_1
X_3149_ _0677_ _1587_ _0676_ VPWR VGND sg13g2_nand2_1
XFILLER_28_847 VPWR VGND sg13g2_decap_8
XFILLER_42_327 VPWR VGND sg13g2_fill_1
XFILLER_23_596 VPWR VGND sg13g2_decap_8
XFILLER_11_769 VPWR VGND sg13g2_decap_8
XFILLER_3_946 VPWR VGND sg13g2_decap_8
Xfanout760 sap_3_inst.controller.stage\[1\] net760 VPWR VGND sg13g2_buf_8
Xfanout782 net784 net782 VPWR VGND sg13g2_buf_8
Xfanout793 net795 net793 VPWR VGND sg13g2_buf_8
Xfanout771 sap_3_inst.controller.opcode\[6\] net771 VPWR VGND sg13g2_buf_8
XFILLER_46_611 VPWR VGND sg13g2_decap_8
XFILLER_19_836 VPWR VGND sg13g2_decap_8
XFILLER_45_121 VPWR VGND sg13g2_fill_2
XFILLER_46_688 VPWR VGND sg13g2_decap_8
XFILLER_14_541 VPWR VGND sg13g2_decap_8
XFILLER_41_393 VPWR VGND sg13g2_fill_1
XFILLER_6_740 VPWR VGND sg13g2_decap_8
X_2520_ sap_3_inst.alu.flags\[4\] net32 _1867_ _0029_ VPWR VGND sg13g2_mux2_1
X_2451_ _1869_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] net645
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2382_ _1739_ _1784_ _1798_ _1802_ VPWR VGND sg13g2_nor3_2
X_4121_ net819 VGND VPWR _0085_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\]
+ clknet_5_5__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4052_ net832 VGND VPWR _0020_ u_ser.shadow_reg\[3\] clknet_3_1__leaf_clk sg13g2_dfrbpq_1
X_3003_ _0557_ _0547_ _0344_ _0546_ _0342_ VPWR VGND sg13g2_a22oi_1
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
XFILLER_37_611 VPWR VGND sg13g2_decap_8
XFILLER_25_806 VPWR VGND sg13g2_decap_8
XFILLER_37_688 VPWR VGND sg13g2_decap_8
XFILLER_20_500 VPWR VGND sg13g2_decap_8
X_3905_ _1336_ _1309_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] _1301_
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_861 VPWR VGND sg13g2_decap_8
X_3836_ _1272_ VPWR _0153_ VGND _1275_ _1276_ sg13g2_o21ai_1
XFILLER_20_577 VPWR VGND sg13g2_decap_8
X_3767_ _1228_ VPWR _1229_ VGND _0908_ _1227_ sg13g2_o21ai_1
X_2718_ VPWR net16 _0289_ VGND sg13g2_inv_1
X_3698_ _1183_ net654 _0943_ VPWR VGND sg13g2_nand2_1
X_2649_ _0236_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] net647
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_0_927 VPWR VGND sg13g2_decap_8
XFILLER_27_110 VPWR VGND sg13g2_decap_8
XFILLER_28_644 VPWR VGND sg13g2_decap_8
XFILLER_43_658 VPWR VGND sg13g2_decap_8
XFILLER_30_319 VPWR VGND sg13g2_fill_2
XFILLER_23_393 VPWR VGND sg13g2_decap_8
XFILLER_11_566 VPWR VGND sg13g2_decap_8
XFILLER_7_537 VPWR VGND sg13g2_decap_8
XFILLER_3_743 VPWR VGND sg13g2_decap_8
XFILLER_47_942 VPWR VGND sg13g2_decap_8
XFILLER_19_633 VPWR VGND sg13g2_decap_8
XFILLER_20_1004 VPWR VGND sg13g2_decap_8
Xfanout590 _0789_ net590 VPWR VGND sg13g2_buf_8
XFILLER_46_485 VPWR VGND sg13g2_decap_8
XFILLER_34_647 VPWR VGND sg13g2_decap_8
Xclkbuf_1_0__f_sap_3_inst.alu.clk clknet_0_sap_3_inst.alu.clk clknet_1_0__leaf_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_15_861 VPWR VGND sg13g2_decap_8
XFILLER_30_842 VPWR VGND sg13g2_decap_8
X_3621_ VGND VPWR net588 net651 _1124_ net600 sg13g2_a21oi_1
X_3552_ VPWR _1066_ _1065_ VGND sg13g2_inv_1
X_2503_ _1917_ net646 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] net722
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3483_ _1002_ _1003_ _0999_ _1005_ VPWR VGND _1004_ sg13g2_nand4_1
X_2434_ _1847_ _1853_ _1854_ VPWR VGND sg13g2_nor2_1
X_2365_ _1623_ _1704_ net764 _1785_ VPWR VGND sg13g2_nand3_1
XFILLER_37_0 VPWR VGND sg13g2_fill_1
X_4104_ net823 VGND VPWR _0068_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[2\]
+ clknet_5_3__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2296_ _1716_ net778 _1518_ VPWR VGND sg13g2_nand2_2
X_4035_ VGND VPWR _1417_ _0186_ _0194_ _1435_ sg13g2_a21oi_1
XFILLER_38_975 VPWR VGND sg13g2_decap_8
XFILLER_25_603 VPWR VGND sg13g2_decap_8
XFILLER_37_485 VPWR VGND sg13g2_decap_8
XFILLER_13_809 VPWR VGND sg13g2_decap_8
XFILLER_24_157 VPWR VGND sg13g2_fill_2
XFILLER_36_1011 VPWR VGND sg13g2_decap_8
XFILLER_40_639 VPWR VGND sg13g2_decap_8
XFILLER_21_886 VPWR VGND sg13g2_decap_8
X_3819_ net11 net608 _1265_ VPWR VGND sg13g2_nor2_1
XFILLER_4_529 VPWR VGND sg13g2_decap_8
XFILLER_43_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_724 VPWR VGND sg13g2_decap_8
XFILLER_48_717 VPWR VGND sg13g2_decap_8
XFILLER_28_441 VPWR VGND sg13g2_decap_4
XFILLER_28_452 VPWR VGND sg13g2_fill_1
XFILLER_29_986 VPWR VGND sg13g2_decap_8
XFILLER_44_967 VPWR VGND sg13g2_decap_8
XFILLER_16_647 VPWR VGND sg13g2_decap_8
XFILLER_43_455 VPWR VGND sg13g2_decap_8
XFILLER_30_138 VPWR VGND sg13g2_fill_1
XFILLER_8_824 VPWR VGND sg13g2_decap_8
XFILLER_7_323 VPWR VGND sg13g2_fill_1
XFILLER_12_875 VPWR VGND sg13g2_decap_8
XFILLER_3_540 VPWR VGND sg13g2_decap_8
X_2150_ _1562_ _1568_ _1528_ _1570_ VPWR VGND sg13g2_nand3_1
XFILLER_46_282 VPWR VGND sg13g2_fill_2
XFILLER_35_934 VPWR VGND sg13g2_decap_8
X_2983_ VPWR VGND _0537_ net627 _0536_ sap_3_inst.alu.act\[6\] _0538_ net707 sg13g2_a221oi_1
X_3604_ _1110_ net602 _1014_ VPWR VGND sg13g2_nand2_2
X_3535_ VPWR VGND net601 _1052_ _0911_ _0700_ _1053_ net596 sg13g2_a221oi_1
X_3466_ VGND VPWR _0742_ _0837_ _0989_ net653 sg13g2_a21oi_1
X_2417_ _1837_ _1836_ net756 _1821_ _1675_ VPWR VGND sg13g2_a22oi_1
X_3397_ _0899_ VPWR _0068_ VGND _0912_ _0919_ sg13g2_o21ai_1
X_2348_ VPWR VGND _1604_ _1728_ _1656_ _1597_ _1768_ _1632_ sg13g2_a221oi_1
X_2279_ _1609_ _1697_ _1698_ _1699_ VPWR VGND sg13g2_nor3_1
X_4018_ u_ser.shadow_reg\[0\] VPWR _1426_ VGND _1437_ u_ser.state\[0\] sg13g2_o21ai_1
XFILLER_25_400 VPWR VGND sg13g2_decap_8
XFILLER_26_912 VPWR VGND sg13g2_decap_8
XFILLER_38_772 VPWR VGND sg13g2_decap_8
XFILLER_13_606 VPWR VGND sg13g2_decap_8
XFILLER_26_989 VPWR VGND sg13g2_decap_8
XFILLER_41_959 VPWR VGND sg13g2_decap_8
XFILLER_25_477 VPWR VGND sg13g2_decap_8
XFILLER_21_683 VPWR VGND sg13g2_decap_8
XFILLER_5_805 VPWR VGND sg13g2_decap_8
XFILLER_0_521 VPWR VGND sg13g2_decap_8
Xclkbuf_4_14_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_14_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_48_514 VPWR VGND sg13g2_decap_8
XFILLER_0_598 VPWR VGND sg13g2_decap_8
XFILLER_29_783 VPWR VGND sg13g2_decap_8
XFILLER_17_956 VPWR VGND sg13g2_decap_8
XFILLER_44_764 VPWR VGND sg13g2_decap_8
XFILLER_32_937 VPWR VGND sg13g2_decap_8
XFILLER_8_621 VPWR VGND sg13g2_decap_8
XFILLER_12_672 VPWR VGND sg13g2_decap_8
XFILLER_8_698 VPWR VGND sg13g2_decap_8
X_3320_ net599 _0847_ _0848_ VPWR VGND sg13g2_nor2_1
XFILLER_4_893 VPWR VGND sg13g2_decap_8
XFILLER_26_1010 VPWR VGND sg13g2_decap_8
X_3251_ net702 net694 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] _0779_
+ VPWR VGND _0688_ sg13g2_nand4_1
X_2202_ net751 _1615_ _1617_ _1620_ _1622_ VPWR VGND sg13g2_and4_1
X_3182_ _0710_ _0706_ _0709_ net672 _1468_ VPWR VGND sg13g2_a22oi_1
X_2133_ net740 _1547_ _1553_ VPWR VGND sg13g2_nor2_1
XFILLER_39_558 VPWR VGND sg13g2_decap_8
X_2064_ VPWR _1486_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_35_731 VPWR VGND sg13g2_decap_8
XFILLER_23_904 VPWR VGND sg13g2_decap_8
XFILLER_22_447 VPWR VGND sg13g2_decap_8
X_2966_ VGND VPWR _0326_ _0497_ _0521_ _0332_ sg13g2_a21oi_1
X_2897_ _0453_ VPWR _0454_ VGND _0336_ _0451_ sg13g2_o21ai_1
XFILLER_2_819 VPWR VGND sg13g2_decap_8
X_3518_ _1038_ VPWR _1039_ VGND _1031_ _1033_ sg13g2_o21ai_1
X_3449_ net660 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] net670 _0972_
+ VPWR VGND sg13g2_a21o_1
XFILLER_27_45 VPWR VGND sg13g2_fill_1
XFILLER_27_78 VPWR VGND sg13g2_fill_2
XFILLER_14_926 VPWR VGND sg13g2_decap_8
XFILLER_26_786 VPWR VGND sg13g2_decap_8
Xclkbuf_4_6_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_6_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_41_756 VPWR VGND sg13g2_decap_8
XFILLER_21_480 VPWR VGND sg13g2_decap_8
XFILLER_5_602 VPWR VGND sg13g2_decap_8
XFILLER_5_679 VPWR VGND sg13g2_decap_8
XFILLER_4_38 VPWR VGND sg13g2_fill_2
XFILLER_4_27 VPWR VGND sg13g2_decap_8
XFILLER_49_834 VPWR VGND sg13g2_decap_8
XFILLER_48_311 VPWR VGND sg13g2_decap_8
XFILLER_1_885 VPWR VGND sg13g2_decap_8
XFILLER_48_388 VPWR VGND sg13g2_decap_8
XFILLER_29_580 VPWR VGND sg13g2_decap_8
XFILLER_36_528 VPWR VGND sg13g2_decap_8
XFILLER_17_753 VPWR VGND sg13g2_decap_8
XFILLER_44_561 VPWR VGND sg13g2_decap_8
XFILLER_32_734 VPWR VGND sg13g2_decap_8
X_2820_ VGND VPWR sap_3_inst.alu.act\[1\] net708 _0380_ net626 sg13g2_a21oi_1
XFILLER_13_970 VPWR VGND sg13g2_decap_8
X_2751_ VGND VPWR net736 _1824_ _0312_ net724 sg13g2_a21oi_1
XFILLER_9_952 VPWR VGND sg13g2_decap_8
X_2682_ net753 _1582_ net730 _0265_ VPWR VGND sg13g2_a21o_1
XFILLER_8_495 VPWR VGND sg13g2_decap_8
XFILLER_4_690 VPWR VGND sg13g2_decap_8
X_3303_ _0831_ net776 _0635_ VPWR VGND sg13g2_nand2_1
X_3234_ _0762_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] net676 VPWR
+ VGND sg13g2_nand2_1
X_3165_ _0693_ _0662_ net686 VPWR VGND sg13g2_nand2_2
X_3096_ _0624_ _1607_ _1622_ _0623_ VPWR VGND sg13g2_and3_1
X_2116_ _1536_ net760 net761 VPWR VGND sg13g2_xnor2_1
XFILLER_27_539 VPWR VGND sg13g2_decap_8
X_2047_ VPWR _1469_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] VGND
+ sg13g2_inv_1
XFILLER_23_701 VPWR VGND sg13g2_decap_8
X_3998_ _1409_ net710 _0515_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_778 VPWR VGND sg13g2_decap_8
X_2949_ VPWR VGND _0504_ net627 _0503_ sap_3_inst.alu.act\[5\] _0505_ net707 sg13g2_a221oi_1
XFILLER_2_616 VPWR VGND sg13g2_decap_8
XFILLER_1_159 VPWR VGND sg13g2_fill_2
XFILLER_18_539 VPWR VGND sg13g2_decap_8
XFILLER_14_723 VPWR VGND sg13g2_decap_8
XFILLER_26_583 VPWR VGND sg13g2_decap_8
XFILLER_41_553 VPWR VGND sg13g2_decap_8
XFILLER_9_204 VPWR VGND sg13g2_fill_1
XFILLER_13_277 VPWR VGND sg13g2_fill_2
XFILLER_6_922 VPWR VGND sg13g2_decap_8
XFILLER_10_984 VPWR VGND sg13g2_decap_8
Xclkload18 VPWR clkload18/Y clknet_5_25__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
XFILLER_6_999 VPWR VGND sg13g2_decap_8
XFILLER_5_476 VPWR VGND sg13g2_decap_8
XFILLER_49_631 VPWR VGND sg13g2_decap_8
XFILLER_1_682 VPWR VGND sg13g2_decap_8
XFILLER_23_1002 VPWR VGND sg13g2_decap_8
XFILLER_17_550 VPWR VGND sg13g2_decap_8
X_3921_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] _1309_
+ _1350_ net808 sg13g2_a21oi_1
XFILLER_32_531 VPWR VGND sg13g2_decap_8
X_3852_ regFile_serial_start net75 _0154_ _0159_ VPWR VGND sg13g2_a21o_1
X_2803_ _1458_ _1550_ _1796_ _0363_ VPWR VGND sg13g2_nor3_1
XFILLER_20_759 VPWR VGND sg13g2_decap_8
X_3783_ _1240_ VPWR _0135_ VGND _0996_ _1241_ sg13g2_o21ai_1
XFILLER_30_1017 VPWR VGND sg13g2_decap_8
X_2734_ net58 sap_3_inst.out\[3\] net813 _0020_ VPWR VGND sg13g2_mux2_1
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
X_2665_ net789 net795 net797 net792 _0251_ VPWR VGND sg13g2_nor4_1
X_2596_ _2000_ _2001_ _1805_ _2006_ VPWR VGND _2005_ sg13g2_nand4_1
XFILLER_5_81 VPWR VGND sg13g2_fill_1
X_3217_ net701 net696 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] _0745_
+ VPWR VGND net686 sg13g2_nand4_1
X_4197_ net846 VGND VPWR _0161_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[0\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
X_3148_ VGND VPWR net735 _1616_ _0676_ _1597_ sg13g2_a21oi_1
XFILLER_27_314 VPWR VGND sg13g2_decap_8
XFILLER_28_826 VPWR VGND sg13g2_decap_8
X_3079_ net752 net777 _0607_ VPWR VGND _0606_ sg13g2_nand3b_1
XFILLER_39_1020 VPWR VGND sg13g2_decap_8
XFILLER_36_892 VPWR VGND sg13g2_decap_8
XFILLER_23_575 VPWR VGND sg13g2_decap_8
XFILLER_11_748 VPWR VGND sg13g2_decap_8
XFILLER_7_719 VPWR VGND sg13g2_decap_8
XFILLER_40_45 VPWR VGND sg13g2_fill_1
XFILLER_3_925 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_46_1024 VPWR VGND sg13g2_decap_4
Xfanout750 _1599_ net750 VPWR VGND sg13g2_buf_8
Xfanout761 sap_3_inst.controller.stage\[0\] net761 VPWR VGND sg13g2_buf_8
Xfanout783 net784 net783 VPWR VGND sg13g2_buf_8
Xfanout772 net773 net772 VPWR VGND sg13g2_buf_8
XFILLER_19_815 VPWR VGND sg13g2_decap_8
Xfanout794 net795 net794 VPWR VGND sg13g2_buf_1
XFILLER_1_39 VPWR VGND sg13g2_fill_2
XFILLER_46_667 VPWR VGND sg13g2_decap_8
XFILLER_34_829 VPWR VGND sg13g2_decap_8
XFILLER_14_520 VPWR VGND sg13g2_decap_8
XFILLER_42_884 VPWR VGND sg13g2_decap_8
XFILLER_14_597 VPWR VGND sg13g2_decap_8
XFILLER_10_781 VPWR VGND sg13g2_decap_8
XFILLER_6_796 VPWR VGND sg13g2_decap_8
X_2450_ sap_3_inst.alu.flags\[7\] net34 _1867_ _0032_ VPWR VGND sg13g2_mux2_1
X_2381_ _1766_ _1784_ _1739_ _1801_ VPWR VGND _1799_ sg13g2_nand4_1
XFILLER_2_980 VPWR VGND sg13g2_decap_8
X_4120_ net830 VGND VPWR _0084_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\]
+ clknet_5_3__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4051_ net836 VGND VPWR _0019_ u_ser.shadow_reg\[2\] clknet_3_3__leaf_clk sg13g2_dfrbpq_1
X_3002_ VGND VPWR net790 _0338_ _0556_ _0555_ sg13g2_a21oi_1
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
XFILLER_37_667 VPWR VGND sg13g2_decap_8
XFILLER_33_840 VPWR VGND sg13g2_decap_8
XFILLER_36_188 VPWR VGND sg13g2_fill_2
X_3904_ _1335_ _1307_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] net810
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] VPWR VGND sg13g2_a22oi_1
X_3835_ net656 VPWR _1276_ VGND net599 _1040_ sg13g2_o21ai_1
XFILLER_20_556 VPWR VGND sg13g2_decap_8
X_3766_ net11 net600 _1228_ VPWR VGND sg13g2_nor2_1
X_2717_ _0289_ net577 _1819_ VPWR VGND sg13g2_nand2_2
X_3697_ _1182_ _0766_ _0835_ VPWR VGND sg13g2_xnor2_1
X_2648_ _0233_ _0234_ _0235_ VPWR VGND sg13g2_and2_1
XFILLER_0_906 VPWR VGND sg13g2_decap_8
X_2579_ _1987_ _1988_ _1989_ VPWR VGND sg13g2_and2_1
XFILLER_28_623 VPWR VGND sg13g2_decap_8
XFILLER_16_829 VPWR VGND sg13g2_decap_8
XFILLER_27_166 VPWR VGND sg13g2_decap_4
XFILLER_43_637 VPWR VGND sg13g2_decap_8
XFILLER_24_895 VPWR VGND sg13g2_decap_8
XFILLER_11_545 VPWR VGND sg13g2_decap_8
XFILLER_7_516 VPWR VGND sg13g2_decap_8
XFILLER_13_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_722 VPWR VGND sg13g2_decap_8
XFILLER_3_799 VPWR VGND sg13g2_decap_8
XFILLER_47_921 VPWR VGND sg13g2_decap_8
Xfanout580 _0321_ net580 VPWR VGND sg13g2_buf_8
XFILLER_19_612 VPWR VGND sg13g2_decap_8
Xfanout591 net592 net591 VPWR VGND sg13g2_buf_8
XFILLER_47_998 VPWR VGND sg13g2_decap_8
XFILLER_46_464 VPWR VGND sg13g2_decap_8
XFILLER_19_689 VPWR VGND sg13g2_decap_8
XFILLER_34_626 VPWR VGND sg13g2_decap_8
XFILLER_15_840 VPWR VGND sg13g2_decap_8
XFILLER_33_136 VPWR VGND sg13g2_fill_2
XFILLER_42_681 VPWR VGND sg13g2_decap_8
XFILLER_30_821 VPWR VGND sg13g2_decap_8
X_3620_ _1121_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] _1123_ _0090_
+ VPWR VGND sg13g2_a21o_1
XFILLER_30_898 VPWR VGND sg13g2_decap_8
X_3551_ _1065_ net603 _1015_ VPWR VGND sg13g2_nand2_2
X_2502_ _1916_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] net636
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3482_ _1004_ net656 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] net681
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_593 VPWR VGND sg13g2_decap_8
X_2433_ _1849_ _1850_ _1848_ _1853_ VPWR VGND _1852_ sg13g2_nand4_1
X_2364_ _1779_ _1778_ _1782_ _1784_ VPWR VGND sg13g2_a21o_2
X_4103_ net823 VGND VPWR _0067_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[1\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
X_2295_ _1441_ net763 _1715_ VPWR VGND sg13g2_nor2_2
X_4034_ VGND VPWR net814 _0186_ _1435_ net70 sg13g2_a21oi_1
XFILLER_38_954 VPWR VGND sg13g2_decap_8
XFILLER_25_659 VPWR VGND sg13g2_decap_8
XFILLER_40_618 VPWR VGND sg13g2_decap_8
XFILLER_21_865 VPWR VGND sg13g2_decap_8
X_3818_ _1263_ VPWR _0147_ VGND _0892_ _1264_ sg13g2_o21ai_1
X_3749_ _1072_ net594 _1214_ VPWR VGND sg13g2_nor2_1
XFILLER_4_508 VPWR VGND sg13g2_decap_8
XFILLER_0_703 VPWR VGND sg13g2_decap_8
XFILLER_29_965 VPWR VGND sg13g2_decap_8
XFILLER_44_946 VPWR VGND sg13g2_decap_8
XFILLER_43_434 VPWR VGND sg13g2_decap_8
XFILLER_16_626 VPWR VGND sg13g2_decap_8
XFILLER_28_497 VPWR VGND sg13g2_decap_8
XFILLER_8_803 VPWR VGND sg13g2_decap_8
XFILLER_12_854 VPWR VGND sg13g2_decap_8
XFILLER_24_692 VPWR VGND sg13g2_decap_8
XFILLER_3_596 VPWR VGND sg13g2_decap_8
X_2080_ VPWR _1502_ net60 VGND sg13g2_inv_1
XFILLER_38_239 VPWR VGND sg13g2_fill_1
XFILLER_19_464 VPWR VGND sg13g2_fill_2
XFILLER_35_913 VPWR VGND sg13g2_decap_8
XFILLER_47_795 VPWR VGND sg13g2_decap_8
XFILLER_34_456 VPWR VGND sg13g2_fill_1
XFILLER_34_467 VPWR VGND sg13g2_fill_2
X_2982_ VGND VPWR net575 _0525_ _0537_ net707 sg13g2_a21oi_1
XFILLER_22_629 VPWR VGND sg13g2_decap_8
XFILLER_21_128 VPWR VGND sg13g2_fill_1
X_3603_ _0087_ _1107_ _1109_ net619 _1482_ VPWR VGND sg13g2_a22oi_1
XFILLER_30_695 VPWR VGND sg13g2_decap_8
XFILLER_7_880 VPWR VGND sg13g2_decap_8
X_3534_ _0921_ net607 net19 _1052_ VPWR VGND sg13g2_a21o_2
X_3465_ _0988_ _0741_ _0838_ VPWR VGND sg13g2_nand2_1
X_2416_ VGND VPWR _1713_ _1832_ _1836_ _1835_ sg13g2_a21oi_1
X_3396_ _0801_ net651 _0832_ _0835_ _0922_ VPWR VGND sg13g2_and4_1
X_2347_ _1767_ _1627_ _1705_ VPWR VGND sg13g2_nand2_1
X_2278_ net744 _1691_ _1698_ VPWR VGND sg13g2_nor2_1
X_4017_ _1415_ _1424_ _1439_ _1425_ VPWR VGND sg13g2_nand3_1
XFILLER_38_751 VPWR VGND sg13g2_decap_8
XFILLER_25_456 VPWR VGND sg13g2_decap_8
XFILLER_26_968 VPWR VGND sg13g2_decap_8
XFILLER_41_938 VPWR VGND sg13g2_decap_8
XFILLER_34_990 VPWR VGND sg13g2_decap_8
XFILLER_12_139 VPWR VGND sg13g2_fill_2
XFILLER_21_662 VPWR VGND sg13g2_decap_8
XFILLER_10_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_500 VPWR VGND sg13g2_decap_8
XFILLER_0_577 VPWR VGND sg13g2_decap_8
XFILLER_29_762 VPWR VGND sg13g2_decap_8
XFILLER_17_935 VPWR VGND sg13g2_decap_8
XFILLER_44_743 VPWR VGND sg13g2_decap_8
XFILLER_32_916 VPWR VGND sg13g2_decap_8
XFILLER_40_982 VPWR VGND sg13g2_decap_8
XFILLER_8_600 VPWR VGND sg13g2_decap_8
XFILLER_12_651 VPWR VGND sg13g2_decap_8
XFILLER_8_677 VPWR VGND sg13g2_decap_8
XFILLER_11_194 VPWR VGND sg13g2_fill_2
XFILLER_4_872 VPWR VGND sg13g2_decap_8
X_3250_ net705 _0659_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] _0778_
+ VPWR VGND sg13g2_nand3_1
X_2201_ _1621_ _1582_ _1619_ VPWR VGND sg13g2_nand2_1
X_3181_ _0691_ _0701_ _0707_ _0708_ _0709_ VPWR VGND sg13g2_and4_1
X_2132_ _1552_ _1550_ _1548_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_537 VPWR VGND sg13g2_decap_8
X_2063_ VPWR _1485_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_47_592 VPWR VGND sg13g2_decap_8
XFILLER_35_710 VPWR VGND sg13g2_decap_8
XFILLER_35_787 VPWR VGND sg13g2_decap_8
XFILLER_16_990 VPWR VGND sg13g2_decap_8
X_2965_ _0520_ _0510_ _0335_ _0509_ _0344_ VPWR VGND sg13g2_a22oi_1
XFILLER_33_1015 VPWR VGND sg13g2_decap_8
X_2896_ _0453_ _0344_ _0450_ VPWR VGND sg13g2_nand2_1
XFILLER_30_492 VPWR VGND sg13g2_decap_8
X_3517_ VGND VPWR net652 _1035_ _1038_ _1037_ sg13g2_a21oi_1
X_3448_ _0971_ net674 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] net680
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] VPWR VGND sg13g2_a22oi_1
X_3379_ _0900_ _0902_ _0903_ _0904_ _0905_ VPWR VGND sg13g2_and4_1
XFILLER_27_24 VPWR VGND sg13g2_fill_1
XFILLER_45_529 VPWR VGND sg13g2_decap_8
XFILLER_14_905 VPWR VGND sg13g2_decap_8
XFILLER_26_765 VPWR VGND sg13g2_decap_8
XFILLER_41_735 VPWR VGND sg13g2_decap_8
XFILLER_22_993 VPWR VGND sg13g2_decap_8
XFILLER_5_658 VPWR VGND sg13g2_decap_8
XFILLER_49_813 VPWR VGND sg13g2_decap_8
XFILLER_1_864 VPWR VGND sg13g2_decap_8
XFILLER_48_367 VPWR VGND sg13g2_decap_8
XFILLER_36_507 VPWR VGND sg13g2_decap_8
XFILLER_17_732 VPWR VGND sg13g2_decap_8
XFILLER_44_540 VPWR VGND sg13g2_decap_8
XFILLER_16_231 VPWR VGND sg13g2_fill_2
XFILLER_32_713 VPWR VGND sg13g2_decap_8
XFILLER_9_931 VPWR VGND sg13g2_decap_8
X_2750_ _0300_ VPWR _0311_ VGND _0309_ _0310_ sg13g2_o21ai_1
X_2681_ _0262_ _0263_ _0261_ _0264_ VPWR VGND sg13g2_nand3_1
X_3302_ _0830_ _0808_ net606 VPWR VGND sg13g2_nand2_1
X_3233_ _0761_ net666 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] net671
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_27_518 VPWR VGND sg13g2_decap_8
X_3164_ net704 net702 _0658_ net689 _0692_ VPWR VGND sg13g2_nor4_1
X_3095_ _0620_ _0621_ _0622_ _0623_ VPWR VGND sg13g2_or3_1
X_2115_ _1535_ _1505_ _1534_ VPWR VGND sg13g2_nand2_2
X_2046_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[0\] _1468_ VPWR VGND
+ sg13g2_inv_4
XFILLER_35_584 VPWR VGND sg13g2_decap_8
XFILLER_23_757 VPWR VGND sg13g2_decap_8
X_3997_ _1406_ VPWR _0182_ VGND net583 _1408_ sg13g2_o21ai_1
X_2948_ VGND VPWR net575 _0488_ _0504_ net707 sg13g2_a21oi_1
X_2879_ _0437_ _0436_ _0326_ _0434_ net625 VPWR VGND sg13g2_a22oi_1
XFILLER_8_8 VPWR VGND sg13g2_fill_2
XFILLER_1_105 VPWR VGND sg13g2_fill_2
XFILLER_46_849 VPWR VGND sg13g2_decap_8
XFILLER_18_518 VPWR VGND sg13g2_decap_8
XFILLER_14_702 VPWR VGND sg13g2_decap_8
XFILLER_26_562 VPWR VGND sg13g2_decap_8
XFILLER_41_532 VPWR VGND sg13g2_decap_8
XFILLER_14_779 VPWR VGND sg13g2_decap_8
XFILLER_22_790 VPWR VGND sg13g2_decap_8
XFILLER_6_901 VPWR VGND sg13g2_decap_8
XFILLER_10_963 VPWR VGND sg13g2_decap_8
Xclkload19 VPWR clkload19/Y clknet_5_29__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
XFILLER_6_978 VPWR VGND sg13g2_decap_8
XFILLER_1_661 VPWR VGND sg13g2_decap_8
XFILLER_49_610 VPWR VGND sg13g2_decap_8
XFILLER_49_687 VPWR VGND sg13g2_decap_8
XFILLER_37_849 VPWR VGND sg13g2_decap_8
X_3920_ net811 net63 _1349_ _0164_ VPWR VGND sg13g2_a21o_1
XFILLER_45_893 VPWR VGND sg13g2_decap_8
X_4045__10 VPWR net46 clknet_leaf_1_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_32_510 VPWR VGND sg13g2_decap_8
X_3851_ VGND VPWR _1440_ _1285_ _0158_ _1282_ sg13g2_a21oi_1
X_3782_ net660 _0984_ _1241_ VPWR VGND _1159_ sg13g2_nand3b_1
X_2802_ net775 _1951_ _1956_ _0355_ _0362_ VPWR VGND sg13g2_nor4_1
XFILLER_20_738 VPWR VGND sg13g2_decap_8
XFILLER_32_587 VPWR VGND sg13g2_decap_8
X_2733_ net64 sap_3_inst.out\[2\] net813 _0019_ VPWR VGND sg13g2_mux2_1
X_2664_ VGND VPWR net17 _0250_ _0239_ sg13g2_or2_1
X_2595_ _2005_ net644 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] net723
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_28_805 VPWR VGND sg13g2_decap_8
X_4196_ net846 VGND VPWR _0160_ regFile_serial clknet_3_6__leaf_clk sg13g2_dfrbpq_1
X_3216_ net704 net698 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] _0744_
+ VPWR VGND net694 sg13g2_nand4_1
X_3147_ VPWR VGND _1630_ _0674_ _0673_ net750 _0675_ _0671_ sg13g2_a221oi_1
XFILLER_43_819 VPWR VGND sg13g2_decap_8
X_3078_ _0606_ _1642_ _1532_ net747 net760 VPWR VGND sg13g2_a22oi_1
XFILLER_36_871 VPWR VGND sg13g2_decap_8
X_2029_ VPWR _1451_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] VGND
+ sg13g2_inv_1
Xclkbuf_5_9__f_sap_3_inst.alu.clk_regs clknet_4_4_0_sap_3_inst.alu.clk_regs clknet_5_9__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_23_554 VPWR VGND sg13g2_decap_8
XFILLER_11_727 VPWR VGND sg13g2_decap_8
XFILLER_3_904 VPWR VGND sg13g2_decap_8
XFILLER_46_1003 VPWR VGND sg13g2_decap_8
Xfanout751 _1596_ net751 VPWR VGND sg13g2_buf_8
Xfanout740 net741 net740 VPWR VGND sg13g2_buf_8
Xfanout784 sap_3_inst.controller.opcode\[1\] net784 VPWR VGND sg13g2_buf_8
Xfanout762 sap_3_inst.alu.flags\[1\] net762 VPWR VGND sg13g2_buf_8
Xfanout773 sap_3_inst.controller.opcode\[5\] net773 VPWR VGND sg13g2_buf_8
Xfanout795 sap_3_inst.alu.acc\[5\] net795 VPWR VGND sg13g2_buf_8
XFILLER_46_646 VPWR VGND sg13g2_decap_8
XFILLER_45_112 VPWR VGND sg13g2_fill_1
XFILLER_34_808 VPWR VGND sg13g2_decap_8
XFILLER_27_882 VPWR VGND sg13g2_decap_8
XFILLER_42_863 VPWR VGND sg13g2_decap_8
XFILLER_14_576 VPWR VGND sg13g2_decap_8
XFILLER_10_760 VPWR VGND sg13g2_decap_8
XFILLER_6_775 VPWR VGND sg13g2_decap_8
X_2380_ _1738_ _1765_ _1783_ _1800_ VGND VPWR _1798_ sg13g2_nor4_2
X_4050_ net832 VGND VPWR _0018_ u_ser.shadow_reg\[1\] clknet_3_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_49_484 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
X_3001_ _0555_ sap_3_inst.alu.flags\[1\] _1957_ net682 VPWR VGND sg13g2_and3_1
XFILLER_37_646 VPWR VGND sg13g2_decap_8
XFILLER_24_307 VPWR VGND sg13g2_fill_1
XFILLER_36_145 VPWR VGND sg13g2_fill_1
XFILLER_45_690 VPWR VGND sg13g2_decap_8
XFILLER_18_882 VPWR VGND sg13g2_decap_8
Xclkbuf_5_16__f_sap_3_inst.alu.clk_regs clknet_4_8_0_sap_3_inst.alu.clk_regs clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3903_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] _1306_
+ _1334_ net808 sg13g2_a21oi_1
XFILLER_33_896 VPWR VGND sg13g2_decap_8
X_3834_ VPWR VGND net712 _1070_ _1274_ _1030_ _1275_ _1273_ sg13g2_a221oi_1
XFILLER_20_535 VPWR VGND sg13g2_decap_8
X_3765_ _1227_ _0872_ _1226_ VPWR VGND sg13g2_nand2_1
X_3696_ _1181_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] net578 VPWR
+ VGND sg13g2_nand2_1
X_2716_ net576 _1876_ net15 VPWR VGND sg13g2_and2_1
X_2647_ _0234_ net637 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] net722
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_10_49 VPWR VGND sg13g2_fill_2
X_2578_ _1988_ net630 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] net639
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_28_602 VPWR VGND sg13g2_decap_8
X_4179_ net825 VGND VPWR _0143_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\]
+ clknet_5_9__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_16_808 VPWR VGND sg13g2_decap_8
XFILLER_43_616 VPWR VGND sg13g2_decap_8
XFILLER_28_679 VPWR VGND sg13g2_decap_8
XFILLER_24_874 VPWR VGND sg13g2_decap_8
XFILLER_11_524 VPWR VGND sg13g2_decap_8
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_3_701 VPWR VGND sg13g2_decap_8
XFILLER_3_778 VPWR VGND sg13g2_decap_8
XFILLER_47_900 VPWR VGND sg13g2_decap_8
Xfanout581 _0321_ net581 VPWR VGND sg13g2_buf_8
Xfanout592 _0788_ net592 VPWR VGND sg13g2_buf_8
XFILLER_46_443 VPWR VGND sg13g2_decap_8
XFILLER_47_977 VPWR VGND sg13g2_decap_8
XFILLER_19_668 VPWR VGND sg13g2_decap_8
XFILLER_34_605 VPWR VGND sg13g2_decap_8
XFILLER_42_660 VPWR VGND sg13g2_decap_8
XFILLER_15_896 VPWR VGND sg13g2_decap_8
XFILLER_30_800 VPWR VGND sg13g2_decap_8
XFILLER_30_877 VPWR VGND sg13g2_decap_8
X_3550_ VGND VPWR net33 _1064_ _1009_ net606 sg13g2_a21oi_2
XFILLER_6_572 VPWR VGND sg13g2_decap_8
X_2501_ _1912_ _1914_ _1915_ VPWR VGND sg13g2_and2_1
X_3481_ _1003_ net660 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] net679
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2432_ net737 _1851_ _1852_ VPWR VGND sg13g2_nor2_1
X_2363_ VGND VPWR _1782_ _1783_ _1779_ _1778_ sg13g2_a21oi_2
X_4102_ net823 VGND VPWR _0066_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[0\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
X_4033_ VGND VPWR net814 _0186_ _0193_ _1434_ sg13g2_a21oi_1
X_2294_ _1714_ _1541_ _1712_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_933 VPWR VGND sg13g2_decap_8
XFILLER_49_281 VPWR VGND sg13g2_decap_8
XFILLER_25_638 VPWR VGND sg13g2_decap_8
XFILLER_21_844 VPWR VGND sg13g2_decap_8
XFILLER_33_693 VPWR VGND sg13g2_decap_8
X_3817_ _0893_ net655 _1264_ VPWR VGND _0887_ sg13g2_nand3b_1
X_3748_ VGND VPWR _1488_ net593 _0128_ _1213_ sg13g2_a21oi_1
X_3679_ net712 VPWR _1168_ VGND _0289_ _1138_ sg13g2_o21ai_1
XFILLER_0_759 VPWR VGND sg13g2_decap_8
XFILLER_47_218 VPWR VGND sg13g2_fill_1
XFILLER_29_944 VPWR VGND sg13g2_decap_8
XFILLER_44_925 VPWR VGND sg13g2_decap_8
XFILLER_16_605 VPWR VGND sg13g2_decap_8
XFILLER_28_476 VPWR VGND sg13g2_decap_8
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_24_671 VPWR VGND sg13g2_decap_8
XFILLER_31_619 VPWR VGND sg13g2_decap_8
XFILLER_12_833 VPWR VGND sg13g2_decap_8
XFILLER_8_859 VPWR VGND sg13g2_decap_8
XFILLER_3_575 VPWR VGND sg13g2_decap_8
XFILLER_39_719 VPWR VGND sg13g2_decap_8
XFILLER_47_774 VPWR VGND sg13g2_decap_8
XFILLER_22_608 VPWR VGND sg13g2_decap_8
XFILLER_35_969 VPWR VGND sg13g2_decap_8
XFILLER_43_980 VPWR VGND sg13g2_decap_8
X_2981_ _0528_ _0535_ _0523_ _0536_ VPWR VGND sg13g2_nand3_1
XFILLER_15_693 VPWR VGND sg13g2_decap_8
XFILLER_30_674 VPWR VGND sg13g2_decap_8
X_3602_ _1109_ _0980_ _1108_ VPWR VGND sg13g2_nand2_1
X_3533_ _0075_ _1049_ _1051_ net584 _1467_ VPWR VGND sg13g2_a22oi_1
XFILLER_42_0 VPWR VGND sg13g2_fill_1
X_3464_ _0987_ _0741_ _0803_ VPWR VGND sg13g2_xnor2_1
X_2415_ VGND VPWR _1514_ _1833_ _1835_ _1834_ sg13g2_a21oi_1
X_3395_ _0920_ VPWR _0921_ VGND net590 _0801_ sg13g2_o21ai_1
X_2346_ _1766_ _1765_ VPWR VGND sg13g2_inv_2
X_2277_ net742 _1629_ _1697_ VPWR VGND sg13g2_nor2_2
XFILLER_38_730 VPWR VGND sg13g2_decap_8
X_4016_ net814 u_ser.shadow_reg\[1\] u_ser.shadow_reg\[2\] u_ser.shadow_reg\[3\] u_ser.shadow_reg\[4\]
+ u_ser.bit_pos\[1\] _1424_ VPWR VGND sg13g2_mux4_1
XFILLER_26_947 VPWR VGND sg13g2_decap_8
XFILLER_41_917 VPWR VGND sg13g2_decap_8
XFILLER_25_435 VPWR VGND sg13g2_decap_8
XFILLER_33_490 VPWR VGND sg13g2_decap_8
XFILLER_21_641 VPWR VGND sg13g2_decap_8
X_4042__7 VPWR net43 clknet_leaf_2_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_10_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_556 VPWR VGND sg13g2_decap_8
XFILLER_48_549 VPWR VGND sg13g2_decap_8
XFILLER_17_914 VPWR VGND sg13g2_decap_8
XFILLER_29_741 VPWR VGND sg13g2_decap_8
XFILLER_44_722 VPWR VGND sg13g2_decap_8
XFILLER_44_799 VPWR VGND sg13g2_decap_8
XFILLER_12_630 VPWR VGND sg13g2_decap_8
XFILLER_40_961 VPWR VGND sg13g2_decap_8
XFILLER_8_656 VPWR VGND sg13g2_decap_8
XFILLER_4_851 VPWR VGND sg13g2_decap_8
X_2200_ _1581_ _1618_ _1620_ VPWR VGND sg13g2_nor2_2
X_3180_ _0708_ net667 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] net678
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_516 VPWR VGND sg13g2_decap_8
X_2131_ _1548_ _1549_ _1551_ VPWR VGND sg13g2_nor2_2
X_2062_ _1484_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[6\] VPWR VGND
+ sg13g2_inv_2
XFILLER_47_571 VPWR VGND sg13g2_decap_8
XFILLER_35_766 VPWR VGND sg13g2_decap_8
XFILLER_23_939 VPWR VGND sg13g2_decap_8
X_2964_ _0519_ _0342_ _0508_ _0340_ net787 VPWR VGND sg13g2_a22oi_1
XFILLER_15_490 VPWR VGND sg13g2_decap_8
XFILLER_8_60 VPWR VGND sg13g2_fill_1
X_2895_ VPWR _0452_ _0451_ VGND sg13g2_inv_1
XFILLER_31_983 VPWR VGND sg13g2_decap_8
X_3516_ VGND VPWR net34 net595 _1037_ _1036_ sg13g2_a21oi_1
X_3447_ _0970_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[5\] net587 VPWR
+ VGND sg13g2_nand2_1
X_3378_ _0904_ net678 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] net680
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2329_ _1581_ _1597_ _1618_ _1749_ VPWR VGND sg13g2_nor3_1
XFILLER_45_508 VPWR VGND sg13g2_decap_8
XFILLER_26_744 VPWR VGND sg13g2_decap_8
XFILLER_41_714 VPWR VGND sg13g2_decap_8
XFILLER_43_68 VPWR VGND sg13g2_fill_2
XFILLER_22_972 VPWR VGND sg13g2_decap_8
XFILLER_40_257 VPWR VGND sg13g2_fill_2
XFILLER_5_637 VPWR VGND sg13g2_decap_8
XFILLER_49_1023 VPWR VGND sg13g2_decap_4
XFILLER_4_158 VPWR VGND sg13g2_fill_1
XFILLER_1_843 VPWR VGND sg13g2_decap_8
XFILLER_49_869 VPWR VGND sg13g2_decap_8
XFILLER_48_346 VPWR VGND sg13g2_decap_8
XFILLER_1_1025 VPWR VGND sg13g2_decap_4
XFILLER_17_711 VPWR VGND sg13g2_decap_8
XFILLER_17_788 VPWR VGND sg13g2_decap_8
XFILLER_44_596 VPWR VGND sg13g2_decap_8
XFILLER_9_910 VPWR VGND sg13g2_decap_8
XFILLER_32_769 VPWR VGND sg13g2_decap_8
XFILLER_12_460 VPWR VGND sg13g2_fill_1
X_2680_ _1608_ VPWR _0263_ VGND net744 _1644_ sg13g2_o21ai_1
XFILLER_9_987 VPWR VGND sg13g2_decap_8
X_3301_ _0829_ net653 net711 VPWR VGND sg13g2_nand2_2
X_3232_ net703 net690 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] _0760_
+ VPWR VGND sg13g2_nand3_1
X_3163_ _0691_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] net674 VPWR
+ VGND sg13g2_nand2_1
X_2114_ net761 net760 _1534_ VPWR VGND sg13g2_nor2b_2
XFILLER_39_346 VPWR VGND sg13g2_fill_2
X_3094_ _1573_ _1575_ _0622_ VPWR VGND sg13g2_nor2_1
X_2045_ VPWR _1467_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] VGND
+ sg13g2_inv_1
XFILLER_35_563 VPWR VGND sg13g2_decap_8
XFILLER_23_736 VPWR VGND sg13g2_decap_8
X_3996_ VGND VPWR _0496_ net710 _1408_ _1407_ sg13g2_a21oi_1
XFILLER_10_408 VPWR VGND sg13g2_fill_2
XFILLER_11_909 VPWR VGND sg13g2_decap_8
XFILLER_22_268 VPWR VGND sg13g2_fill_2
X_2947_ net575 _0481_ _0499_ _0502_ _0503_ VPWR VGND sg13g2_or4_1
XFILLER_31_780 VPWR VGND sg13g2_decap_8
X_2878_ _0434_ _0389_ _0435_ _0436_ VPWR VGND sg13g2_a21o_1
XFILLER_46_828 VPWR VGND sg13g2_decap_8
XFILLER_39_880 VPWR VGND sg13g2_decap_8
XFILLER_26_541 VPWR VGND sg13g2_decap_8
XFILLER_41_511 VPWR VGND sg13g2_decap_8
XFILLER_14_758 VPWR VGND sg13g2_decap_8
XFILLER_16_1011 VPWR VGND sg13g2_decap_8
XFILLER_41_588 VPWR VGND sg13g2_decap_8
XFILLER_13_279 VPWR VGND sg13g2_fill_1
XFILLER_10_942 VPWR VGND sg13g2_decap_8
XFILLER_6_957 VPWR VGND sg13g2_decap_8
XFILLER_1_640 VPWR VGND sg13g2_decap_8
XFILLER_49_666 VPWR VGND sg13g2_decap_8
XFILLER_37_828 VPWR VGND sg13g2_decap_8
XFILLER_45_872 VPWR VGND sg13g2_decap_8
XFILLER_44_393 VPWR VGND sg13g2_decap_8
XFILLER_17_585 VPWR VGND sg13g2_decap_8
XFILLER_32_566 VPWR VGND sg13g2_decap_8
X_3850_ _1282_ _1284_ _1286_ _0157_ VPWR VGND sg13g2_nor3_1
X_3781_ _1240_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] net611 VPWR
+ VGND sg13g2_nand2_1
Xclkbuf_0_sap_3_inst.alu.clk sap_3_inst.alu.clk clknet_0_sap_3_inst.alu.clk VPWR VGND
+ sg13g2_buf_8
X_2801_ _0361_ _0348_ _0359_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_717 VPWR VGND sg13g2_decap_8
X_2732_ net59 sap_3_inst.out\[1\] net813 _0018_ VPWR VGND sg13g2_mux2_1
XFILLER_9_784 VPWR VGND sg13g2_decap_8
X_2663_ _0243_ VPWR _0250_ VGND _1673_ _0249_ sg13g2_o21ai_1
X_2594_ _2004_ _2002_ _2003_ VPWR VGND sg13g2_nand2_1
X_3215_ net698 net691 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] _0743_
+ VPWR VGND net686 sg13g2_nand4_1
X_4195_ net846 VGND VPWR net76 regFile_serial_start clknet_3_6__leaf_clk sg13g2_dfrbpq_1
X_3146_ _0674_ net730 net726 _1620_ net749 VPWR VGND sg13g2_a22oi_1
X_3077_ _0604_ VPWR _0605_ VGND _1594_ _1850_ sg13g2_o21ai_1
X_2028_ VPWR _1450_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_36_850 VPWR VGND sg13g2_decap_8
XFILLER_23_533 VPWR VGND sg13g2_decap_8
XFILLER_11_706 VPWR VGND sg13g2_decap_8
X_3979_ VGND VPWR _0359_ net709 _1395_ _1394_ sg13g2_a21oi_1
XFILLER_40_14 VPWR VGND sg13g2_fill_1
Xfanout730 _1633_ net730 VPWR VGND sg13g2_buf_8
Xfanout741 net742 net741 VPWR VGND sg13g2_buf_8
Xfanout752 _1595_ net752 VPWR VGND sg13g2_buf_8
Xfanout785 net786 net785 VPWR VGND sg13g2_buf_8
Xfanout774 net775 net774 VPWR VGND sg13g2_buf_8
Xfanout763 net764 net763 VPWR VGND sg13g2_buf_8
XFILLER_46_625 VPWR VGND sg13g2_decap_8
Xfanout796 net797 net796 VPWR VGND sg13g2_buf_8
XFILLER_27_861 VPWR VGND sg13g2_decap_8
XFILLER_42_842 VPWR VGND sg13g2_decap_8
XFILLER_14_555 VPWR VGND sg13g2_decap_8
XFILLER_6_754 VPWR VGND sg13g2_decap_8
XFILLER_7_1020 VPWR VGND sg13g2_decap_8
XFILLER_49_463 VPWR VGND sg13g2_decap_8
X_3000_ _0332_ _0552_ _0554_ VPWR VGND sg13g2_and2_1
XFILLER_37_625 VPWR VGND sg13g2_decap_8
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
XFILLER_18_861 VPWR VGND sg13g2_decap_8
X_3902_ _1333_ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] _1314_
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_514 VPWR VGND sg13g2_decap_8
XFILLER_33_875 VPWR VGND sg13g2_decap_8
X_3833_ net656 net653 _0289_ _1274_ VPWR VGND sg13g2_nand3_1
X_3764_ _1226_ _0888_ _0907_ VPWR VGND sg13g2_nand2_1
XFILLER_9_581 VPWR VGND sg13g2_decap_8
X_3695_ net578 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] _1180_ _0108_
+ VPWR VGND sg13g2_a21o_1
X_2715_ VPWR net14 _0288_ VGND sg13g2_inv_1
X_2646_ _0233_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] net638
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2577_ _1987_ net633 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] net635
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] VPWR VGND sg13g2_a22oi_1
X_4178_ net842 VGND VPWR _0142_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_658 VPWR VGND sg13g2_decap_8
X_3129_ _0654_ _0656_ _0657_ VPWR VGND sg13g2_and2_1
XFILLER_24_853 VPWR VGND sg13g2_decap_8
XFILLER_11_503 VPWR VGND sg13g2_decap_8
XFILLER_23_352 VPWR VGND sg13g2_fill_1
XFILLER_3_757 VPWR VGND sg13g2_decap_8
Xfanout582 _1390_ net582 VPWR VGND sg13g2_buf_8
Xfanout593 _1208_ net593 VPWR VGND sg13g2_buf_8
XFILLER_47_956 VPWR VGND sg13g2_decap_8
XFILLER_46_422 VPWR VGND sg13g2_decap_8
XFILLER_19_647 VPWR VGND sg13g2_decap_8
XFILLER_20_1018 VPWR VGND sg13g2_decap_8
XFILLER_46_499 VPWR VGND sg13g2_decap_8
XFILLER_15_875 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_2_sap_3_inst.alu.clk clknet_1_0__leaf_sap_3_inst.alu.clk clknet_leaf_2_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_30_856 VPWR VGND sg13g2_decap_8
X_3480_ _1002_ net665 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] net668
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_551 VPWR VGND sg13g2_decap_8
X_2500_ _1914_ net630 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] net644
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] VPWR VGND sg13g2_a22oi_1
X_2431_ _1504_ net766 _1524_ _1558_ _1851_ VPWR VGND sg13g2_nor4_1
XFILLER_29_1021 VPWR VGND sg13g2_decap_8
X_2362_ _1762_ _1781_ net757 _1782_ VPWR VGND sg13g2_nand3_1
X_2293_ _1712_ _1541_ _1713_ VPWR VGND sg13g2_nor2b_2
X_4101_ net818 VGND VPWR _0065_ sap_3_inst.controller.opcode\[7\] clknet_5_1__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_4032_ net814 _1415_ _1434_ VPWR VGND sg13g2_nor2_1
XFILLER_38_912 VPWR VGND sg13g2_decap_8
XFILLER_38_989 VPWR VGND sg13g2_decap_8
XFILLER_25_617 VPWR VGND sg13g2_decap_8
XFILLER_37_499 VPWR VGND sg13g2_decap_8
XFILLER_21_823 VPWR VGND sg13g2_decap_8
XFILLER_33_672 VPWR VGND sg13g2_decap_8
XFILLER_36_1025 VPWR VGND sg13g2_decap_4
X_3816_ _1263_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] net610 VPWR
+ VGND sg13g2_nand2_1
X_3747_ net593 _1212_ _1213_ VPWR VGND sg13g2_nor2_1
X_3678_ _1161_ VPWR _0104_ VGND _1164_ _1167_ sg13g2_o21ai_1
X_2629_ _0218_ _0215_ _0217_ _1858_ net2 VPWR VGND sg13g2_a22oi_1
XFILLER_0_738 VPWR VGND sg13g2_decap_8
XFILLER_47_208 VPWR VGND sg13g2_fill_1
XFILLER_29_923 VPWR VGND sg13g2_decap_8
XFILLER_44_904 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_12_812 VPWR VGND sg13g2_decap_8
XFILLER_24_650 VPWR VGND sg13g2_decap_8
XFILLER_30_119 VPWR VGND sg13g2_fill_1
XFILLER_11_311 VPWR VGND sg13g2_fill_2
XFILLER_8_838 VPWR VGND sg13g2_decap_8
XFILLER_12_889 VPWR VGND sg13g2_decap_8
XFILLER_3_554 VPWR VGND sg13g2_decap_8
XFILLER_11_82 VPWR VGND sg13g2_fill_2
XFILLER_4_1012 VPWR VGND sg13g2_decap_8
XFILLER_47_753 VPWR VGND sg13g2_decap_8
XFILLER_19_466 VPWR VGND sg13g2_fill_1
XFILLER_35_948 VPWR VGND sg13g2_decap_8
XFILLER_36_90 VPWR VGND sg13g2_fill_1
X_2980_ _0533_ _0534_ _1944_ _0535_ VPWR VGND sg13g2_nand3_1
XFILLER_15_672 VPWR VGND sg13g2_decap_8
XFILLER_34_469 VPWR VGND sg13g2_fill_1
XFILLER_30_653 VPWR VGND sg13g2_decap_8
X_3601_ VGND VPWR net619 _0981_ _1108_ net599 sg13g2_a21oi_1
X_3532_ net18 _1050_ _1051_ VPWR VGND sg13g2_nor2_1
X_3463_ net587 _0983_ _0985_ _0986_ VPWR VGND sg13g2_or3_1
X_2414_ net724 VPWR _1834_ VGND _1543_ net732 sg13g2_o21ai_1
X_3394_ net589 net591 _0775_ _0920_ VPWR VGND sg13g2_a21o_1
XFILLER_35_0 VPWR VGND sg13g2_fill_1
X_2345_ VGND VPWR _1763_ _1765_ _1759_ net756 sg13g2_a21oi_2
X_2276_ _1567_ VPWR _1696_ VGND _1579_ _1599_ sg13g2_o21ai_1
X_4015_ _1415_ _1422_ u_ser.bit_pos\[2\] _1423_ VPWR VGND sg13g2_nand3_1
XFILLER_25_414 VPWR VGND sg13g2_decap_8
XFILLER_26_926 VPWR VGND sg13g2_decap_8
XFILLER_38_786 VPWR VGND sg13g2_decap_8
XFILLER_21_620 VPWR VGND sg13g2_decap_8
XFILLER_40_439 VPWR VGND sg13g2_decap_4
XFILLER_21_697 VPWR VGND sg13g2_decap_8
XFILLER_5_819 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_535 VPWR VGND sg13g2_decap_8
XFILLER_48_528 VPWR VGND sg13g2_decap_8
XFILLER_29_720 VPWR VGND sg13g2_decap_8
XFILLER_44_701 VPWR VGND sg13g2_decap_8
XFILLER_43_200 VPWR VGND sg13g2_fill_2
XFILLER_29_797 VPWR VGND sg13g2_decap_8
XFILLER_44_778 VPWR VGND sg13g2_decap_8
XFILLER_25_981 VPWR VGND sg13g2_decap_8
XFILLER_40_940 VPWR VGND sg13g2_decap_8
XFILLER_8_635 VPWR VGND sg13g2_decap_8
XFILLER_12_686 VPWR VGND sg13g2_decap_8
XFILLER_11_196 VPWR VGND sg13g2_fill_1
XFILLER_4_830 VPWR VGND sg13g2_decap_8
XFILLER_26_1024 VPWR VGND sg13g2_decap_4
X_2130_ _1523_ net781 _1550_ VPWR VGND net783 sg13g2_nand3b_1
XFILLER_47_550 VPWR VGND sg13g2_decap_8
X_2061_ VPWR _1483_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] VGND
+ sg13g2_inv_1
XFILLER_19_285 VPWR VGND sg13g2_fill_2
XFILLER_35_745 VPWR VGND sg13g2_decap_8
XFILLER_23_918 VPWR VGND sg13g2_decap_8
XFILLER_34_266 VPWR VGND sg13g2_fill_2
X_2963_ VGND VPWR net794 net683 _0518_ _0517_ sg13g2_a21oi_1
XFILLER_31_962 VPWR VGND sg13g2_decap_8
X_2894_ _0451_ net797 sap_3_inst.alu.tmp\[4\] VPWR VGND sg13g2_xnor2_1
XFILLER_30_450 VPWR VGND sg13g2_fill_1
X_3515_ net712 VPWR _1036_ VGND _0289_ net595 sg13g2_o21ai_1
X_3446_ _0969_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[4\] net586 _0070_
+ VPWR VGND sg13g2_mux2_1
X_3377_ _0903_ net657 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] net667
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2328_ VGND VPWR _1593_ _1638_ _1748_ _1576_ sg13g2_a21oi_1
X_2259_ VGND VPWR _1676_ net729 _1679_ _1539_ sg13g2_a21oi_1
XFILLER_26_723 VPWR VGND sg13g2_decap_8
XFILLER_38_583 VPWR VGND sg13g2_decap_8
XFILLER_22_951 VPWR VGND sg13g2_decap_8
XFILLER_21_494 VPWR VGND sg13g2_decap_8
XFILLER_5_616 VPWR VGND sg13g2_decap_8
XFILLER_49_1002 VPWR VGND sg13g2_decap_8
XFILLER_1_822 VPWR VGND sg13g2_decap_8
XFILLER_49_848 VPWR VGND sg13g2_decap_8
XFILLER_48_325 VPWR VGND sg13g2_decap_8
XFILLER_1_899 VPWR VGND sg13g2_decap_8
XFILLER_1_1004 VPWR VGND sg13g2_decap_8
XFILLER_29_594 VPWR VGND sg13g2_decap_8
XFILLER_44_575 VPWR VGND sg13g2_decap_8
XFILLER_17_767 VPWR VGND sg13g2_decap_8
XFILLER_32_748 VPWR VGND sg13g2_decap_8
XFILLER_13_984 VPWR VGND sg13g2_decap_8
XFILLER_9_966 VPWR VGND sg13g2_decap_8
XFILLER_12_483 VPWR VGND sg13g2_decap_8
XFILLER_33_91 VPWR VGND sg13g2_fill_1
X_3300_ net651 net712 _0828_ VPWR VGND sg13g2_nor2_2
X_3231_ _0759_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] net690 net687
+ VPWR VGND sg13g2_and3_1
X_3162_ _0690_ net690 net686 VPWR VGND sg13g2_nand2_2
X_2113_ _1533_ _1505_ _1532_ VPWR VGND sg13g2_nand2_2
X_3093_ _1570_ net726 _0621_ VPWR VGND sg13g2_nor2_1
XFILLER_48_892 VPWR VGND sg13g2_decap_8
X_2044_ VPWR _1466_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] VGND
+ sg13g2_inv_1
XFILLER_23_715 VPWR VGND sg13g2_decap_8
XFILLER_35_542 VPWR VGND sg13g2_decap_8
XFILLER_22_203 VPWR VGND sg13g2_fill_2
X_3995_ net710 net793 _1407_ VPWR VGND sg13g2_nor2b_1
X_2946_ _0501_ VPWR _0502_ VGND _0328_ _0490_ sg13g2_o21ai_1
X_2877_ _0348_ _0359_ _0384_ _0435_ VGND VPWR _0422_ sg13g2_nor4_2
XFILLER_1_107 VPWR VGND sg13g2_fill_1
X_3429_ _0953_ _0949_ _0952_ net671 _1474_ VPWR VGND sg13g2_a22oi_1
XFILLER_46_807 VPWR VGND sg13g2_decap_8
XFILLER_26_520 VPWR VGND sg13g2_decap_8
XFILLER_14_737 VPWR VGND sg13g2_decap_8
XFILLER_26_597 VPWR VGND sg13g2_decap_8
XFILLER_41_567 VPWR VGND sg13g2_decap_8
XFILLER_13_247 VPWR VGND sg13g2_fill_2
XFILLER_10_921 VPWR VGND sg13g2_decap_8
XFILLER_6_936 VPWR VGND sg13g2_decap_8
XFILLER_5_435 VPWR VGND sg13g2_fill_2
XFILLER_10_998 VPWR VGND sg13g2_decap_8
Xclkbuf_5_24__f_sap_3_inst.alu.clk_regs clknet_4_12_0_sap_3_inst.alu.clk_regs clknet_5_24__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_0_162 VPWR VGND sg13g2_fill_1
XFILLER_1_696 VPWR VGND sg13g2_decap_8
XFILLER_49_645 VPWR VGND sg13g2_decap_8
XFILLER_0_184 VPWR VGND sg13g2_fill_2
XFILLER_23_1016 VPWR VGND sg13g2_decap_8
XFILLER_23_1027 VPWR VGND sg13g2_fill_2
XFILLER_37_807 VPWR VGND sg13g2_decap_8
XFILLER_45_851 VPWR VGND sg13g2_decap_8
XFILLER_17_564 VPWR VGND sg13g2_decap_8
XFILLER_44_372 VPWR VGND sg13g2_decap_8
XFILLER_32_545 VPWR VGND sg13g2_decap_8
X_2800_ _0348_ _0359_ _0360_ VPWR VGND sg13g2_nor2_1
X_3780_ _0134_ _1099_ _1239_ net613 _1477_ VPWR VGND sg13g2_a22oi_1
X_2731_ net69 sap_3_inst.out\[0\] net813 _0017_ VPWR VGND sg13g2_mux2_1
XFILLER_9_763 VPWR VGND sg13g2_decap_8
XFILLER_13_781 VPWR VGND sg13g2_decap_8
X_2662_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] _0248_
+ net638 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] _0249_ net645 sg13g2_a221oi_1
X_2593_ _2003_ net630 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] net639
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_980 VPWR VGND sg13g2_decap_8
X_3214_ _0735_ _0738_ _0734_ _0742_ VPWR VGND _0740_ sg13g2_nand4_1
X_4194_ net847 VGND VPWR _0158_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_2
X_3145_ _0673_ _0670_ _0672_ _1614_ _1609_ VPWR VGND sg13g2_a22oi_1
X_3076_ _0604_ _1851_ _1746_ VPWR VGND sg13g2_nand2b_1
X_2027_ VPWR _1449_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_23_512 VPWR VGND sg13g2_decap_8
X_3978_ _1458_ net709 _1394_ VPWR VGND sg13g2_nor2_1
XFILLER_23_589 VPWR VGND sg13g2_decap_8
X_2929_ _0482_ _0484_ _0485_ VPWR VGND sg13g2_and2_1
XFILLER_3_939 VPWR VGND sg13g2_decap_8
XFILLER_49_35 VPWR VGND sg13g2_decap_4
Xfanout720 net721 net720 VPWR VGND sg13g2_buf_8
Xfanout731 _1577_ net731 VPWR VGND sg13g2_buf_8
Xfanout742 _1510_ net742 VPWR VGND sg13g2_buf_8
Xfanout753 _1588_ net753 VPWR VGND sg13g2_buf_8
Xfanout764 _1519_ net764 VPWR VGND sg13g2_buf_8
Xfanout775 sap_3_inst.controller.opcode\[4\] net775 VPWR VGND sg13g2_buf_8
XFILLER_46_604 VPWR VGND sg13g2_decap_8
Xfanout786 sap_3_inst.controller.opcode\[0\] net786 VPWR VGND sg13g2_buf_8
XFILLER_19_829 VPWR VGND sg13g2_decap_8
Xfanout797 sap_3_inst.alu.acc\[4\] net797 VPWR VGND sg13g2_buf_8
XFILLER_27_840 VPWR VGND sg13g2_decap_8
XFILLER_42_821 VPWR VGND sg13g2_decap_8
XFILLER_41_342 VPWR VGND sg13g2_fill_1
XFILLER_14_534 VPWR VGND sg13g2_decap_8
XFILLER_26_394 VPWR VGND sg13g2_decap_8
XFILLER_42_898 VPWR VGND sg13g2_decap_8
XFILLER_6_733 VPWR VGND sg13g2_decap_8
XFILLER_10_795 VPWR VGND sg13g2_decap_8
XFILLER_2_994 VPWR VGND sg13g2_decap_8
XFILLER_49_442 VPWR VGND sg13g2_decap_8
XFILLER_1_493 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
XFILLER_37_604 VPWR VGND sg13g2_decap_8
XFILLER_18_840 VPWR VGND sg13g2_decap_8
X_3901_ net811 net55 _1332_ _0162_ VPWR VGND sg13g2_a21o_1
XFILLER_33_854 VPWR VGND sg13g2_decap_8
X_3832_ VGND VPWR net610 _1032_ _1273_ net605 sg13g2_a21oi_1
XFILLER_9_560 VPWR VGND sg13g2_decap_8
X_3763_ _1225_ net660 _0910_ VPWR VGND sg13g2_nand2_1
X_3694_ net578 _1178_ _1179_ _1180_ VPWR VGND sg13g2_nor3_1
X_2714_ _0288_ net576 _1899_ VPWR VGND sg13g2_nand2_2
X_2645_ _0232_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] net643
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2576_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[2\] net648 _1986_ VPWR
+ VGND sg13g2_nor2_1
X_4177_ net833 VGND VPWR _0141_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\]
+ clknet_5_18__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3128_ net729 _0655_ net778 _0656_ VPWR VGND sg13g2_nand3_1
XFILLER_28_637 VPWR VGND sg13g2_decap_8
X_3059_ sap_3_inst.alu.tmp\[5\] net22 net715 _0055_ VPWR VGND sg13g2_mux2_1
XFILLER_24_832 VPWR VGND sg13g2_decap_8
XFILLER_23_386 VPWR VGND sg13g2_decap_8
XFILLER_11_559 VPWR VGND sg13g2_decap_8
XFILLER_13_1026 VPWR VGND sg13g2_fill_2
XFILLER_3_736 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
Xfanout583 _1390_ net583 VPWR VGND sg13g2_buf_8
Xfanout572 _1982_ net572 VPWR VGND sg13g2_buf_8
XFILLER_47_935 VPWR VGND sg13g2_decap_8
XFILLER_46_401 VPWR VGND sg13g2_decap_8
XFILLER_19_626 VPWR VGND sg13g2_decap_8
Xfanout594 _1208_ net594 VPWR VGND sg13g2_buf_8
XFILLER_18_147 VPWR VGND sg13g2_fill_2
XFILLER_46_478 VPWR VGND sg13g2_decap_8
XFILLER_15_854 VPWR VGND sg13g2_decap_8
XFILLER_33_128 VPWR VGND sg13g2_fill_2
XFILLER_42_695 VPWR VGND sg13g2_decap_8
XFILLER_30_835 VPWR VGND sg13g2_decap_8
XFILLER_6_530 VPWR VGND sg13g2_decap_8
XFILLER_10_592 VPWR VGND sg13g2_decap_8
X_2430_ _1850_ _1569_ _1576_ VPWR VGND sg13g2_nand2_1
XFILLER_29_1000 VPWR VGND sg13g2_decap_8
X_2361_ _1781_ _1520_ _1780_ VPWR VGND sg13g2_nand2_1
XFILLER_2_791 VPWR VGND sg13g2_decap_8
X_2292_ _1515_ VPWR _1712_ VGND _1584_ _1591_ sg13g2_o21ai_1
X_4100_ net818 VGND VPWR _0064_ sap_3_inst.controller.opcode\[6\] clknet_5_4__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_2_52 VPWR VGND sg13g2_fill_2
X_4031_ VPWR _0192_ _1433_ VGND sg13g2_inv_1
XFILLER_38_968 VPWR VGND sg13g2_decap_8
XFILLER_37_478 VPWR VGND sg13g2_decap_8
XFILLER_24_128 VPWR VGND sg13g2_fill_1
XFILLER_21_802 VPWR VGND sg13g2_decap_8
XFILLER_33_651 VPWR VGND sg13g2_decap_8
XFILLER_36_1004 VPWR VGND sg13g2_decap_8
XFILLER_32_183 VPWR VGND sg13g2_fill_2
X_3815_ _1262_ VPWR _0146_ VGND _1469_ net658 sg13g2_o21ai_1
XFILLER_20_356 VPWR VGND sg13g2_fill_2
XFILLER_21_879 VPWR VGND sg13g2_decap_8
X_3746_ _1212_ _1064_ _1065_ VPWR VGND sg13g2_nand2_1
X_3677_ _1166_ VPWR _1167_ VGND net599 _1014_ sg13g2_o21ai_1
X_2628_ _0217_ net629 _0216_ VPWR VGND sg13g2_nand2_1
XFILLER_0_717 VPWR VGND sg13g2_decap_8
X_2559_ _1971_ _1970_ _1723_ VPWR VGND sg13g2_nand2b_1
XFILLER_43_1008 VPWR VGND sg13g2_decap_8
XFILLER_29_902 VPWR VGND sg13g2_decap_8
X_4229_ net844 VGND VPWR _0192_ sap_3_inst.reg_file.array_serializer_inst.word_index\[3\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_29_979 VPWR VGND sg13g2_decap_8
XFILLER_43_448 VPWR VGND sg13g2_decap_8
XFILLER_8_817 VPWR VGND sg13g2_decap_8
XFILLER_12_868 VPWR VGND sg13g2_decap_8
XFILLER_11_389 VPWR VGND sg13g2_fill_1
XFILLER_3_533 VPWR VGND sg13g2_decap_8
XFILLER_47_732 VPWR VGND sg13g2_decap_8
XFILLER_19_423 VPWR VGND sg13g2_fill_1
XFILLER_35_927 VPWR VGND sg13g2_decap_8
XFILLER_15_651 VPWR VGND sg13g2_decap_8
XFILLER_30_632 VPWR VGND sg13g2_decap_8
XFILLER_42_492 VPWR VGND sg13g2_decap_8
X_3600_ VPWR VGND _1106_ net618 _1105_ net606 _1107_ _0993_ sg13g2_a221oi_1
X_3531_ net605 _0898_ _1050_ VPWR VGND sg13g2_nor2_1
XFILLER_7_894 VPWR VGND sg13g2_decap_8
X_3462_ _0985_ _0869_ _0984_ net595 net22 VPWR VGND sg13g2_a22oi_1
X_2413_ net740 _1676_ _1833_ VPWR VGND sg13g2_nor2_1
X_3393_ VGND VPWR _0835_ _0918_ _0919_ _0917_ sg13g2_a21oi_1
X_2344_ _1762_ VPWR _1764_ VGND net766 _1521_ sg13g2_o21ai_1
X_2275_ VGND VPWR _1606_ _1680_ _1695_ _1694_ sg13g2_a21oi_1
X_4014_ _1419_ VPWR _1422_ VGND u_ser.bit_pos\[1\] _1421_ sg13g2_o21ai_1
XFILLER_26_905 VPWR VGND sg13g2_decap_8
XFILLER_38_765 VPWR VGND sg13g2_decap_8
XFILLER_19_990 VPWR VGND sg13g2_decap_8
XFILLER_20_153 VPWR VGND sg13g2_decap_4
XFILLER_21_676 VPWR VGND sg13g2_decap_8
X_3729_ _1204_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] net617 VPWR
+ VGND sg13g2_nand2_1
XFILLER_0_514 VPWR VGND sg13g2_decap_8
XFILLER_48_507 VPWR VGND sg13g2_decap_8
XFILLER_29_776 VPWR VGND sg13g2_decap_8
XFILLER_44_757 VPWR VGND sg13g2_decap_8
XFILLER_17_949 VPWR VGND sg13g2_decap_8
XFILLER_25_960 VPWR VGND sg13g2_decap_8
XFILLER_43_278 VPWR VGND sg13g2_fill_2
XFILLER_40_996 VPWR VGND sg13g2_decap_8
XFILLER_8_614 VPWR VGND sg13g2_decap_8
XFILLER_12_665 VPWR VGND sg13g2_decap_8
XFILLER_11_175 VPWR VGND sg13g2_fill_1
XFILLER_4_886 VPWR VGND sg13g2_decap_8
XFILLER_26_1003 VPWR VGND sg13g2_decap_8
X_2060_ VPWR _1482_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] VGND
+ sg13g2_inv_1
XFILLER_35_724 VPWR VGND sg13g2_decap_8
X_2962_ net790 _0324_ _0517_ VPWR VGND sg13g2_nor2_1
XFILLER_31_941 VPWR VGND sg13g2_decap_8
X_2893_ _1460_ _1473_ _0450_ VPWR VGND sg13g2_nor2_1
XFILLER_7_691 VPWR VGND sg13g2_decap_8
X_3514_ _0827_ _1034_ net621 _1035_ VPWR VGND sg13g2_nand3_1
X_3445_ _0966_ _0968_ _0960_ _0969_ VPWR VGND sg13g2_nand3_1
X_3376_ _0902_ net663 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] net666
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2327_ net740 _1746_ _1747_ VPWR VGND sg13g2_nor2_1
X_2258_ _1678_ net758 net754 VPWR VGND sg13g2_nand2_2
XFILLER_26_702 VPWR VGND sg13g2_decap_8
XFILLER_38_562 VPWR VGND sg13g2_decap_8
X_2189_ _1525_ _1562_ net781 _1609_ VPWR VGND sg13g2_nand3_1
XFILLER_25_201 VPWR VGND sg13g2_fill_1
XFILLER_14_919 VPWR VGND sg13g2_decap_8
XFILLER_26_779 VPWR VGND sg13g2_decap_8
XFILLER_43_37 VPWR VGND sg13g2_fill_2
XFILLER_41_749 VPWR VGND sg13g2_decap_8
XFILLER_13_418 VPWR VGND sg13g2_fill_2
XFILLER_22_930 VPWR VGND sg13g2_decap_8
XFILLER_40_259 VPWR VGND sg13g2_fill_1
XFILLER_21_451 VPWR VGND sg13g2_fill_1
XFILLER_1_801 VPWR VGND sg13g2_decap_8
XFILLER_1_878 VPWR VGND sg13g2_decap_8
XFILLER_49_827 VPWR VGND sg13g2_decap_8
XFILLER_48_304 VPWR VGND sg13g2_decap_8
XFILLER_29_573 VPWR VGND sg13g2_decap_8
XFILLER_17_746 VPWR VGND sg13g2_decap_8
XFILLER_44_554 VPWR VGND sg13g2_decap_8
XFILLER_32_727 VPWR VGND sg13g2_decap_8
XFILLER_13_963 VPWR VGND sg13g2_decap_8
XFILLER_9_945 VPWR VGND sg13g2_decap_8
XFILLER_40_793 VPWR VGND sg13g2_decap_8
XFILLER_8_488 VPWR VGND sg13g2_decap_8
XFILLER_4_683 VPWR VGND sg13g2_decap_8
X_3230_ net701 net692 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] _0758_
+ VPWR VGND net687 sg13g2_nand4_1
X_3161_ _0659_ net686 _0689_ VPWR VGND sg13g2_and2_1
X_2112_ net760 net761 _1532_ VPWR VGND sg13g2_nor2b_2
XFILLER_39_337 VPWR VGND sg13g2_fill_1
XFILLER_48_871 VPWR VGND sg13g2_decap_8
X_3092_ _1442_ net773 _1570_ net731 _0620_ VPWR VGND sg13g2_nor4_1
X_2043_ VPWR _1465_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] VGND
+ sg13g2_inv_1
XFILLER_35_521 VPWR VGND sg13g2_decap_8
XFILLER_22_215 VPWR VGND sg13g2_fill_2
XFILLER_35_598 VPWR VGND sg13g2_decap_8
X_3994_ _1406_ sap_3_inst.alu.act\[5\] net583 VPWR VGND sg13g2_nand2_1
X_2945_ _0496_ VPWR _0501_ VGND net625 _0500_ sg13g2_o21ai_1
Xclkbuf_4_9_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_9_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2876_ _0434_ _0423_ _0432_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_609 VPWR VGND sg13g2_decap_8
X_3428_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] _0951_
+ net663 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] _0952_ net666 sg13g2_a221oi_1
X_3359_ _0886_ _0807_ _0884_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_716 VPWR VGND sg13g2_decap_8
XFILLER_26_576 VPWR VGND sg13g2_decap_8
XFILLER_41_546 VPWR VGND sg13g2_decap_8
XFILLER_10_900 VPWR VGND sg13g2_decap_8
XFILLER_6_915 VPWR VGND sg13g2_decap_8
XFILLER_10_977 VPWR VGND sg13g2_decap_8
XFILLER_49_624 VPWR VGND sg13g2_decap_8
XFILLER_1_675 VPWR VGND sg13g2_decap_8
XFILLER_45_830 VPWR VGND sg13g2_decap_8
XFILLER_17_543 VPWR VGND sg13g2_decap_8
XFILLER_32_524 VPWR VGND sg13g2_decap_8
XFILLER_13_760 VPWR VGND sg13g2_decap_8
XFILLER_40_590 VPWR VGND sg13g2_decap_8
X_2730_ u_ser.state\[1\] u_ser.state\[0\] _0185_ VPWR VGND sg13g2_nor2_2
XFILLER_9_742 VPWR VGND sg13g2_decap_8
X_2661_ _0245_ _0246_ _0244_ _0248_ VPWR VGND _0247_ sg13g2_nand4_1
XFILLER_8_241 VPWR VGND sg13g2_fill_1
X_2592_ _2002_ net636 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] net646
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_4_480 VPWR VGND sg13g2_decap_8
X_3213_ _0734_ _0735_ _0738_ _0740_ _0741_ VPWR VGND sg13g2_and4_1
X_4193_ net847 VGND VPWR net57 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\]
+ clknet_3_6__leaf_clk sg13g2_dfrbpq_2
X_3144_ _1608_ VPWR _0672_ VGND _1632_ _0671_ sg13g2_o21ai_1
XFILLER_28_819 VPWR VGND sg13g2_decap_8
X_3075_ VGND VPWR _1615_ _1749_ _0603_ net731 sg13g2_a21oi_1
X_2026_ VPWR _1448_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_36_885 VPWR VGND sg13g2_decap_8
XFILLER_39_1013 VPWR VGND sg13g2_decap_8
X_3977_ _1393_ VPWR _0177_ VGND net582 _1392_ sg13g2_o21ai_1
XFILLER_23_568 VPWR VGND sg13g2_decap_8
X_2928_ VGND VPWR _0484_ sap_3_inst.alu.tmp\[5\] net794 sg13g2_or2_1
X_2859_ VGND VPWR _0412_ _0415_ _0417_ _0416_ sg13g2_a21oi_1
XFILLER_3_918 VPWR VGND sg13g2_decap_8
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_1017 VPWR VGND sg13g2_decap_8
XFILLER_6_8 VPWR VGND sg13g2_decap_8
Xfanout721 _1953_ net721 VPWR VGND sg13g2_buf_8
Xfanout710 _1389_ net710 VPWR VGND sg13g2_buf_8
Xfanout732 _1572_ net732 VPWR VGND sg13g2_buf_8
Xfanout754 _1557_ net754 VPWR VGND sg13g2_buf_8
Xfanout743 net744 net743 VPWR VGND sg13g2_buf_8
Xfanout765 _1518_ net765 VPWR VGND sg13g2_buf_8
Xfanout776 net779 net776 VPWR VGND sg13g2_buf_8
Xfanout787 net788 net787 VPWR VGND sg13g2_buf_2
Xfanout798 net800 net798 VPWR VGND sg13g2_buf_8
XFILLER_19_808 VPWR VGND sg13g2_decap_8
XFILLER_42_800 VPWR VGND sg13g2_decap_8
XFILLER_14_513 VPWR VGND sg13g2_decap_8
XFILLER_27_896 VPWR VGND sg13g2_decap_8
XFILLER_42_877 VPWR VGND sg13g2_decap_8
XFILLER_6_712 VPWR VGND sg13g2_decap_8
XFILLER_5_200 VPWR VGND sg13g2_fill_1
XFILLER_10_774 VPWR VGND sg13g2_decap_8
XFILLER_6_789 VPWR VGND sg13g2_decap_8
XFILLER_2_973 VPWR VGND sg13g2_decap_8
XFILLER_49_421 VPWR VGND sg13g2_decap_8
XFILLER_1_472 VPWR VGND sg13g2_decap_8
XFILLER_49_498 VPWR VGND sg13g2_decap_8
XFILLER_18_896 VPWR VGND sg13g2_decap_8
X_3900_ VPWR VGND _1331_ net812 _1326_ _1461_ _1332_ net807 sg13g2_a221oi_1
XFILLER_32_332 VPWR VGND sg13g2_fill_1
XFILLER_33_833 VPWR VGND sg13g2_decap_8
X_3831_ _1272_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] net610 VPWR
+ VGND sg13g2_nand2_1
XFILLER_20_549 VPWR VGND sg13g2_decap_8
X_3762_ _1224_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] net611 VPWR
+ VGND sg13g2_nand2_1
XFILLER_32_387 VPWR VGND sg13g2_fill_2
X_3693_ VGND VPWR _0666_ _0911_ _1179_ net598 sg13g2_a21oi_1
X_2713_ net577 _1919_ net13 VPWR VGND sg13g2_and2_1
X_2644_ _0231_ sap_3_inst.alu.flags\[0\] _0230_ VPWR VGND sg13g2_nand2_1
X_2575_ _1985_ sap_3_inst.alu.flags\[2\] _1961_ VPWR VGND sg13g2_nand2_1
X_4176_ net841 VGND VPWR _0140_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\]
+ clknet_5_28__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_616 VPWR VGND sg13g2_decap_8
X_3127_ net769 net767 _1518_ _0655_ VPWR VGND sg13g2_nor3_1
X_3058_ _0597_ VPWR _0054_ VGND _1473_ net716 sg13g2_o21ai_1
XFILLER_24_811 VPWR VGND sg13g2_decap_8
XFILLER_36_682 VPWR VGND sg13g2_decap_8
XFILLER_24_888 VPWR VGND sg13g2_decap_8
XFILLER_11_538 VPWR VGND sg13g2_decap_8
XFILLER_7_509 VPWR VGND sg13g2_decap_8
XFILLER_13_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_715 VPWR VGND sg13g2_decap_8
XFILLER_47_914 VPWR VGND sg13g2_decap_8
Xfanout584 net585 net584 VPWR VGND sg13g2_buf_8
XFILLER_19_605 VPWR VGND sg13g2_decap_8
Xfanout573 net573 net22 VPWR VGND sg13g2_buf_8
XFILLER_18_115 VPWR VGND sg13g2_fill_2
Xfanout595 net596 net595 VPWR VGND sg13g2_buf_8
XFILLER_46_457 VPWR VGND sg13g2_decap_8
XFILLER_34_619 VPWR VGND sg13g2_decap_8
XFILLER_15_833 VPWR VGND sg13g2_decap_8
XFILLER_27_693 VPWR VGND sg13g2_decap_8
XFILLER_42_674 VPWR VGND sg13g2_decap_8
XFILLER_30_814 VPWR VGND sg13g2_decap_8
XFILLER_10_571 VPWR VGND sg13g2_decap_8
XFILLER_6_586 VPWR VGND sg13g2_decap_8
X_2360_ _1676_ net729 net783 _1780_ VPWR VGND sg13g2_nand3_1
XFILLER_2_770 VPWR VGND sg13g2_decap_8
X_2291_ _1584_ _1591_ _1711_ VPWR VGND sg13g2_nor2_1
XFILLER_2_31 VPWR VGND sg13g2_decap_8
X_4030_ _1433_ _1430_ net815 _1429_ net810 VPWR VGND sg13g2_a22oi_1
XFILLER_38_947 VPWR VGND sg13g2_decap_8
XFILLER_49_295 VPWR VGND sg13g2_decap_8
XFILLER_18_693 VPWR VGND sg13g2_decap_8
XFILLER_33_630 VPWR VGND sg13g2_decap_8
XFILLER_21_858 VPWR VGND sg13g2_decap_8
X_3814_ _1261_ VPWR _1262_ VGND _0874_ _1260_ sg13g2_o21ai_1
X_3745_ _1211_ VPWR _0127_ VGND _1192_ net593 sg13g2_o21ai_1
XFILLER_9_380 VPWR VGND sg13g2_fill_1
X_3676_ net624 _1165_ _1166_ VPWR VGND sg13g2_nor2_1
X_2627_ _0216_ net762 _1839_ VPWR VGND sg13g2_nand2_1
X_2558_ _1970_ _1966_ _1969_ net649 _1446_ VPWR VGND sg13g2_a22oi_1
X_2489_ _1905_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] net645
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4228_ net844 VGND VPWR _0191_ sap_3_inst.reg_file.array_serializer_inst.word_index\[2\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
X_4159_ net820 VGND VPWR _0123_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\]
+ clknet_5_6__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_958 VPWR VGND sg13g2_decap_8
XFILLER_44_939 VPWR VGND sg13g2_decap_8
XFILLER_16_619 VPWR VGND sg13g2_decap_8
XFILLER_43_427 VPWR VGND sg13g2_decap_8
XFILLER_15_118 VPWR VGND sg13g2_decap_4
XFILLER_11_313 VPWR VGND sg13g2_fill_1
XFILLER_12_847 VPWR VGND sg13g2_decap_8
XFILLER_24_685 VPWR VGND sg13g2_decap_8
XFILLER_3_512 VPWR VGND sg13g2_decap_8
XFILLER_3_589 VPWR VGND sg13g2_decap_8
XFILLER_47_711 VPWR VGND sg13g2_decap_8
XFILLER_35_906 VPWR VGND sg13g2_decap_8
XFILLER_47_788 VPWR VGND sg13g2_decap_8
XFILLER_28_980 VPWR VGND sg13g2_decap_8
XFILLER_15_630 VPWR VGND sg13g2_decap_8
XFILLER_27_490 VPWR VGND sg13g2_decap_8
XFILLER_43_994 VPWR VGND sg13g2_decap_8
XFILLER_42_471 VPWR VGND sg13g2_decap_8
XFILLER_30_611 VPWR VGND sg13g2_decap_8
XFILLER_30_688 VPWR VGND sg13g2_decap_8
X_3530_ VGND VPWR net600 _0898_ _1049_ net584 sg13g2_a21oi_1
XFILLER_7_873 VPWR VGND sg13g2_decap_8
X_3461_ _0984_ _0288_ net597 VPWR VGND sg13g2_nand2_1
X_2412_ _1831_ VPWR _1832_ VGND _1551_ _1823_ sg13g2_o21ai_1
X_3392_ _0800_ _0873_ _0918_ VPWR VGND sg13g2_nor2_1
X_2343_ _1761_ _1762_ _1530_ _1763_ VPWR VGND sg13g2_nand3_1
X_2274_ _1689_ _1693_ _1684_ _1694_ VPWR VGND sg13g2_nand3_1
X_4013_ _1420_ VPWR _1421_ VGND u_ser.bit_pos\[0\] u_ser.shadow_reg\[5\] sg13g2_o21ai_1
XFILLER_38_744 VPWR VGND sg13g2_decap_8
XFILLER_25_449 VPWR VGND sg13g2_decap_8
XFILLER_18_490 VPWR VGND sg13g2_decap_8
XFILLER_34_983 VPWR VGND sg13g2_decap_8
XFILLER_21_655 VPWR VGND sg13g2_decap_8
XFILLER_32_28 VPWR VGND sg13g2_fill_1
XFILLER_10_1019 VPWR VGND sg13g2_decap_8
X_3728_ _0118_ _1099_ _1203_ net616 _1478_ VPWR VGND sg13g2_a22oi_1
X_3659_ _1152_ _1149_ _0287_ net684 net572 VPWR VGND sg13g2_a22oi_1
XFILLER_29_755 VPWR VGND sg13g2_decap_8
XFILLER_17_928 VPWR VGND sg13g2_decap_8
XFILLER_44_736 VPWR VGND sg13g2_decap_8
XFILLER_43_202 VPWR VGND sg13g2_fill_1
XFILLER_19_1011 VPWR VGND sg13g2_decap_8
XFILLER_32_909 VPWR VGND sg13g2_decap_8
XFILLER_12_644 VPWR VGND sg13g2_decap_8
XFILLER_24_482 VPWR VGND sg13g2_decap_8
XFILLER_40_975 VPWR VGND sg13g2_decap_8
XFILLER_4_865 VPWR VGND sg13g2_decap_8
XFILLER_35_703 VPWR VGND sg13g2_decap_8
XFILLER_47_585 VPWR VGND sg13g2_decap_8
XFILLER_34_246 VPWR VGND sg13g2_fill_1
X_2961_ _0497_ _0515_ _0516_ VPWR VGND sg13g2_nor2_1
XFILLER_16_983 VPWR VGND sg13g2_decap_8
XFILLER_31_920 VPWR VGND sg13g2_decap_8
XFILLER_34_268 VPWR VGND sg13g2_fill_1
XFILLER_43_791 VPWR VGND sg13g2_decap_8
XFILLER_33_1008 VPWR VGND sg13g2_decap_8
X_2892_ net714 VPWR _0449_ VGND _0446_ _0447_ sg13g2_o21ai_1
XFILLER_31_997 VPWR VGND sg13g2_decap_8
XFILLER_30_485 VPWR VGND sg13g2_decap_8
XFILLER_7_670 VPWR VGND sg13g2_decap_8
X_3513_ _1034_ _0722_ _0840_ VPWR VGND sg13g2_xnor2_1
X_3444_ _0967_ VPWR _0968_ VGND net13 net596 sg13g2_o21ai_1
XFILLER_40_0 VPWR VGND sg13g2_fill_2
X_3375_ _0901_ net661 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] net676
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2326_ net773 VPWR _1746_ VGND _1441_ _1442_ sg13g2_o21ai_1
X_2257_ _1504_ _1558_ _1677_ VPWR VGND sg13g2_nor2_2
XFILLER_38_541 VPWR VGND sg13g2_decap_8
X_2188_ net785 net782 _1564_ _1608_ VPWR VGND sg13g2_nor3_2
XFILLER_26_758 VPWR VGND sg13g2_decap_8
XFILLER_41_728 VPWR VGND sg13g2_decap_8
XFILLER_34_780 VPWR VGND sg13g2_decap_8
XFILLER_22_986 VPWR VGND sg13g2_decap_8
XFILLER_49_806 VPWR VGND sg13g2_decap_8
XFILLER_1_857 VPWR VGND sg13g2_decap_8
XFILLER_29_552 VPWR VGND sg13g2_decap_8
XFILLER_44_533 VPWR VGND sg13g2_decap_8
XFILLER_17_725 VPWR VGND sg13g2_decap_8
XFILLER_32_706 VPWR VGND sg13g2_decap_8
XFILLER_13_942 VPWR VGND sg13g2_decap_8
XFILLER_24_290 VPWR VGND sg13g2_fill_1
XFILLER_40_772 VPWR VGND sg13g2_decap_8
XFILLER_9_924 VPWR VGND sg13g2_decap_8
XFILLER_12_474 VPWR VGND sg13g2_fill_1
XFILLER_4_662 VPWR VGND sg13g2_decap_8
X_3160_ VPWR VGND _0686_ _0684_ _0685_ _0617_ _0688_ _0618_ sg13g2_a221oi_1
X_2111_ _1529_ VPWR _1531_ VGND net767 net756 sg13g2_o21ai_1
X_3091_ _0617_ _0618_ _0619_ VPWR VGND sg13g2_and2_1
Xhold1 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[4\] VPWR VGND net50 sg13g2_dlygate4sd3_1
XFILLER_48_850 VPWR VGND sg13g2_decap_8
X_2042_ VPWR _1464_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] VGND
+ sg13g2_inv_1
XFILLER_47_382 VPWR VGND sg13g2_decap_8
XFILLER_35_500 VPWR VGND sg13g2_decap_8
XFILLER_35_577 VPWR VGND sg13g2_decap_8
X_3993_ _1405_ VPWR _0181_ VGND net583 _1404_ sg13g2_o21ai_1
XFILLER_16_780 VPWR VGND sg13g2_decap_8
X_2944_ _0326_ _0464_ _0500_ VPWR VGND sg13g2_and2_1
X_2875_ _0422_ _0432_ _0433_ VPWR VGND sg13g2_nor2_1
XFILLER_30_271 VPWR VGND sg13g2_fill_2
XFILLER_31_794 VPWR VGND sg13g2_decap_8
X_3427_ _0951_ _0947_ _0950_ VPWR VGND sg13g2_nand2_1
X_3358_ _0710_ _0722_ _0805_ _0885_ VGND VPWR _0883_ sg13g2_nor4_2
X_2309_ _1729_ _1534_ _1642_ VPWR VGND sg13g2_nand2_1
X_3289_ VPWR VGND _0812_ _0815_ _1703_ _1613_ _0817_ _1697_ sg13g2_a221oi_1
XFILLER_39_894 VPWR VGND sg13g2_decap_8
XFILLER_26_555 VPWR VGND sg13g2_decap_8
XFILLER_41_525 VPWR VGND sg13g2_decap_8
XFILLER_16_1025 VPWR VGND sg13g2_decap_4
XFILLER_22_783 VPWR VGND sg13g2_decap_8
XFILLER_10_956 VPWR VGND sg13g2_decap_8
XFILLER_49_603 VPWR VGND sg13g2_decap_8
XFILLER_1_654 VPWR VGND sg13g2_decap_8
XFILLER_17_522 VPWR VGND sg13g2_decap_8
XFILLER_36_319 VPWR VGND sg13g2_fill_2
XFILLER_45_886 VPWR VGND sg13g2_decap_8
XFILLER_32_503 VPWR VGND sg13g2_decap_8
XFILLER_17_599 VPWR VGND sg13g2_decap_8
XFILLER_9_721 VPWR VGND sg13g2_decap_8
X_2660_ _0247_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] net647
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_9_798 VPWR VGND sg13g2_decap_8
X_2591_ _2001_ net635 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] net649
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] VPWR VGND sg13g2_a22oi_1
X_3212_ _0740_ _0736_ _0737_ _0739_ VPWR VGND sg13g2_and3_1
X_4192_ net847 VGND VPWR _0156_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[0\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
X_3143_ _1536_ _1642_ _0671_ VPWR VGND sg13g2_and2_1
X_3074_ VGND VPWR _1443_ net739 _0065_ _0602_ sg13g2_a21oi_1
X_2025_ VPWR _1447_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_36_864 VPWR VGND sg13g2_decap_8
XFILLER_23_547 VPWR VGND sg13g2_decap_8
X_3976_ _1393_ sap_3_inst.alu.act\[0\] net582 VPWR VGND sg13g2_nand2_1
XFILLER_10_208 VPWR VGND sg13g2_fill_1
X_2927_ net794 sap_3_inst.alu.tmp\[5\] _0483_ VPWR VGND sg13g2_nor2_1
XFILLER_31_591 VPWR VGND sg13g2_decap_8
X_2858_ net714 VPWR _0416_ VGND _0412_ _0415_ sg13g2_o21ai_1
X_2789_ _0346_ VPWR _0350_ VGND net805 _0325_ sg13g2_o21ai_1
XFILLER_2_429 VPWR VGND sg13g2_fill_2
Xfanout700 _0645_ net700 VPWR VGND sg13g2_buf_8
Xfanout733 _1572_ net733 VPWR VGND sg13g2_buf_1
Xfanout711 _0827_ net711 VPWR VGND sg13g2_buf_8
Xfanout722 net723 net722 VPWR VGND sg13g2_buf_8
Xfanout755 _1532_ net755 VPWR VGND sg13g2_buf_8
Xfanout744 net745 net744 VPWR VGND sg13g2_buf_8
Xfanout766 net767 net766 VPWR VGND sg13g2_buf_8
Xfanout777 net779 net777 VPWR VGND sg13g2_buf_8
Xfanout788 net789 net788 VPWR VGND sg13g2_buf_2
Xfanout799 net800 net799 VPWR VGND sg13g2_buf_1
XFILLER_46_639 VPWR VGND sg13g2_decap_8
XFILLER_39_691 VPWR VGND sg13g2_decap_8
XFILLER_27_875 VPWR VGND sg13g2_decap_8
Xclkbuf_5_29__f_sap_3_inst.alu.clk_regs clknet_4_14_0_sap_3_inst.alu.clk_regs clknet_5_29__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_42_856 VPWR VGND sg13g2_decap_8
XFILLER_41_355 VPWR VGND sg13g2_fill_2
XFILLER_14_569 VPWR VGND sg13g2_decap_8
XFILLER_22_580 VPWR VGND sg13g2_decap_8
XFILLER_10_753 VPWR VGND sg13g2_decap_8
XFILLER_6_768 VPWR VGND sg13g2_decap_8
XFILLER_2_952 VPWR VGND sg13g2_decap_8
XFILLER_49_400 VPWR VGND sg13g2_decap_8
XFILLER_49_477 VPWR VGND sg13g2_decap_8
XFILLER_37_639 VPWR VGND sg13g2_decap_8
XFILLER_18_875 VPWR VGND sg13g2_decap_8
XFILLER_33_812 VPWR VGND sg13g2_decap_8
XFILLER_45_683 VPWR VGND sg13g2_decap_8
X_3830_ _0152_ _1110_ _1271_ net610 _1485_ VPWR VGND sg13g2_a22oi_1
XFILLER_33_889 VPWR VGND sg13g2_decap_8
XFILLER_20_528 VPWR VGND sg13g2_decap_8
X_3761_ net611 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] _1223_ _0131_
+ VPWR VGND sg13g2_a21o_1
X_2712_ VPWR net12 _0287_ VGND sg13g2_inv_1
XFILLER_9_595 VPWR VGND sg13g2_decap_8
X_3692_ net604 _0922_ _1052_ _1178_ VPWR VGND sg13g2_nor3_1
X_2643_ _0230_ _1946_ _1786_ VPWR VGND sg13g2_nand2b_1
X_2574_ _1962_ VPWR _0028_ VGND _1961_ _1984_ sg13g2_o21ai_1
X_4175_ net820 VGND VPWR _0139_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\]
+ clknet_5_6__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3126_ net757 VPWR _0654_ VGND _0647_ _0653_ sg13g2_o21ai_1
XFILLER_43_609 VPWR VGND sg13g2_decap_8
X_3057_ _0597_ net32 net716 VPWR VGND sg13g2_nand2_1
XFILLER_36_661 VPWR VGND sg13g2_decap_8
XFILLER_24_867 VPWR VGND sg13g2_decap_8
XFILLER_11_517 VPWR VGND sg13g2_decap_8
X_3959_ _1125_ _1126_ net655 _1383_ VPWR VGND sg13g2_nand3_1
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
Xfanout574 _0334_ net574 VPWR VGND sg13g2_buf_8
Xfanout585 _1044_ net585 VPWR VGND sg13g2_buf_8
Xfanout596 _0868_ net596 VPWR VGND sg13g2_buf_8
XFILLER_46_436 VPWR VGND sg13g2_decap_8
XFILLER_18_127 VPWR VGND sg13g2_fill_2
XFILLER_15_812 VPWR VGND sg13g2_decap_8
XFILLER_27_672 VPWR VGND sg13g2_decap_8
XFILLER_42_653 VPWR VGND sg13g2_decap_8
XFILLER_15_889 VPWR VGND sg13g2_decap_8
XFILLER_10_550 VPWR VGND sg13g2_decap_8
XFILLER_6_565 VPWR VGND sg13g2_decap_8
X_2290_ _1709_ VPWR _1710_ VGND _1607_ _1695_ sg13g2_o21ai_1
XFILLER_49_274 VPWR VGND sg13g2_decap_8
XFILLER_2_54 VPWR VGND sg13g2_fill_1
XFILLER_38_926 VPWR VGND sg13g2_decap_8
XFILLER_18_672 VPWR VGND sg13g2_decap_8
XFILLER_45_480 VPWR VGND sg13g2_decap_8
XFILLER_17_160 VPWR VGND sg13g2_fill_1
XFILLER_21_837 VPWR VGND sg13g2_decap_8
XFILLER_33_686 VPWR VGND sg13g2_decap_8
X_3813_ net609 _1083_ _1261_ VPWR VGND sg13g2_nor2_1
X_3744_ _1211_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] net593 VPWR
+ VGND sg13g2_nand2_1
X_3675_ VPWR VGND net15 _0850_ _1137_ net33 _1165_ net684 sg13g2_a221oi_1
X_2626_ VGND VPWR _0215_ net629 net803 sg13g2_or2_1
X_2557_ net648 _1964_ _1967_ _1968_ _1969_ VPWR VGND sg13g2_and4_1
X_2488_ _1904_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] net650
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4227_ net844 VGND VPWR _0190_ sap_3_inst.reg_file.array_serializer_inst.word_index\[1\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_2
XFILLER_29_937 VPWR VGND sg13g2_decap_8
X_4158_ net843 VGND VPWR _0122_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\]
+ clknet_5_27__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_44_918 VPWR VGND sg13g2_decap_8
XFILLER_43_406 VPWR VGND sg13g2_decap_8
X_3109_ net741 _1515_ _1715_ _0637_ VPWR VGND sg13g2_nor3_1
X_4089_ net838 VGND VPWR _0053_ sap_3_inst.alu.tmp\[3\] clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_28_469 VPWR VGND sg13g2_decap_8
XFILLER_24_664 VPWR VGND sg13g2_decap_8
XFILLER_12_826 VPWR VGND sg13g2_decap_8
XFILLER_23_141 VPWR VGND sg13g2_fill_1
XFILLER_11_336 VPWR VGND sg13g2_fill_1
XFILLER_20_892 VPWR VGND sg13g2_decap_8
XFILLER_11_41 VPWR VGND sg13g2_fill_1
XFILLER_3_568 VPWR VGND sg13g2_decap_8
XFILLER_4_1026 VPWR VGND sg13g2_fill_2
XFILLER_47_767 VPWR VGND sg13g2_decap_8
XFILLER_43_973 VPWR VGND sg13g2_decap_8
XFILLER_42_450 VPWR VGND sg13g2_decap_8
XFILLER_15_686 VPWR VGND sg13g2_decap_8
XFILLER_30_667 VPWR VGND sg13g2_decap_8
XFILLER_7_852 VPWR VGND sg13g2_decap_8
XFILLER_11_881 VPWR VGND sg13g2_decap_8
X_3460_ VGND VPWR net669 _0980_ _0983_ _0982_ sg13g2_a21oi_1
X_2411_ _1831_ _1826_ _1830_ VPWR VGND sg13g2_nand2_1
X_3391_ VPWR VGND _0916_ _0872_ _0915_ net711 _0917_ _0914_ sg13g2_a221oi_1
X_2342_ _1762_ _1505_ _1508_ VPWR VGND sg13g2_nand2_2
XFILLER_42_1010 VPWR VGND sg13g2_decap_8
X_2273_ VGND VPWR net750 _1691_ _1693_ _1692_ sg13g2_a21oi_1
X_4012_ _1420_ net814 u_ser.shadow_reg\[6\] VPWR VGND sg13g2_nand2b_1
XFILLER_38_723 VPWR VGND sg13g2_decap_8
XFILLER_37_244 VPWR VGND sg13g2_fill_2
XFILLER_25_428 VPWR VGND sg13g2_decap_8
XFILLER_34_962 VPWR VGND sg13g2_decap_8
XFILLER_21_634 VPWR VGND sg13g2_decap_8
XFILLER_33_483 VPWR VGND sg13g2_decap_8
X_3727_ net616 _1187_ _1203_ VPWR VGND sg13g2_nor2_1
X_3658_ _0100_ _1147_ _1151_ _0664_ _1456_ VPWR VGND sg13g2_a22oi_1
X_2609_ _0027_ _1985_ _0198_ VPWR VGND sg13g2_nand2_1
X_3589_ _0085_ _0935_ _1097_ net618 _1452_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_549 VPWR VGND sg13g2_decap_8
XFILLER_29_734 VPWR VGND sg13g2_decap_8
XFILLER_44_715 VPWR VGND sg13g2_decap_8
XFILLER_17_907 VPWR VGND sg13g2_decap_8
XFILLER_24_461 VPWR VGND sg13g2_decap_8
XFILLER_25_995 VPWR VGND sg13g2_decap_8
XFILLER_40_954 VPWR VGND sg13g2_decap_8
XFILLER_12_623 VPWR VGND sg13g2_decap_8
XFILLER_8_649 VPWR VGND sg13g2_decap_8
XFILLER_7_137 VPWR VGND sg13g2_fill_2
XFILLER_4_844 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_39_509 VPWR VGND sg13g2_decap_8
XFILLER_47_564 VPWR VGND sg13g2_decap_8
XFILLER_16_962 VPWR VGND sg13g2_decap_8
XFILLER_35_759 VPWR VGND sg13g2_decap_8
XFILLER_43_770 VPWR VGND sg13g2_decap_8
X_2960_ _0515_ _0510_ _0514_ VPWR VGND sg13g2_xnor2_1
X_2891_ _0446_ _0447_ _0448_ VPWR VGND sg13g2_and2_1
XFILLER_31_976 VPWR VGND sg13g2_decap_8
Xclkbuf_5_3__f_sap_3_inst.alu.clk_regs clknet_4_1_0_sap_3_inst.alu.clk_regs clknet_5_3__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3512_ net606 VPWR _1033_ VGND net669 _1032_ sg13g2_o21ai_1
X_3443_ _0967_ net596 net32 VPWR VGND sg13g2_nand2b_1
X_3374_ _0900_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] net675 VPWR
+ VGND sg13g2_nand2_1
X_2325_ _1566_ _1744_ _1745_ VPWR VGND sg13g2_and2_1
X_2256_ net786 net783 net781 _1676_ VPWR VGND sg13g2_nand3_1
XFILLER_38_520 VPWR VGND sg13g2_decap_8
X_2187_ _1589_ _1606_ _1607_ VPWR VGND sg13g2_and2_1
XFILLER_26_737 VPWR VGND sg13g2_decap_8
XFILLER_38_597 VPWR VGND sg13g2_decap_8
XFILLER_41_707 VPWR VGND sg13g2_decap_8
XFILLER_22_965 VPWR VGND sg13g2_decap_8
XFILLER_49_1016 VPWR VGND sg13g2_decap_8
XFILLER_49_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_836 VPWR VGND sg13g2_decap_8
XFILLER_48_339 VPWR VGND sg13g2_decap_8
XFILLER_29_531 VPWR VGND sg13g2_decap_8
XFILLER_17_704 VPWR VGND sg13g2_decap_8
XFILLER_44_512 VPWR VGND sg13g2_decap_8
XFILLER_1_1018 VPWR VGND sg13g2_decap_8
XFILLER_16_203 VPWR VGND sg13g2_fill_2
XFILLER_44_589 VPWR VGND sg13g2_decap_8
XFILLER_9_903 VPWR VGND sg13g2_decap_8
XFILLER_13_921 VPWR VGND sg13g2_decap_8
XFILLER_25_792 VPWR VGND sg13g2_decap_8
XFILLER_31_239 VPWR VGND sg13g2_fill_1
Xclkbuf_5_10__f_sap_3_inst.alu.clk_regs clknet_4_5_0_sap_3_inst.alu.clk_regs clknet_5_10__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_40_751 VPWR VGND sg13g2_decap_8
XFILLER_12_497 VPWR VGND sg13g2_decap_8
XFILLER_13_998 VPWR VGND sg13g2_decap_8
XFILLER_4_641 VPWR VGND sg13g2_decap_8
X_2110_ _1522_ _1529_ _1530_ VPWR VGND sg13g2_nor2b_2
X_3090_ VGND VPWR _1516_ _1746_ _0618_ _1842_ sg13g2_a21oi_1
Xhold2 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[5\] VPWR VGND net51 sg13g2_dlygate4sd3_1
X_2041_ VPWR _1463_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] VGND
+ sg13g2_inv_1
XFILLER_47_361 VPWR VGND sg13g2_decap_8
XFILLER_35_556 VPWR VGND sg13g2_decap_8
X_3992_ _1405_ sap_3_inst.alu.act\[4\] net583 VPWR VGND sg13g2_nand2_1
XFILLER_23_729 VPWR VGND sg13g2_decap_8
X_2943_ _0492_ _0494_ _0491_ _0499_ VPWR VGND _0498_ sg13g2_nand4_1
X_2874_ VGND VPWR net802 _1471_ _0432_ _0387_ sg13g2_a21oi_1
XFILLER_31_773 VPWR VGND sg13g2_decap_8
X_3426_ _0950_ net667 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] net681
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3357_ VGND VPWR _0884_ _0882_ _0881_ sg13g2_or2_1
X_2308_ VGND VPWR _1600_ _1609_ _1728_ _1648_ sg13g2_a21oi_1
X_3288_ _0816_ _1613_ _1697_ VPWR VGND sg13g2_nand2_1
X_2239_ net734 _1603_ _1659_ VPWR VGND sg13g2_nor2_1
XFILLER_39_873 VPWR VGND sg13g2_decap_8
XFILLER_26_534 VPWR VGND sg13g2_decap_8
XFILLER_41_504 VPWR VGND sg13g2_decap_8
XFILLER_16_1004 VPWR VGND sg13g2_decap_8
XFILLER_22_762 VPWR VGND sg13g2_decap_8
XFILLER_10_935 VPWR VGND sg13g2_decap_8
XFILLER_1_633 VPWR VGND sg13g2_decap_8
XFILLER_49_659 VPWR VGND sg13g2_decap_8
XFILLER_0_198 VPWR VGND sg13g2_fill_2
XFILLER_17_501 VPWR VGND sg13g2_decap_8
XFILLER_45_865 VPWR VGND sg13g2_decap_8
XFILLER_17_578 VPWR VGND sg13g2_decap_8
XFILLER_44_386 VPWR VGND sg13g2_decap_8
XFILLER_9_700 VPWR VGND sg13g2_decap_8
XFILLER_32_559 VPWR VGND sg13g2_decap_8
XFILLER_8_210 VPWR VGND sg13g2_fill_2
XFILLER_13_795 VPWR VGND sg13g2_decap_8
XFILLER_9_777 VPWR VGND sg13g2_decap_8
X_2590_ _2000_ net633 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] net641
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_994 VPWR VGND sg13g2_decap_8
XFILLER_5_54 VPWR VGND sg13g2_fill_1
X_3211_ _0739_ net660 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] net680
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4191_ net846 VGND VPWR _0155_ sap_3_inst.reg_file.array_serializer_inst.state\[1\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_1
X_3142_ net742 net726 _0670_ VPWR VGND sg13g2_and2_1
X_3073_ net739 net34 _0602_ VPWR VGND sg13g2_nor2_1
XFILLER_27_309 VPWR VGND sg13g2_fill_2
X_2024_ _1446_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[3\] VPWR VGND
+ sg13g2_inv_2
XFILLER_36_843 VPWR VGND sg13g2_decap_8
XFILLER_23_526 VPWR VGND sg13g2_decap_8
X_3975_ VGND VPWR _0323_ net709 _1392_ _1391_ sg13g2_a21oi_1
X_2926_ _0482_ net793 sap_3_inst.alu.tmp\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_31_570 VPWR VGND sg13g2_decap_8
X_2857_ _0415_ net798 net720 VPWR VGND sg13g2_xnor2_1
X_2788_ _0323_ net762 _0349_ VPWR VGND sg13g2_xor2_1
Xfanout723 _1730_ net723 VPWR VGND sg13g2_buf_8
Xfanout712 _0826_ net712 VPWR VGND sg13g2_buf_8
X_3409_ _0934_ _0933_ _0932_ VPWR VGND sg13g2_nand2b_1
Xfanout701 _0644_ net701 VPWR VGND sg13g2_buf_8
Xfanout745 _1509_ net745 VPWR VGND sg13g2_buf_8
Xfanout734 _1560_ net734 VPWR VGND sg13g2_buf_8
Xfanout756 _1521_ net756 VPWR VGND sg13g2_buf_8
Xfanout767 _1513_ net767 VPWR VGND sg13g2_buf_8
Xfanout778 net779 net778 VPWR VGND sg13g2_buf_2
Xfanout789 sap_3_inst.alu.acc\[7\] net789 VPWR VGND sg13g2_buf_8
XFILLER_46_618 VPWR VGND sg13g2_decap_8
Xclkbuf_4_10_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_10_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_39_670 VPWR VGND sg13g2_decap_8
XFILLER_27_854 VPWR VGND sg13g2_decap_8
XFILLER_38_191 VPWR VGND sg13g2_fill_2
XFILLER_42_835 VPWR VGND sg13g2_decap_8
XFILLER_14_548 VPWR VGND sg13g2_decap_8
XFILLER_14_41 VPWR VGND sg13g2_fill_1
XFILLER_10_732 VPWR VGND sg13g2_decap_8
XFILLER_6_747 VPWR VGND sg13g2_decap_8
XFILLER_2_931 VPWR VGND sg13g2_decap_8
XFILLER_7_1013 VPWR VGND sg13g2_decap_8
XFILLER_49_456 VPWR VGND sg13g2_decap_8
XFILLER_37_618 VPWR VGND sg13g2_decap_8
XFILLER_18_854 VPWR VGND sg13g2_decap_8
XFILLER_45_662 VPWR VGND sg13g2_decap_8
XFILLER_17_342 VPWR VGND sg13g2_fill_2
XFILLER_33_868 VPWR VGND sg13g2_decap_8
XFILLER_20_507 VPWR VGND sg13g2_decap_8
X_3760_ net611 _0892_ _1222_ _1223_ VPWR VGND sg13g2_nor3_1
XFILLER_13_592 VPWR VGND sg13g2_decap_8
X_2711_ _0287_ net576 _1970_ VPWR VGND sg13g2_nand2_2
XFILLER_9_574 VPWR VGND sg13g2_decap_8
X_3691_ _1177_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] net578 _0107_
+ VPWR VGND sg13g2_mux2_1
X_2642_ _0205_ VPWR _0026_ VGND _0228_ _0229_ sg13g2_o21ai_1
X_2573_ _1983_ VPWR _1984_ VGND net789 _1867_ sg13g2_o21ai_1
XFILLER_5_791 VPWR VGND sg13g2_decap_8
X_4174_ net844 VGND VPWR _0138_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\]
+ clknet_5_27__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3125_ _0650_ _0652_ _0648_ _0653_ VPWR VGND sg13g2_nand3_1
X_3056_ VGND VPWR net572 net716 _0053_ _0596_ sg13g2_a21oi_1
XFILLER_27_139 VPWR VGND sg13g2_decap_4
XFILLER_36_640 VPWR VGND sg13g2_decap_8
XFILLER_24_846 VPWR VGND sg13g2_decap_8
X_3958_ net609 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] _1382_ _0169_
+ VPWR VGND sg13g2_a21o_1
Xclkbuf_4_2_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_2_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2909_ _0466_ net625 _0463_ VPWR VGND sg13g2_nand2_1
X_3889_ _1318_ _1320_ _1315_ _1322_ VPWR VGND _1321_ sg13g2_nand4_1
Xfanout575 _0334_ net575 VPWR VGND sg13g2_buf_2
XFILLER_47_949 VPWR VGND sg13g2_decap_8
XFILLER_46_415 VPWR VGND sg13g2_decap_8
Xfanout597 _0849_ net597 VPWR VGND sg13g2_buf_8
Xfanout586 _0863_ net586 VPWR VGND sg13g2_buf_8
XFILLER_27_651 VPWR VGND sg13g2_decap_8
XFILLER_42_632 VPWR VGND sg13g2_decap_8
XFILLER_15_868 VPWR VGND sg13g2_decap_8
XFILLER_14_367 VPWR VGND sg13g2_fill_1
XFILLER_23_890 VPWR VGND sg13g2_decap_8
XFILLER_30_849 VPWR VGND sg13g2_decap_8
XFILLER_6_544 VPWR VGND sg13g2_decap_8
XFILLER_29_1014 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_4
XFILLER_38_905 VPWR VGND sg13g2_decap_8
XFILLER_18_651 VPWR VGND sg13g2_decap_8
XFILLER_46_982 VPWR VGND sg13g2_decap_8
XFILLER_33_665 VPWR VGND sg13g2_decap_8
XFILLER_36_1018 VPWR VGND sg13g2_decap_8
XFILLER_21_816 VPWR VGND sg13g2_decap_8
X_3812_ VGND VPWR _1080_ _1259_ _1260_ _1077_ sg13g2_a21oi_1
X_3743_ _1189_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] net594 _0126_
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_371 VPWR VGND sg13g2_fill_2
X_3674_ VPWR _1164_ _1163_ VGND sg13g2_inv_1
X_2625_ _0214_ _0213_ _1723_ VPWR VGND sg13g2_nand2b_1
X_2556_ _1968_ net633 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] net635
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2487_ VGND VPWR net629 _1902_ _1903_ _1901_ sg13g2_a21oi_1
X_4226_ net844 VGND VPWR _0189_ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_2
X_4157_ net828 VGND VPWR _0121_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\]
+ clknet_5_14__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_916 VPWR VGND sg13g2_decap_8
X_3108_ _0636_ net743 _1711_ VPWR VGND sg13g2_nand2_1
XFILLER_28_448 VPWR VGND sg13g2_decap_4
X_4088_ net834 VGND VPWR _0052_ sap_3_inst.alu.tmp\[2\] clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3039_ _0584_ net775 _0317_ VPWR VGND sg13g2_nand2_1
XFILLER_37_982 VPWR VGND sg13g2_decap_8
XFILLER_24_643 VPWR VGND sg13g2_decap_8
XFILLER_12_805 VPWR VGND sg13g2_decap_8
XFILLER_20_871 VPWR VGND sg13g2_decap_8
XFILLER_3_547 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_4_1005 VPWR VGND sg13g2_decap_8
XFILLER_47_746 VPWR VGND sg13g2_decap_8
XFILLER_46_278 VPWR VGND sg13g2_decap_4
XFILLER_36_61 VPWR VGND sg13g2_fill_2
XFILLER_43_952 VPWR VGND sg13g2_decap_8
XFILLER_14_142 VPWR VGND sg13g2_fill_2
XFILLER_15_665 VPWR VGND sg13g2_decap_8
XFILLER_30_646 VPWR VGND sg13g2_decap_8
XFILLER_11_860 VPWR VGND sg13g2_decap_8
XFILLER_7_831 VPWR VGND sg13g2_decap_8
X_2410_ net737 _1828_ _1829_ _1830_ VPWR VGND sg13g2_nor3_1
X_3390_ _0869_ VPWR _0916_ VGND net11 _0850_ sg13g2_o21ai_1
X_2341_ VGND VPWR _1761_ _1760_ _1539_ sg13g2_or2_1
X_2272_ net776 net751 _1648_ _1692_ VPWR VGND sg13g2_nor3_1
X_4011_ u_ser.shadow_reg\[7\] u_ser.bit_pos\[1\] _1419_ VPWR VGND net814 sg13g2_nand3b_1
XFILLER_38_702 VPWR VGND sg13g2_decap_8
XFILLER_25_407 VPWR VGND sg13g2_decap_8
XFILLER_26_919 VPWR VGND sg13g2_decap_8
XFILLER_38_779 VPWR VGND sg13g2_decap_8
XFILLER_34_941 VPWR VGND sg13g2_decap_8
XFILLER_21_613 VPWR VGND sg13g2_decap_8
X_3726_ _0117_ _0935_ _1202_ net616 _1449_ VPWR VGND sg13g2_a22oi_1
X_3657_ VGND VPWR _1148_ _1150_ _1151_ net624 sg13g2_a21oi_1
X_2608_ _0197_ VPWR _0198_ VGND _1868_ net19 sg13g2_o21ai_1
X_3588_ net618 _0938_ _1096_ _1097_ VPWR VGND sg13g2_nor3_1
X_2539_ _1951_ _1949_ VPWR VGND _1947_ sg13g2_nand2b_2
XFILLER_0_528 VPWR VGND sg13g2_decap_8
XFILLER_29_713 VPWR VGND sg13g2_decap_8
X_4209_ net845 VGND VPWR _0173_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\]
+ clknet_5_25__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_43_259 VPWR VGND sg13g2_fill_2
XFILLER_12_602 VPWR VGND sg13g2_decap_8
XFILLER_24_440 VPWR VGND sg13g2_decap_8
XFILLER_25_974 VPWR VGND sg13g2_decap_8
XFILLER_40_933 VPWR VGND sg13g2_decap_8
XFILLER_11_101 VPWR VGND sg13g2_fill_2
XFILLER_8_628 VPWR VGND sg13g2_decap_8
XFILLER_11_145 VPWR VGND sg13g2_fill_2
XFILLER_12_679 VPWR VGND sg13g2_decap_8
XFILLER_4_823 VPWR VGND sg13g2_decap_8
XFILLER_26_1017 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_543 VPWR VGND sg13g2_decap_8
XFILLER_47_71 VPWR VGND sg13g2_fill_1
XFILLER_35_738 VPWR VGND sg13g2_decap_8
XFILLER_16_941 VPWR VGND sg13g2_decap_8
X_2890_ VGND VPWR _0412_ _0413_ _0447_ _0414_ sg13g2_a21oi_1
XFILLER_31_955 VPWR VGND sg13g2_decap_8
XFILLER_8_10 VPWR VGND sg13g2_fill_1
X_3511_ _1032_ _0721_ _0805_ VPWR VGND sg13g2_xnor2_1
X_3442_ _0965_ VPWR _0966_ VGND net622 _0962_ sg13g2_o21ai_1
X_3373_ _0899_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[2\] net586 VPWR
+ VGND sg13g2_nand2_1
X_2324_ _1744_ net734 net733 VPWR VGND sg13g2_nand2_1
XFILLER_26_0 VPWR VGND sg13g2_fill_2
X_2255_ _1444_ _1584_ _1675_ VPWR VGND sg13g2_nor2_1
X_2186_ _1592_ net750 _1604_ _1606_ VPWR VGND sg13g2_nor3_1
XFILLER_26_716 VPWR VGND sg13g2_decap_8
XFILLER_38_576 VPWR VGND sg13g2_decap_8
XFILLER_22_944 VPWR VGND sg13g2_decap_8
XFILLER_21_487 VPWR VGND sg13g2_decap_8
XFILLER_5_609 VPWR VGND sg13g2_decap_8
X_3709_ _1192_ _1190_ _1191_ VPWR VGND sg13g2_nand2_1
XFILLER_1_815 VPWR VGND sg13g2_decap_8
XFILLER_48_318 VPWR VGND sg13g2_decap_8
XFILLER_29_510 VPWR VGND sg13g2_decap_8
XFILLER_29_587 VPWR VGND sg13g2_decap_8
XFILLER_44_568 VPWR VGND sg13g2_decap_8
XFILLER_13_900 VPWR VGND sg13g2_decap_8
XFILLER_25_771 VPWR VGND sg13g2_decap_8
XFILLER_40_730 VPWR VGND sg13g2_decap_8
XFILLER_13_977 VPWR VGND sg13g2_decap_8
XFILLER_8_436 VPWR VGND sg13g2_fill_1
XFILLER_9_959 VPWR VGND sg13g2_decap_8
XFILLER_32_1021 VPWR VGND sg13g2_decap_8
XFILLER_33_84 VPWR VGND sg13g2_fill_1
XFILLER_4_620 VPWR VGND sg13g2_decap_8
XFILLER_4_697 VPWR VGND sg13g2_decap_8
XFILLER_0_892 VPWR VGND sg13g2_decap_8
Xhold3 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[7\] VPWR VGND net52 sg13g2_dlygate4sd3_1
XFILLER_47_340 VPWR VGND sg13g2_decap_8
X_2040_ VPWR _1462_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] VGND
+ sg13g2_inv_1
XFILLER_48_885 VPWR VGND sg13g2_decap_8
X_4048__13 VPWR net49 clknet_leaf_1_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_35_535 VPWR VGND sg13g2_decap_8
X_3991_ VGND VPWR _0463_ net710 _1404_ _1403_ sg13g2_a21oi_1
XFILLER_23_708 VPWR VGND sg13g2_decap_8
X_2942_ VGND VPWR _0498_ _0497_ _0327_ sg13g2_or2_1
XFILLER_31_752 VPWR VGND sg13g2_decap_8
X_2873_ VPWR VGND net796 _0430_ net682 net801 _0431_ net683 sg13g2_a221oi_1
XFILLER_30_251 VPWR VGND sg13g2_fill_1
XFILLER_8_992 VPWR VGND sg13g2_decap_8
X_3425_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] _0948_
+ net657 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\] _0949_ net661 sg13g2_a221oi_1
X_3356_ _0881_ _0882_ _0883_ VPWR VGND sg13g2_nor2_2
X_2307_ _1598_ net749 _1589_ _1727_ VPWR VGND sg13g2_nand3_1
X_3287_ VGND VPWR _0815_ _0814_ _0667_ sg13g2_or2_1
X_2238_ net748 _1657_ _1658_ VPWR VGND sg13g2_nor2_1
XFILLER_39_852 VPWR VGND sg13g2_decap_8
XFILLER_26_513 VPWR VGND sg13g2_decap_8
X_2169_ _1589_ _1582_ _1587_ net753 VPWR VGND sg13g2_and3_1
XFILLER_22_741 VPWR VGND sg13g2_decap_8
XFILLER_10_914 VPWR VGND sg13g2_decap_8
XFILLER_6_929 VPWR VGND sg13g2_decap_8
XFILLER_5_406 VPWR VGND sg13g2_fill_1
XFILLER_1_612 VPWR VGND sg13g2_decap_8
XFILLER_49_638 VPWR VGND sg13g2_decap_8
XFILLER_1_689 VPWR VGND sg13g2_decap_8
XFILLER_23_1009 VPWR VGND sg13g2_decap_8
XFILLER_48_148 VPWR VGND sg13g2_fill_2
XFILLER_28_40 VPWR VGND sg13g2_fill_1
XFILLER_45_844 VPWR VGND sg13g2_decap_8
XFILLER_44_365 VPWR VGND sg13g2_decap_8
XFILLER_17_557 VPWR VGND sg13g2_decap_8
XFILLER_32_538 VPWR VGND sg13g2_decap_8
XFILLER_13_774 VPWR VGND sg13g2_decap_8
XFILLER_9_756 VPWR VGND sg13g2_decap_8
XFILLER_5_973 VPWR VGND sg13g2_decap_8
XFILLER_4_494 VPWR VGND sg13g2_decap_8
X_3210_ _0738_ net665 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] net679
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4190_ net846 VGND VPWR _0154_ sap_3_inst.reg_file.array_serializer_inst.state\[0\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_1
X_3141_ VGND VPWR _1623_ _0668_ _0669_ _0275_ sg13g2_a21oi_1
X_3072_ net33 net770 net738 _0064_ VPWR VGND sg13g2_mux2_1
XFILLER_36_822 VPWR VGND sg13g2_decap_8
XFILLER_48_682 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk_div_out clk_div_out clknet_0_clk_div_out VPWR VGND sg13g2_buf_8
X_2023_ _1445_ net800 VPWR VGND sg13g2_inv_2
XFILLER_35_332 VPWR VGND sg13g2_fill_1
XFILLER_23_505 VPWR VGND sg13g2_decap_8
XFILLER_39_1027 VPWR VGND sg13g2_fill_2
XFILLER_36_899 VPWR VGND sg13g2_decap_8
X_3974_ _1459_ net709 _1391_ VPWR VGND sg13g2_nor2_1
X_2925_ VGND VPWR _0477_ _0479_ _0481_ _0480_ sg13g2_a21oi_1
X_2856_ net798 net720 _0414_ VPWR VGND sg13g2_nor2_1
X_2787_ _0348_ net762 VPWR VGND _0323_ sg13g2_nand2b_2
XFILLER_49_28 VPWR VGND sg13g2_decap_8
XFILLER_49_39 VPWR VGND sg13g2_fill_2
Xfanout724 net725 net724 VPWR VGND sg13g2_buf_8
Xfanout713 _0826_ net713 VPWR VGND sg13g2_buf_8
X_3408_ _0908_ _0930_ net590 _0933_ VPWR VGND sg13g2_nand3_1
Xfanout702 _0644_ net702 VPWR VGND sg13g2_buf_2
Xfanout735 _1559_ net735 VPWR VGND sg13g2_buf_8
Xfanout746 _1631_ net746 VPWR VGND sg13g2_buf_8
Xfanout757 _1517_ net757 VPWR VGND sg13g2_buf_8
X_3339_ VGND VPWR _0669_ _0866_ _0867_ _0685_ sg13g2_a21oi_1
Xfanout768 sap_3_inst.controller.opcode\[7\] net768 VPWR VGND sg13g2_buf_8
Xfanout779 sap_3_inst.controller.opcode\[3\] net779 VPWR VGND sg13g2_buf_8
XFILLER_27_833 VPWR VGND sg13g2_decap_8
XFILLER_42_814 VPWR VGND sg13g2_decap_8
XFILLER_14_527 VPWR VGND sg13g2_decap_8
XFILLER_41_335 VPWR VGND sg13g2_decap_8
XFILLER_10_711 VPWR VGND sg13g2_decap_8
XFILLER_14_86 VPWR VGND sg13g2_fill_1
XFILLER_6_726 VPWR VGND sg13g2_decap_8
XFILLER_10_788 VPWR VGND sg13g2_decap_8
XFILLER_2_910 VPWR VGND sg13g2_decap_8
XFILLER_2_987 VPWR VGND sg13g2_decap_8
XFILLER_1_486 VPWR VGND sg13g2_decap_8
XFILLER_49_435 VPWR VGND sg13g2_decap_8
XFILLER_39_61 VPWR VGND sg13g2_fill_1
XFILLER_18_833 VPWR VGND sg13g2_decap_8
XFILLER_45_641 VPWR VGND sg13g2_decap_8
XFILLER_33_847 VPWR VGND sg13g2_decap_8
XFILLER_13_571 VPWR VGND sg13g2_decap_8
XFILLER_9_553 VPWR VGND sg13g2_decap_8
X_2710_ _1673_ _1994_ net11 VPWR VGND sg13g2_nor2_2
X_3690_ _1177_ _1176_ _1050_ VPWR VGND sg13g2_nand2b_1
X_2641_ _0227_ _1867_ _0204_ _0229_ VPWR VGND sg13g2_a21o_1
X_2572_ _1983_ _1867_ _1982_ VPWR VGND sg13g2_nand2_1
XFILLER_5_770 VPWR VGND sg13g2_decap_8
X_4173_ net829 VGND VPWR _0137_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\]
+ clknet_5_15__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3124_ _0652_ _0651_ net728 _1685_ _1621_ VPWR VGND sg13g2_a22oi_1
X_3055_ sap_3_inst.alu.tmp\[3\] net715 _0596_ VPWR VGND sg13g2_nor2_1
XFILLER_24_825 VPWR VGND sg13g2_decap_8
XFILLER_36_696 VPWR VGND sg13g2_decap_8
X_3957_ net608 _1046_ _1047_ _1382_ VPWR VGND sg13g2_nor3_1
X_2908_ _0463_ _0435_ _0465_ VPWR VGND sg13g2_xor2_1
XFILLER_13_1019 VPWR VGND sg13g2_decap_8
X_3888_ _1321_ _1306_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] _1301_
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2839_ _0355_ VPWR _0398_ VGND _0322_ _0357_ sg13g2_o21ai_1
XFILLER_3_729 VPWR VGND sg13g2_decap_8
XFILLER_47_928 VPWR VGND sg13g2_decap_8
XFILLER_19_619 VPWR VGND sg13g2_decap_8
Xfanout576 _1674_ net576 VPWR VGND sg13g2_buf_8
Xfanout598 _0834_ net598 VPWR VGND sg13g2_buf_8
Xfanout587 _0863_ net587 VPWR VGND sg13g2_buf_1
XFILLER_27_630 VPWR VGND sg13g2_decap_8
XFILLER_26_140 VPWR VGND sg13g2_fill_1
XFILLER_42_611 VPWR VGND sg13g2_decap_8
XFILLER_15_847 VPWR VGND sg13g2_decap_8
XFILLER_42_688 VPWR VGND sg13g2_decap_8
XFILLER_30_828 VPWR VGND sg13g2_decap_8
XFILLER_41_51 VPWR VGND sg13g2_fill_1
XFILLER_6_523 VPWR VGND sg13g2_decap_8
XFILLER_10_585 VPWR VGND sg13g2_decap_8
XFILLER_2_784 VPWR VGND sg13g2_decap_8
XFILLER_2_45 VPWR VGND sg13g2_decap_8
XFILLER_46_961 VPWR VGND sg13g2_decap_8
XFILLER_18_630 VPWR VGND sg13g2_decap_8
XFILLER_33_644 VPWR VGND sg13g2_decap_8
X_3811_ _1259_ net609 net592 VPWR VGND sg13g2_nand2_1
XFILLER_14_891 VPWR VGND sg13g2_decap_8
X_3742_ _1185_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] net593 _0125_
+ VPWR VGND sg13g2_mux2_1
X_3673_ net607 VPWR _1163_ VGND _1008_ _1162_ sg13g2_o21ai_1
X_2624_ _0213_ _0208_ _0212_ net649 _1461_ VPWR VGND sg13g2_a22oi_1
X_2555_ _1967_ net636 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] net641
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2486_ _1902_ sap_3_inst.alu.flags\[5\] _1839_ VPWR VGND sg13g2_nand2_1
X_4225_ net831 VGND VPWR net73 sap_3_outputReg_start_sync clknet_3_0__leaf_clk sg13g2_dfrbpq_1
X_4156_ net825 VGND VPWR _0120_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3107_ net743 _1711_ _0635_ VPWR VGND sg13g2_and2_1
X_4087_ net834 VGND VPWR _0051_ sap_3_inst.alu.tmp\[1\] clknet_5_28__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_37_961 VPWR VGND sg13g2_decap_8
X_3038_ _0326_ net625 _0583_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_1_sap_3_inst.alu.clk clknet_1_1__leaf_sap_3_inst.alu.clk clknet_leaf_1_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_24_622 VPWR VGND sg13g2_decap_8
XFILLER_36_493 VPWR VGND sg13g2_decap_8
XFILLER_24_699 VPWR VGND sg13g2_decap_8
XFILLER_20_850 VPWR VGND sg13g2_decap_8
XFILLER_3_526 VPWR VGND sg13g2_decap_8
XFILLER_47_725 VPWR VGND sg13g2_decap_8
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
XFILLER_28_994 VPWR VGND sg13g2_decap_8
XFILLER_43_931 VPWR VGND sg13g2_decap_8
XFILLER_15_644 VPWR VGND sg13g2_decap_8
XFILLER_42_485 VPWR VGND sg13g2_decap_8
XFILLER_30_625 VPWR VGND sg13g2_decap_8
XFILLER_7_810 VPWR VGND sg13g2_decap_8
XFILLER_7_887 VPWR VGND sg13g2_decap_8
X_2340_ net727 _1740_ _1760_ VPWR VGND sg13g2_nor2_1
X_2271_ _1645_ _1690_ net733 _1691_ VPWR VGND sg13g2_nand3_1
XFILLER_2_581 VPWR VGND sg13g2_decap_8
X_4010_ _1418_ VPWR _0186_ VGND u_ser.state\[1\] _1438_ sg13g2_o21ai_1
XFILLER_37_246 VPWR VGND sg13g2_fill_1
XFILLER_38_758 VPWR VGND sg13g2_decap_8
XFILLER_19_983 VPWR VGND sg13g2_decap_8
XFILLER_34_920 VPWR VGND sg13g2_decap_8
XFILLER_45_290 VPWR VGND sg13g2_fill_1
XFILLER_33_463 VPWR VGND sg13g2_fill_2
XFILLER_34_997 VPWR VGND sg13g2_decap_8
XFILLER_20_146 VPWR VGND sg13g2_decap_8
XFILLER_20_157 VPWR VGND sg13g2_fill_1
XFILLER_21_669 VPWR VGND sg13g2_decap_8
X_3725_ net616 _1054_ _1202_ VPWR VGND sg13g2_nor2_1
X_3656_ _1149_ VPWR _1150_ VGND _1673_ _1994_ sg13g2_o21ai_1
X_2607_ VGND VPWR _1868_ _0196_ _0197_ _1961_ sg13g2_a21oi_1
X_3587_ VPWR VGND _0287_ _0850_ _1075_ net572 _1096_ net684 sg13g2_a221oi_1
X_2538_ VGND VPWR _1950_ _1949_ _1947_ sg13g2_or2_1
XFILLER_0_507 VPWR VGND sg13g2_decap_8
X_2469_ _1887_ net640 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] net645
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] VPWR VGND sg13g2_a22oi_1
X_4208_ net821 VGND VPWR _0172_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\]
+ clknet_5_18__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4139_ net824 VGND VPWR _0103_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\]
+ clknet_5_11__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_257 VPWR VGND sg13g2_fill_2
XFILLER_29_769 VPWR VGND sg13g2_decap_8
XFILLER_43_238 VPWR VGND sg13g2_fill_1
XFILLER_25_953 VPWR VGND sg13g2_decap_8
XFILLER_40_912 VPWR VGND sg13g2_decap_8
XFILLER_19_1025 VPWR VGND sg13g2_decap_4
XFILLER_24_496 VPWR VGND sg13g2_decap_8
XFILLER_40_989 VPWR VGND sg13g2_decap_8
XFILLER_8_607 VPWR VGND sg13g2_decap_8
XFILLER_12_658 VPWR VGND sg13g2_decap_8
XFILLER_4_802 VPWR VGND sg13g2_decap_8
XFILLER_4_879 VPWR VGND sg13g2_decap_8
XFILLER_47_522 VPWR VGND sg13g2_decap_8
XFILLER_47_599 VPWR VGND sg13g2_decap_8
XFILLER_35_717 VPWR VGND sg13g2_decap_8
XFILLER_16_920 VPWR VGND sg13g2_decap_8
XFILLER_28_791 VPWR VGND sg13g2_decap_8
XFILLER_42_271 VPWR VGND sg13g2_fill_1
XFILLER_16_997 VPWR VGND sg13g2_decap_8
XFILLER_31_934 VPWR VGND sg13g2_decap_8
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_30_499 VPWR VGND sg13g2_decap_8
X_3510_ net621 _1028_ _1029_ _1031_ VPWR VGND sg13g2_nor3_1
XFILLER_7_684 VPWR VGND sg13g2_decap_8
X_3441_ VPWR _0965_ _0964_ VGND sg13g2_inv_1
X_3372_ net586 sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[1\] _0895_ _0067_
+ VPWR VGND sg13g2_a21o_1
XFILLER_3_890 VPWR VGND sg13g2_decap_8
X_2323_ _1742_ VPWR _1743_ VGND _1554_ _1740_ sg13g2_o21ai_1
X_2254_ VPWR _1674_ _1673_ VGND sg13g2_inv_1
X_2185_ _1605_ _1590_ VPWR VGND _1580_ sg13g2_nand2b_2
XFILLER_38_555 VPWR VGND sg13g2_decap_8
XFILLER_19_780 VPWR VGND sg13g2_decap_8
XFILLER_22_923 VPWR VGND sg13g2_decap_8
XFILLER_34_794 VPWR VGND sg13g2_decap_8
X_3708_ _1191_ net597 net22 VPWR VGND sg13g2_nand2b_1
X_3639_ _1135_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] net624 VPWR
+ VGND sg13g2_nand2_1
XFILLER_29_566 VPWR VGND sg13g2_decap_8
XFILLER_44_547 VPWR VGND sg13g2_decap_8
XFILLER_16_238 VPWR VGND sg13g2_fill_2
XFILLER_17_739 VPWR VGND sg13g2_decap_8
XFILLER_25_750 VPWR VGND sg13g2_decap_8
XFILLER_13_956 VPWR VGND sg13g2_decap_8
XFILLER_40_786 VPWR VGND sg13g2_decap_8
XFILLER_9_938 VPWR VGND sg13g2_decap_8
XFILLER_12_466 VPWR VGND sg13g2_fill_1
XFILLER_32_1000 VPWR VGND sg13g2_decap_8
XFILLER_4_676 VPWR VGND sg13g2_decap_8
XFILLER_3_164 VPWR VGND sg13g2_fill_2
Xclkbuf_5_8__f_sap_3_inst.alu.clk_regs clknet_4_4_0_sap_3_inst.alu.clk_regs clknet_5_8__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_0_871 VPWR VGND sg13g2_decap_8
Xhold4 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[6\] VPWR VGND net53 sg13g2_dlygate4sd3_1
XFILLER_48_864 VPWR VGND sg13g2_decap_8
XFILLER_35_514 VPWR VGND sg13g2_decap_8
XFILLER_47_396 VPWR VGND sg13g2_decap_8
X_3990_ _1460_ _1389_ _1403_ VPWR VGND sg13g2_nor2_1
X_2941_ VGND VPWR _0497_ _0485_ _0464_ sg13g2_or2_1
XFILLER_16_794 VPWR VGND sg13g2_decap_8
XFILLER_31_731 VPWR VGND sg13g2_decap_8
X_2872_ _1951_ _0331_ _0421_ _0430_ VPWR VGND sg13g2_nor3_1
XFILLER_8_971 VPWR VGND sg13g2_decap_8
X_3424_ net676 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] net671 _0948_
+ VPWR VGND sg13g2_a21o_1
X_3355_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[1\] net621 _0882_ VPWR
+ VGND sg13g2_nor2_1
X_2306_ _1726_ _1640_ _1724_ VPWR VGND sg13g2_nand2_1
X_3286_ _0681_ VPWR _0814_ VGND net751 _1687_ sg13g2_o21ai_1
X_2237_ _1657_ _1507_ net746 VPWR VGND sg13g2_nand2_2
XFILLER_39_831 VPWR VGND sg13g2_decap_8
X_2168_ _1528_ _1568_ _1523_ _1588_ VPWR VGND sg13g2_nand3_1
XFILLER_14_709 VPWR VGND sg13g2_decap_8
X_2099_ _1519_ net774 net772 VPWR VGND sg13g2_nand2_1
XFILLER_26_569 VPWR VGND sg13g2_decap_8
XFILLER_41_539 VPWR VGND sg13g2_decap_8
XFILLER_22_720 VPWR VGND sg13g2_decap_8
XFILLER_34_591 VPWR VGND sg13g2_decap_8
XFILLER_6_908 VPWR VGND sg13g2_decap_8
XFILLER_22_797 VPWR VGND sg13g2_decap_8
Xclkbuf_5_15__f_sap_3_inst.alu.clk_regs clknet_4_7_0_sap_3_inst.alu.clk_regs clknet_5_15__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_1_668 VPWR VGND sg13g2_decap_8
XFILLER_49_617 VPWR VGND sg13g2_decap_8
XFILLER_28_30 VPWR VGND sg13g2_fill_1
XFILLER_29_352 VPWR VGND sg13g2_fill_2
XFILLER_45_823 VPWR VGND sg13g2_decap_8
XFILLER_17_536 VPWR VGND sg13g2_decap_8
XFILLER_28_96 VPWR VGND sg13g2_fill_1
XFILLER_32_517 VPWR VGND sg13g2_decap_8
XFILLER_13_753 VPWR VGND sg13g2_decap_8
XFILLER_8_212 VPWR VGND sg13g2_fill_1
XFILLER_9_735 VPWR VGND sg13g2_decap_8
XFILLER_40_583 VPWR VGND sg13g2_decap_8
XFILLER_5_952 VPWR VGND sg13g2_decap_8
X_3140_ _0622_ _0667_ _0668_ VPWR VGND sg13g2_nor2_1
XFILLER_48_661 VPWR VGND sg13g2_decap_8
X_3071_ net22 net772 net738 _0063_ VPWR VGND sg13g2_mux2_1
XFILLER_36_801 VPWR VGND sg13g2_decap_8
X_2022_ net780 _1444_ VPWR VGND sg13g2_inv_4
XFILLER_36_878 VPWR VGND sg13g2_decap_8
XFILLER_39_1006 VPWR VGND sg13g2_decap_8
XFILLER_35_366 VPWR VGND sg13g2_fill_1
X_3973_ _0316_ net709 _1390_ VPWR VGND sg13g2_nor2b_2
XFILLER_16_591 VPWR VGND sg13g2_decap_8
X_2924_ net714 VPWR _0480_ VGND _0477_ _0479_ sg13g2_o21ai_1
X_2855_ _0413_ net798 net720 VPWR VGND sg13g2_nand2_1
X_2786_ _0347_ net762 _0323_ VPWR VGND sg13g2_nand2_1
Xfanout714 _1944_ net714 VPWR VGND sg13g2_buf_8
X_3407_ VGND VPWR net590 _0908_ _0932_ _0930_ sg13g2_a21oi_1
Xfanout703 net706 net703 VPWR VGND sg13g2_buf_8
Xfanout736 _1552_ net736 VPWR VGND sg13g2_buf_8
X_3338_ _0675_ _0865_ _1624_ _0866_ VPWR VGND sg13g2_nand3_1
Xfanout758 _1503_ net758 VPWR VGND sg13g2_buf_8
Xfanout747 _1631_ net747 VPWR VGND sg13g2_buf_1
Xfanout725 _1714_ net725 VPWR VGND sg13g2_buf_8
Xfanout769 sap_3_inst.controller.opcode\[7\] net769 VPWR VGND sg13g2_buf_1
XFILLER_22_1021 VPWR VGND sg13g2_decap_8
XFILLER_27_812 VPWR VGND sg13g2_decap_8
X_3269_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] _0790_
+ net655 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] _0797_ net679 sg13g2_a221oi_1
XFILLER_14_506 VPWR VGND sg13g2_decap_8
XFILLER_27_889 VPWR VGND sg13g2_decap_8
XFILLER_22_594 VPWR VGND sg13g2_decap_8
XFILLER_6_705 VPWR VGND sg13g2_decap_8
XFILLER_10_767 VPWR VGND sg13g2_decap_8
XFILLER_2_966 VPWR VGND sg13g2_decap_8
XFILLER_49_414 VPWR VGND sg13g2_decap_8
XFILLER_18_812 VPWR VGND sg13g2_decap_8
XFILLER_45_620 VPWR VGND sg13g2_decap_8
XFILLER_44_141 VPWR VGND sg13g2_fill_2
XFILLER_45_697 VPWR VGND sg13g2_decap_8
XFILLER_18_889 VPWR VGND sg13g2_decap_8
XFILLER_32_314 VPWR VGND sg13g2_fill_2
XFILLER_33_826 VPWR VGND sg13g2_decap_8
XFILLER_13_550 VPWR VGND sg13g2_decap_8
XFILLER_9_532 VPWR VGND sg13g2_decap_8
X_2640_ sap_3_inst.alu.carry _1867_ _0228_ VPWR VGND sg13g2_nor2_1
X_2571_ net20 net572 VPWR VGND sg13g2_inv_2
X_4172_ net825 VGND VPWR _0136_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3123_ _1588_ VPWR _0651_ VGND net765 _1570_ sg13g2_o21ai_1
XFILLER_28_609 VPWR VGND sg13g2_decap_8
XFILLER_49_981 VPWR VGND sg13g2_decap_8
X_3054_ _0595_ VPWR _0052_ VGND _1471_ net715 sg13g2_o21ai_1
XFILLER_24_804 VPWR VGND sg13g2_decap_8
XFILLER_36_675 VPWR VGND sg13g2_decap_8
X_3956_ net812 net52 _1381_ _0168_ VPWR VGND sg13g2_a21o_1
X_2907_ _0464_ _0435_ _0451_ VPWR VGND sg13g2_nand2_1
XFILLER_32_881 VPWR VGND sg13g2_decap_8
X_3887_ _1320_ _1309_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] net810
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2838_ VGND VPWR _0393_ _0394_ _0397_ _0396_ sg13g2_a21oi_1
XFILLER_3_708 VPWR VGND sg13g2_decap_8
X_2769_ _0330_ _0327_ _0328_ VPWR VGND sg13g2_nand2_1
XFILLER_47_907 VPWR VGND sg13g2_decap_8
Xfanout577 _1674_ net577 VPWR VGND sg13g2_buf_1
Xfanout588 _0799_ net588 VPWR VGND sg13g2_buf_8
Xfanout599 _0834_ net599 VPWR VGND sg13g2_buf_8
XFILLER_15_826 VPWR VGND sg13g2_decap_8
XFILLER_27_686 VPWR VGND sg13g2_decap_8
XFILLER_42_667 VPWR VGND sg13g2_decap_8
XFILLER_30_807 VPWR VGND sg13g2_decap_8
XFILLER_6_502 VPWR VGND sg13g2_decap_8
XFILLER_10_564 VPWR VGND sg13g2_decap_8
XFILLER_6_579 VPWR VGND sg13g2_decap_8
XFILLER_2_763 VPWR VGND sg13g2_decap_8
XFILLER_49_222 VPWR VGND sg13g2_decap_8
XFILLER_49_288 VPWR VGND sg13g2_decap_8
XFILLER_37_417 VPWR VGND sg13g2_fill_1
XFILLER_46_940 VPWR VGND sg13g2_decap_8
XFILLER_18_686 VPWR VGND sg13g2_decap_8
XFILLER_45_494 VPWR VGND sg13g2_decap_8
XFILLER_33_623 VPWR VGND sg13g2_decap_8
X_3810_ VGND VPWR _1495_ net614 _0145_ _1258_ sg13g2_a21oi_1
XFILLER_14_870 VPWR VGND sg13g2_decap_8
X_3741_ _1210_ VPWR _0124_ VGND _1129_ net594 sg13g2_o21ai_1
X_3672_ net679 _1009_ _1162_ VPWR VGND sg13g2_nor2_1
X_2623_ net648 _0209_ _0210_ _0211_ _0212_ VPWR VGND sg13g2_and4_1
X_2554_ _1963_ _1965_ _1966_ VPWR VGND sg13g2_and2_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
X_2485_ net795 net628 _1901_ VPWR VGND sg13g2_nor2_1
X_4224_ net831 VGND VPWR _0187_ sap_3_outputReg_serial clknet_3_0__leaf_clk sg13g2_dfrbpq_1
X_4155_ net824 VGND VPWR _0119_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\]
+ clknet_5_10__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3106_ _0631_ _0632_ _0630_ _0634_ VPWR VGND _0633_ sg13g2_nand4_1
X_4086_ net834 VGND VPWR _0050_ sap_3_inst.alu.tmp\[0\] clknet_5_28__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_37_940 VPWR VGND sg13g2_decap_8
X_3037_ _0581_ VPWR _0582_ VGND _0551_ _0580_ sg13g2_o21ai_1
XFILLER_24_601 VPWR VGND sg13g2_decap_8
XFILLER_23_111 VPWR VGND sg13g2_fill_2
XFILLER_24_678 VPWR VGND sg13g2_decap_8
X_3939_ _1366_ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] _1306_
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_3_505 VPWR VGND sg13g2_decap_8
XFILLER_47_704 VPWR VGND sg13g2_decap_8
XFILLER_43_910 VPWR VGND sg13g2_decap_8
XFILLER_28_973 VPWR VGND sg13g2_decap_8
XFILLER_36_63 VPWR VGND sg13g2_fill_1
XFILLER_14_100 VPWR VGND sg13g2_fill_2
XFILLER_15_623 VPWR VGND sg13g2_decap_8
XFILLER_27_483 VPWR VGND sg13g2_decap_8
XFILLER_43_987 VPWR VGND sg13g2_decap_8
XFILLER_42_464 VPWR VGND sg13g2_decap_8
XFILLER_14_144 VPWR VGND sg13g2_fill_1
XFILLER_30_604 VPWR VGND sg13g2_decap_8
XFILLER_10_361 VPWR VGND sg13g2_fill_1
XFILLER_11_895 VPWR VGND sg13g2_decap_8
XFILLER_7_866 VPWR VGND sg13g2_decap_8
XFILLER_2_560 VPWR VGND sg13g2_decap_8
X_2270_ _1690_ _1504_ _1642_ VPWR VGND sg13g2_nand2_1
XFILLER_42_1024 VPWR VGND sg13g2_decap_4
XFILLER_38_737 VPWR VGND sg13g2_decap_8
XFILLER_19_962 VPWR VGND sg13g2_decap_8
XFILLER_34_976 VPWR VGND sg13g2_decap_8
XFILLER_33_497 VPWR VGND sg13g2_decap_8
XFILLER_21_648 VPWR VGND sg13g2_decap_8
X_3724_ VGND VPWR _1455_ net616 _0116_ _1201_ sg13g2_a21oi_1
X_3655_ _1149_ _0849_ _1138_ VPWR VGND sg13g2_nand2_2
X_2606_ _0196_ _2011_ _2014_ VPWR VGND sg13g2_xnor2_1
X_3586_ net618 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] _1095_ _0084_
+ VPWR VGND sg13g2_a21o_1
X_2537_ _1948_ net773 _1949_ VPWR VGND sg13g2_nor2b_2
X_2468_ _1886_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] net632
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] VPWR VGND sg13g2_a22oi_1
X_4207_ net841 VGND VPWR _0171_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\]
+ clknet_5_31__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2399_ _1819_ _1815_ _1818_ net650 _1494_ VPWR VGND sg13g2_a22oi_1
XFILLER_29_748 VPWR VGND sg13g2_decap_8
X_4138_ net842 VGND VPWR _0102_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\]
+ clknet_5_30__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_44_729 VPWR VGND sg13g2_decap_8
X_4069_ net832 VGND VPWR _0033_ sap_3_inst.alu.acc\[0\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_25_932 VPWR VGND sg13g2_decap_8
XFILLER_19_1004 VPWR VGND sg13g2_decap_8
XFILLER_11_103 VPWR VGND sg13g2_fill_1
XFILLER_12_637 VPWR VGND sg13g2_decap_8
XFILLER_24_475 VPWR VGND sg13g2_decap_8
XFILLER_40_968 VPWR VGND sg13g2_decap_8
XFILLER_4_858 VPWR VGND sg13g2_decap_8
XFILLER_47_501 VPWR VGND sg13g2_decap_8
XFILLER_47_578 VPWR VGND sg13g2_decap_8
XFILLER_28_770 VPWR VGND sg13g2_decap_8
XFILLER_16_976 VPWR VGND sg13g2_decap_8
XFILLER_27_291 VPWR VGND sg13g2_fill_1
XFILLER_43_784 VPWR VGND sg13g2_decap_8
XFILLER_31_913 VPWR VGND sg13g2_decap_8
XFILLER_15_497 VPWR VGND sg13g2_decap_8
XFILLER_30_478 VPWR VGND sg13g2_decap_8
XFILLER_11_692 VPWR VGND sg13g2_decap_8
XFILLER_7_663 VPWR VGND sg13g2_decap_8
X_3440_ net607 VPWR _0964_ VGND net671 _0963_ sg13g2_o21ai_1
X_3371_ _0898_ net590 net588 VPWR VGND sg13g2_xnor2_1
X_2322_ _1742_ net743 _1604_ VPWR VGND sg13g2_nand2_1
X_2253_ _1673_ _1538_ _1672_ _1505_ net758 VPWR VGND sg13g2_a22oi_1
X_2184_ _1580_ _1591_ _1604_ VPWR VGND sg13g2_nor2_2
XFILLER_38_534 VPWR VGND sg13g2_decap_8
XFILLER_22_902 VPWR VGND sg13g2_decap_8
XFILLER_34_773 VPWR VGND sg13g2_decap_8
XFILLER_22_979 VPWR VGND sg13g2_decap_8
X_3707_ _1190_ net602 _0981_ VPWR VGND sg13g2_nand2_1
X_3638_ _0097_ _1134_ _1069_ _1121_ _1499_ VPWR VGND sg13g2_a22oi_1
X_3569_ _1080_ VPWR _1081_ VGND _0695_ net590 sg13g2_o21ai_1
XFILLER_29_545 VPWR VGND sg13g2_decap_8
XFILLER_17_718 VPWR VGND sg13g2_decap_8
XFILLER_44_526 VPWR VGND sg13g2_decap_8
XFILLER_13_935 VPWR VGND sg13g2_decap_8
XFILLER_9_917 VPWR VGND sg13g2_decap_8
XFILLER_40_765 VPWR VGND sg13g2_decap_8
XFILLER_33_75 VPWR VGND sg13g2_fill_2
XFILLER_4_655 VPWR VGND sg13g2_decap_8
XFILLER_0_850 VPWR VGND sg13g2_decap_8
XFILLER_48_843 VPWR VGND sg13g2_decap_8
Xhold5 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[0\] VPWR VGND net54 sg13g2_dlygate4sd3_1
XFILLER_47_375 VPWR VGND sg13g2_decap_8
X_2940_ _0495_ _0485_ _0496_ VPWR VGND sg13g2_xor2_1
XFILLER_16_773 VPWR VGND sg13g2_decap_8
XFILLER_31_710 VPWR VGND sg13g2_decap_8
XFILLER_43_581 VPWR VGND sg13g2_decap_8
X_2871_ VPWR VGND _0329_ _0420_ _0428_ _0335_ _0429_ _0422_ sg13g2_a221oi_1
XFILLER_31_787 VPWR VGND sg13g2_decap_8
XFILLER_8_950 VPWR VGND sg13g2_decap_8
X_3423_ _0947_ net675 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] net678
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3354_ _0877_ _0880_ _0881_ VPWR VGND sg13g2_nor2_1
XFILLER_31_0 VPWR VGND sg13g2_fill_1
X_2305_ VPWR _1725_ _1724_ VGND sg13g2_inv_1
X_3285_ net751 _1687_ _0813_ VPWR VGND sg13g2_nor2_1
XFILLER_39_810 VPWR VGND sg13g2_decap_8
X_2236_ _1507_ net746 _1656_ VPWR VGND sg13g2_and2_1
XFILLER_39_887 VPWR VGND sg13g2_decap_8
X_2167_ _1528_ _1562_ _1526_ _1587_ VPWR VGND _1583_ sg13g2_nand4_1
XFILLER_38_397 VPWR VGND sg13g2_fill_2
X_2098_ net774 net772 _1518_ VPWR VGND sg13g2_and2_1
XFILLER_26_548 VPWR VGND sg13g2_decap_8
XFILLER_41_518 VPWR VGND sg13g2_decap_8
XFILLER_34_570 VPWR VGND sg13g2_decap_8
XFILLER_16_1018 VPWR VGND sg13g2_decap_8
XFILLER_22_776 VPWR VGND sg13g2_decap_8
XFILLER_10_949 VPWR VGND sg13g2_decap_8
Xclkbuf_regs_0_clk_div_two sap_3_inst.alu.clk sap_3_inst.alu.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_1_647 VPWR VGND sg13g2_decap_8
XFILLER_45_802 VPWR VGND sg13g2_decap_8
XFILLER_17_515 VPWR VGND sg13g2_decap_8
XFILLER_29_386 VPWR VGND sg13g2_fill_2
XFILLER_45_879 VPWR VGND sg13g2_decap_8
XFILLER_13_732 VPWR VGND sg13g2_decap_8
XFILLER_40_562 VPWR VGND sg13g2_decap_8
XFILLER_9_714 VPWR VGND sg13g2_decap_8
XFILLER_8_257 VPWR VGND sg13g2_fill_2
XFILLER_5_931 VPWR VGND sg13g2_decap_8
X_3070_ VGND VPWR _1442_ net738 _0062_ _0601_ sg13g2_a21oi_1
XFILLER_48_640 VPWR VGND sg13g2_decap_8
X_2021_ _1443_ net768 VPWR VGND sg13g2_inv_2
XFILLER_36_857 VPWR VGND sg13g2_decap_8
XFILLER_16_570 VPWR VGND sg13g2_decap_8
XFILLER_44_890 VPWR VGND sg13g2_decap_8
X_3972_ _1856_ _1388_ _1389_ VPWR VGND sg13g2_nor2_2
X_2923_ _0479_ net793 net720 VPWR VGND sg13g2_xnor2_1
X_2854_ VGND VPWR net801 net721 _0412_ _0395_ sg13g2_a21oi_1
XFILLER_31_584 VPWR VGND sg13g2_decap_8
X_2785_ _0339_ _0341_ _0343_ _0345_ _0346_ VPWR VGND sg13g2_and4_1
Xfanout715 _0593_ net715 VPWR VGND sg13g2_buf_8
X_3406_ _0931_ _0930_ VPWR VGND sg13g2_inv_2
Xfanout704 net705 net704 VPWR VGND sg13g2_buf_8
Xfanout737 _1552_ net737 VPWR VGND sg13g2_buf_1
Xfanout748 _1605_ net748 VPWR VGND sg13g2_buf_8
Xfanout726 _1702_ net726 VPWR VGND sg13g2_buf_8
X_3337_ _0266_ _0678_ _0813_ _0864_ _0865_ VPWR VGND sg13g2_nor4_1
Xfanout759 sap_3_inst.controller.stage\[2\] net759 VPWR VGND sg13g2_buf_8
XFILLER_22_1000 VPWR VGND sg13g2_decap_8
X_3268_ _0796_ net665 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] net668
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] VPWR VGND sg13g2_a22oi_1
X_3199_ _0725_ VPWR _0727_ VGND _1488_ net617 sg13g2_o21ai_1
X_2219_ _1639_ net758 net747 VPWR VGND sg13g2_nand2_2
XFILLER_39_684 VPWR VGND sg13g2_decap_8
XFILLER_27_868 VPWR VGND sg13g2_decap_8
XFILLER_42_849 VPWR VGND sg13g2_decap_8
XFILLER_14_55 VPWR VGND sg13g2_fill_1
XFILLER_22_573 VPWR VGND sg13g2_decap_8
XFILLER_10_746 VPWR VGND sg13g2_decap_8
XFILLER_2_945 VPWR VGND sg13g2_decap_8
XFILLER_7_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_334 VPWR VGND sg13g2_fill_1
XFILLER_18_868 VPWR VGND sg13g2_decap_8
XFILLER_45_676 VPWR VGND sg13g2_decap_8
XFILLER_32_304 VPWR VGND sg13g2_fill_1
XFILLER_33_805 VPWR VGND sg13g2_decap_8
XFILLER_41_882 VPWR VGND sg13g2_decap_8
XFILLER_9_511 VPWR VGND sg13g2_decap_8
XFILLER_9_588 VPWR VGND sg13g2_decap_8
X_2570_ _1971_ _1981_ _1982_ VPWR VGND sg13g2_and2_1
X_4240_ regFile_serial_start net30 VPWR VGND sg13g2_buf_8
X_4171_ net824 VGND VPWR _0135_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\]
+ clknet_5_9__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3122_ VPWR VGND net777 _0649_ _1823_ _1571_ _0650_ _1604_ sg13g2_a221oi_1
XFILLER_49_960 VPWR VGND sg13g2_decap_8
X_3053_ _0595_ net19 net715 VPWR VGND sg13g2_nand2_1
XFILLER_36_654 VPWR VGND sg13g2_decap_8
XFILLER_35_142 VPWR VGND sg13g2_fill_1
XFILLER_32_860 VPWR VGND sg13g2_decap_8
X_3955_ VPWR VGND _1380_ net812 _1375_ _1494_ _1381_ net808 sg13g2_a221oi_1
X_2906_ _0463_ _0451_ _0461_ VPWR VGND sg13g2_xnor2_1
X_3886_ _1319_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] _1307_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2837_ _0396_ net714 _0395_ VPWR VGND sg13g2_nand2b_1
X_2768_ _0329_ _0328_ VPWR VGND sg13g2_inv_2
XFILLER_2_208 VPWR VGND sg13g2_fill_1
X_2699_ _0280_ _0281_ _0282_ VPWR VGND sg13g2_nor2_1
Xfanout589 _0799_ net589 VPWR VGND sg13g2_buf_1
Xfanout578 _1174_ net578 VPWR VGND sg13g2_buf_8
XFILLER_46_429 VPWR VGND sg13g2_decap_8
XFILLER_39_481 VPWR VGND sg13g2_decap_8
XFILLER_15_805 VPWR VGND sg13g2_decap_8
XFILLER_27_665 VPWR VGND sg13g2_decap_8
XFILLER_42_646 VPWR VGND sg13g2_decap_8
XFILLER_41_112 VPWR VGND sg13g2_fill_1
XFILLER_10_543 VPWR VGND sg13g2_decap_8
XFILLER_6_558 VPWR VGND sg13g2_decap_8
XFILLER_2_742 VPWR VGND sg13g2_decap_8
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_201 VPWR VGND sg13g2_fill_1
XFILLER_38_919 VPWR VGND sg13g2_decap_8
XFILLER_49_267 VPWR VGND sg13g2_decap_8
XFILLER_46_996 VPWR VGND sg13g2_decap_8
XFILLER_45_473 VPWR VGND sg13g2_decap_8
XFILLER_18_665 VPWR VGND sg13g2_decap_8
XFILLER_33_602 VPWR VGND sg13g2_decap_8
XFILLER_32_145 VPWR VGND sg13g2_fill_2
XFILLER_33_679 VPWR VGND sg13g2_decap_8
X_3740_ _1210_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] net593 VPWR
+ VGND sg13g2_nand2_1
X_3671_ _1161_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] net623 VPWR
+ VGND sg13g2_nand2_1
X_2622_ _0211_ net633 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] net723
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2553_ _1965_ net642 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] net723
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2484_ _1723_ _1890_ _1898_ _1900_ VPWR VGND sg13g2_nor3_1
X_4223_ net831 VGND VPWR _0186_ u_ser.state\[1\] clknet_3_0__leaf_clk sg13g2_dfrbpq_2
X_4154_ net829 VGND VPWR _0118_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\]
+ clknet_5_25__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3105_ net725 _1769_ _1828_ _0625_ _0633_ VPWR VGND sg13g2_nor4_1
X_4085_ net838 VGND VPWR _0049_ sap_3_inst.alu.carry clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3036_ _0581_ net787 sap_3_inst.alu.tmp\[7\] VPWR VGND sg13g2_nand2b_1
XFILLER_37_996 VPWR VGND sg13g2_decap_8
XFILLER_12_819 VPWR VGND sg13g2_decap_8
XFILLER_24_657 VPWR VGND sg13g2_decap_8
X_3938_ net811 net51 _1365_ _0166_ VPWR VGND sg13g2_a21o_1
XFILLER_20_885 VPWR VGND sg13g2_decap_8
X_3869_ _1302_ sap_3_inst.reg_file.array_serializer_inst.word_index\[1\] sap_3_inst.reg_file.array_serializer_inst.word_index\[0\]
+ VPWR VGND sg13g2_nand2_2
XFILLER_4_1019 VPWR VGND sg13g2_decap_8
XFILLER_28_952 VPWR VGND sg13g2_decap_8
XFILLER_15_602 VPWR VGND sg13g2_decap_8
XFILLER_27_462 VPWR VGND sg13g2_decap_8
XFILLER_43_966 VPWR VGND sg13g2_decap_8
XFILLER_42_443 VPWR VGND sg13g2_decap_8
XFILLER_15_679 VPWR VGND sg13g2_decap_8
XFILLER_11_874 VPWR VGND sg13g2_decap_8
XFILLER_7_845 VPWR VGND sg13g2_decap_8
XFILLER_42_1003 VPWR VGND sg13g2_decap_8
XFILLER_38_716 VPWR VGND sg13g2_decap_8
XFILLER_19_941 VPWR VGND sg13g2_decap_8
XFILLER_46_793 VPWR VGND sg13g2_decap_8
XFILLER_34_955 VPWR VGND sg13g2_decap_8
XFILLER_21_627 VPWR VGND sg13g2_decap_8
XFILLER_33_465 VPWR VGND sg13g2_fill_1
X_3723_ net617 _1052_ _1146_ _1201_ VPWR VGND sg13g2_nor3_1
XFILLER_9_182 VPWR VGND sg13g2_fill_2
X_3654_ _1148_ _2008_ net685 VPWR VGND sg13g2_nand2_1
X_2605_ _2014_ _2012_ _2013_ VPWR VGND sg13g2_xnor2_1
X_3585_ VPWR VGND _1094_ net618 _1092_ net600 _1095_ _0909_ sg13g2_a221oi_1
X_2536_ _1948_ _1935_ _1551_ _1559_ _1545_ VPWR VGND sg13g2_a22oi_1
X_2467_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] net643
+ net647 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] _1885_ net722 sg13g2_a221oi_1
X_4206_ net820 VGND VPWR _0170_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\]
+ clknet_5_1__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2398_ net648 _1813_ _1816_ _1817_ _1818_ VPWR VGND sg13g2_and4_1
XFILLER_29_727 VPWR VGND sg13g2_decap_8
X_4137_ net819 VGND VPWR _0101_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\]
+ clknet_5_5__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_248 VPWR VGND sg13g2_fill_1
XFILLER_44_708 VPWR VGND sg13g2_decap_8
X_4068_ net834 VGND VPWR _0032_ sap_3_inst.alu.flags\[7\] net49 sg13g2_dfrbpq_1
XFILLER_25_911 VPWR VGND sg13g2_decap_8
X_3019_ _0571_ sap_3_inst.out\[1\] net717 VPWR VGND sg13g2_nand2_1
XFILLER_37_793 VPWR VGND sg13g2_decap_8
XFILLER_24_454 VPWR VGND sg13g2_decap_8
XFILLER_12_616 VPWR VGND sg13g2_decap_8
XFILLER_25_988 VPWR VGND sg13g2_decap_8
XFILLER_40_947 VPWR VGND sg13g2_decap_8
XFILLER_20_682 VPWR VGND sg13g2_decap_8
XFILLER_22_66 VPWR VGND sg13g2_fill_1
XFILLER_4_837 VPWR VGND sg13g2_decap_8
XFILLER_47_557 VPWR VGND sg13g2_decap_8
XFILLER_43_763 VPWR VGND sg13g2_decap_8
XFILLER_16_955 VPWR VGND sg13g2_decap_8
XFILLER_31_969 VPWR VGND sg13g2_decap_8
XFILLER_7_642 VPWR VGND sg13g2_decap_8
XFILLER_11_671 VPWR VGND sg13g2_decap_8
XFILLER_6_163 VPWR VGND sg13g2_fill_2
X_3370_ net591 net589 _0897_ VPWR VGND sg13g2_nor2_1
X_2321_ net725 VPWR _1741_ VGND net740 _1740_ sg13g2_o21ai_1
X_2252_ _1672_ net757 _1671_ VPWR VGND sg13g2_nand2_1
XFILLER_33_4 VPWR VGND sg13g2_fill_2
XFILLER_38_513 VPWR VGND sg13g2_decap_8
X_2183_ _1511_ _1590_ _1603_ VPWR VGND net772 sg13g2_nand3b_1
XFILLER_46_590 VPWR VGND sg13g2_decap_8
Xclkbuf_5_23__f_sap_3_inst.alu.clk_regs clknet_4_11_0_sap_3_inst.alu.clk_regs clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_34_752 VPWR VGND sg13g2_decap_8
XFILLER_22_958 VPWR VGND sg13g2_decap_8
X_3706_ _1189_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] net579 _0110_
+ VPWR VGND sg13g2_mux2_1
XFILLER_49_1009 VPWR VGND sg13g2_decap_8
X_3637_ _1072_ _1121_ _1134_ VPWR VGND sg13g2_nor2_1
X_3568_ _0808_ net713 _1080_ VPWR VGND sg13g2_nor2_1
XFILLER_1_829 VPWR VGND sg13g2_decap_8
X_2519_ _1921_ _1924_ _1920_ net21 VPWR VGND _1932_ sg13g2_nand4_1
X_3499_ _0072_ _1018_ _1020_ net587 _1484_ VPWR VGND sg13g2_a22oi_1
XFILLER_29_524 VPWR VGND sg13g2_decap_8
XFILLER_44_505 VPWR VGND sg13g2_decap_8
XFILLER_37_590 VPWR VGND sg13g2_decap_8
XFILLER_13_914 VPWR VGND sg13g2_decap_8
XFILLER_24_262 VPWR VGND sg13g2_fill_2
XFILLER_25_785 VPWR VGND sg13g2_decap_8
XFILLER_40_744 VPWR VGND sg13g2_decap_8
XFILLER_21_991 VPWR VGND sg13g2_decap_8
XFILLER_4_634 VPWR VGND sg13g2_decap_8
XFILLER_48_822 VPWR VGND sg13g2_decap_8
Xhold6 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[1\] VPWR VGND net55 sg13g2_dlygate4sd3_1
XFILLER_47_354 VPWR VGND sg13g2_decap_8
XFILLER_48_899 VPWR VGND sg13g2_decap_8
XFILLER_16_752 VPWR VGND sg13g2_decap_8
XFILLER_35_549 VPWR VGND sg13g2_decap_8
XFILLER_43_560 VPWR VGND sg13g2_decap_8
X_2870_ _0428_ _0400_ _0425_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_766 VPWR VGND sg13g2_decap_8
XFILLER_12_980 VPWR VGND sg13g2_decap_8
X_3422_ _0069_ _0935_ _0941_ net586 _1446_ VPWR VGND sg13g2_a22oi_1
X_3353_ _0875_ _0878_ net621 _0880_ VPWR VGND _0879_ sg13g2_nand4_1
X_2304_ VGND VPWR _1724_ _1612_ _1608_ sg13g2_or2_1
X_3284_ _1620_ _0676_ net749 _0812_ VPWR VGND sg13g2_nand3_1
X_2235_ VPWR _1655_ _1654_ VGND sg13g2_inv_1
X_2166_ _1526_ _1528_ _1562_ _1583_ _1586_ VPWR VGND sg13g2_and4_1
XFILLER_39_866 VPWR VGND sg13g2_decap_8
XFILLER_0_1011 VPWR VGND sg13g2_decap_8
XFILLER_26_527 VPWR VGND sg13g2_decap_8
X_2097_ _1517_ _1514_ VPWR VGND net766 sg13g2_nand2b_2
XFILLER_10_928 VPWR VGND sg13g2_decap_8
XFILLER_22_755 VPWR VGND sg13g2_decap_8
X_2999_ _0553_ _0516_ _0552_ VPWR VGND sg13g2_xnor2_1
XFILLER_1_626 VPWR VGND sg13g2_decap_8
X_4038__3 VPWR net39 clknet_leaf_1_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_45_858 VPWR VGND sg13g2_decap_8
XFILLER_44_379 VPWR VGND sg13g2_decap_8
XFILLER_13_711 VPWR VGND sg13g2_decap_8
XFILLER_25_582 VPWR VGND sg13g2_decap_8
XFILLER_40_541 VPWR VGND sg13g2_decap_8
XFILLER_13_788 VPWR VGND sg13g2_decap_8
XFILLER_5_910 VPWR VGND sg13g2_decap_8
XFILLER_5_987 VPWR VGND sg13g2_decap_8
X_2020_ sap_3_inst.controller.opcode\[4\] _1442_ VPWR VGND sg13g2_inv_4
XFILLER_48_696 VPWR VGND sg13g2_decap_8
XFILLER_35_302 VPWR VGND sg13g2_fill_1
XFILLER_36_836 VPWR VGND sg13g2_decap_8
X_3971_ net724 _0301_ _0303_ _1388_ VPWR VGND sg13g2_nor3_1
XFILLER_23_519 VPWR VGND sg13g2_decap_8
X_2922_ _0478_ net793 net720 VPWR VGND sg13g2_nand2_1
XFILLER_31_563 VPWR VGND sg13g2_decap_8
X_2853_ net580 net801 _0411_ _0035_ VPWR VGND sg13g2_a21o_1
X_2784_ _0345_ _0344_ _0322_ VPWR VGND sg13g2_nand2b_1
X_3405_ _0930_ _0925_ _0929_ net671 _1446_ VPWR VGND sg13g2_a22oi_1
Xfanout705 net706 net705 VPWR VGND sg13g2_buf_8
Xfanout749 _1600_ net749 VPWR VGND sg13g2_buf_8
Xfanout727 _1678_ net727 VPWR VGND sg13g2_buf_8
X_3336_ VGND VPWR net730 net726 _0864_ net753 sg13g2_a21oi_1
Xfanout738 net739 net738 VPWR VGND sg13g2_buf_8
Xfanout716 _0593_ net716 VPWR VGND sg13g2_buf_1
X_3267_ net697 net692 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] _0795_
+ VPWR VGND net688 sg13g2_nand4_1
XFILLER_39_663 VPWR VGND sg13g2_decap_8
X_3198_ _0726_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] net670 VPWR
+ VGND sg13g2_nand2_1
X_2218_ net758 net746 _1638_ VPWR VGND sg13g2_and2_1
XFILLER_26_302 VPWR VGND sg13g2_fill_2
X_2149_ _1569_ _1528_ _1562_ _1568_ VPWR VGND sg13g2_and3_2
XFILLER_26_324 VPWR VGND sg13g2_decap_4
XFILLER_27_847 VPWR VGND sg13g2_decap_8
XFILLER_42_828 VPWR VGND sg13g2_decap_8
XFILLER_22_552 VPWR VGND sg13g2_decap_8
XFILLER_10_725 VPWR VGND sg13g2_decap_8
XFILLER_2_924 VPWR VGND sg13g2_decap_8
XFILLER_7_1006 VPWR VGND sg13g2_decap_8
XFILLER_49_449 VPWR VGND sg13g2_decap_8
XFILLER_45_655 VPWR VGND sg13g2_decap_8
XFILLER_18_847 VPWR VGND sg13g2_decap_8
XFILLER_26_891 VPWR VGND sg13g2_decap_8
XFILLER_41_861 VPWR VGND sg13g2_decap_8
XFILLER_13_585 VPWR VGND sg13g2_decap_8
XFILLER_9_567 VPWR VGND sg13g2_decap_8
XFILLER_5_784 VPWR VGND sg13g2_decap_8
XFILLER_45_1012 VPWR VGND sg13g2_decap_8
X_4170_ net829 VGND VPWR _0134_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\]
+ clknet_5_25__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3121_ _1512_ _1591_ _1593_ net727 _0649_ VPWR VGND sg13g2_nor4_1
XFILLER_1_990 VPWR VGND sg13g2_decap_8
X_3052_ VGND VPWR _0227_ net715 _0051_ _0594_ sg13g2_a21oi_1
XFILLER_48_493 VPWR VGND sg13g2_decap_8
XFILLER_35_121 VPWR VGND sg13g2_fill_2
XFILLER_36_633 VPWR VGND sg13g2_decap_8
Xclkbuf_4_13_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_13_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_23_316 VPWR VGND sg13g2_fill_1
XFILLER_24_839 VPWR VGND sg13g2_decap_8
X_3954_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] _1379_
+ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] _1380_ net810 sg13g2_a221oi_1
X_2905_ _0452_ _0461_ _0462_ VPWR VGND sg13g2_nor2_1
X_3885_ _1318_ net809 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] _1300_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2836_ _0393_ _0394_ _0395_ VPWR VGND sg13g2_nor2_1
X_2767_ VGND VPWR _0328_ _0319_ _0201_ sg13g2_or2_1
X_2698_ VGND VPWR net745 _1712_ _0281_ _1834_ sg13g2_a21oi_1
X_3319_ _0847_ _0710_ _0846_ VPWR VGND sg13g2_xnor2_1
Xfanout579 _1174_ net579 VPWR VGND sg13g2_buf_8
XFILLER_46_408 VPWR VGND sg13g2_decap_8
XFILLER_39_460 VPWR VGND sg13g2_decap_8
XFILLER_27_644 VPWR VGND sg13g2_decap_8
XFILLER_42_625 VPWR VGND sg13g2_decap_8
XFILLER_14_338 VPWR VGND sg13g2_fill_2
XFILLER_23_883 VPWR VGND sg13g2_decap_8
XFILLER_10_522 VPWR VGND sg13g2_decap_8
XFILLER_6_537 VPWR VGND sg13g2_decap_8
XFILLER_10_599 VPWR VGND sg13g2_decap_8
XFILLER_2_721 VPWR VGND sg13g2_decap_8
XFILLER_29_1007 VPWR VGND sg13g2_decap_8
XFILLER_2_798 VPWR VGND sg13g2_decap_8
XFILLER_18_644 VPWR VGND sg13g2_decap_8
XFILLER_46_975 VPWR VGND sg13g2_decap_8
XFILLER_45_452 VPWR VGND sg13g2_decap_8
XFILLER_21_809 VPWR VGND sg13g2_decap_8
XFILLER_33_658 VPWR VGND sg13g2_decap_8
X_3670_ _1157_ VPWR _0103_ VGND _0996_ _1160_ sg13g2_o21ai_1
Xclkbuf_4_5_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_5_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_40_190 VPWR VGND sg13g2_fill_1
XFILLER_12_1022 VPWR VGND sg13g2_decap_8
X_2621_ _0210_ net636 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] net642
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2552_ _1964_ net630 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] net639
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_581 VPWR VGND sg13g2_decap_8
X_4222_ net835 VGND VPWR net813 u_ser.state\[0\] clknet_3_1__leaf_clk sg13g2_dfrbpq_2
X_2483_ _1890_ _1898_ _1899_ VPWR VGND sg13g2_nor2_1
X_4153_ net821 VGND VPWR _0117_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\]
+ clknet_5_7__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_909 VPWR VGND sg13g2_decap_8
X_4084_ net840 VGND VPWR _0048_ sap_3_inst.out\[7\] clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3104_ VGND VPWR _1576_ _1753_ _0632_ _0626_ sg13g2_a21oi_1
X_3035_ net787 sap_3_inst.alu.tmp\[7\] _0580_ VPWR VGND sg13g2_nor2b_1
XFILLER_48_290 VPWR VGND sg13g2_decap_8
XFILLER_37_975 VPWR VGND sg13g2_decap_8
XFILLER_24_636 VPWR VGND sg13g2_decap_8
X_3937_ VPWR VGND _1364_ net812 _1359_ _1480_ _1365_ net807 sg13g2_a221oi_1
XFILLER_20_864 VPWR VGND sg13g2_decap_8
X_3868_ sap_3_inst.reg_file.array_serializer_inst.word_index\[1\] sap_3_inst.reg_file.array_serializer_inst.word_index\[0\]
+ _1298_ _1301_ VPWR VGND sg13g2_nor3_2
X_2819_ _0378_ VPWR _0379_ VGND net574 _0377_ sg13g2_o21ai_1
X_3799_ VGND VPWR net661 _1129_ _0140_ _1252_ sg13g2_a21oi_1
XFILLER_47_739 VPWR VGND sg13g2_decap_8
XFILLER_46_249 VPWR VGND sg13g2_fill_1
XFILLER_28_931 VPWR VGND sg13g2_decap_8
XFILLER_27_441 VPWR VGND sg13g2_decap_8
XFILLER_43_945 VPWR VGND sg13g2_decap_8
XFILLER_42_422 VPWR VGND sg13g2_decap_8
XFILLER_15_658 VPWR VGND sg13g2_decap_8
XFILLER_35_1011 VPWR VGND sg13g2_decap_8
XFILLER_42_499 VPWR VGND sg13g2_decap_8
XFILLER_23_680 VPWR VGND sg13g2_decap_8
XFILLER_30_639 VPWR VGND sg13g2_decap_8
XFILLER_7_824 VPWR VGND sg13g2_decap_8
XFILLER_11_853 VPWR VGND sg13g2_decap_8
XFILLER_2_595 VPWR VGND sg13g2_decap_8
XFILLER_19_920 VPWR VGND sg13g2_decap_8
XFILLER_46_772 VPWR VGND sg13g2_decap_8
XFILLER_45_260 VPWR VGND sg13g2_fill_2
XFILLER_19_997 VPWR VGND sg13g2_decap_8
XFILLER_34_934 VPWR VGND sg13g2_decap_8
XFILLER_21_606 VPWR VGND sg13g2_decap_8
X_3722_ _0115_ _1085_ _1200_ net617 _1463_ VPWR VGND sg13g2_a22oi_1
X_3653_ _1093_ _1146_ _1147_ VPWR VGND sg13g2_nor2_2
X_2604_ net801 net800 _2013_ VPWR VGND sg13g2_xor2_1
X_3584_ _1093_ VPWR _1094_ VGND net668 _0921_ sg13g2_o21ai_1
X_2535_ net745 _1786_ _1947_ VPWR VGND sg13g2_and2_1
X_2466_ _1884_ _1882_ _1883_ VPWR VGND sg13g2_nand2_1
X_4205_ net844 VGND VPWR _0169_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2397_ _1817_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] net645
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4136_ net833 VGND VPWR _0100_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\]
+ clknet_5_28__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_205 VPWR VGND sg13g2_fill_2
XFILLER_29_706 VPWR VGND sg13g2_decap_8
X_4067_ net834 VGND VPWR _0031_ sap_3_inst.alu.flags\[6\] net48 sg13g2_dfrbpq_1
X_3018_ _0570_ VPWR _0041_ VGND _1459_ net717 sg13g2_o21ai_1
XFILLER_37_772 VPWR VGND sg13g2_decap_8
XFILLER_24_433 VPWR VGND sg13g2_decap_8
XFILLER_25_967 VPWR VGND sg13g2_decap_8
XFILLER_40_926 VPWR VGND sg13g2_decap_8
XFILLER_11_138 VPWR VGND sg13g2_fill_1
XFILLER_20_661 VPWR VGND sg13g2_decap_8
XFILLER_4_816 VPWR VGND sg13g2_decap_8
XFILLER_3_348 VPWR VGND sg13g2_fill_2
XFILLER_47_536 VPWR VGND sg13g2_decap_8
XFILLER_16_934 VPWR VGND sg13g2_decap_8
XFILLER_27_271 VPWR VGND sg13g2_fill_2
XFILLER_43_742 VPWR VGND sg13g2_decap_8
XFILLER_42_252 VPWR VGND sg13g2_fill_1
XFILLER_31_948 VPWR VGND sg13g2_decap_8
XFILLER_8_58 VPWR VGND sg13g2_fill_2
XFILLER_11_650 VPWR VGND sg13g2_decap_8
XFILLER_7_621 VPWR VGND sg13g2_decap_8
XFILLER_7_698 VPWR VGND sg13g2_decap_8
XFILLER_6_197 VPWR VGND sg13g2_fill_2
X_2320_ _1740_ net781 _1584_ VPWR VGND sg13g2_nand2_2
X_2251_ _1539_ VPWR _1671_ VGND _1544_ _1670_ sg13g2_o21ai_1
X_2182_ net773 _1512_ _1591_ _1602_ VPWR VGND sg13g2_nor3_1
XFILLER_26_709 VPWR VGND sg13g2_decap_8
XFILLER_38_569 VPWR VGND sg13g2_decap_8
XFILLER_19_794 VPWR VGND sg13g2_decap_8
XFILLER_34_731 VPWR VGND sg13g2_decap_8
XFILLER_22_937 VPWR VGND sg13g2_decap_8
X_3705_ VGND VPWR _1189_ _1188_ _1187_ sg13g2_or2_1
X_3636_ _0096_ _1133_ _1065_ _1121_ _1491_ VPWR VGND sg13g2_a22oi_1
XFILLER_1_808 VPWR VGND sg13g2_decap_8
X_3567_ _1076_ net31 _1078_ _1079_ VPWR VGND sg13g2_a21o_1
X_2518_ net576 VPWR _1932_ VGND _1927_ _1931_ sg13g2_o21ai_1
X_3498_ net587 _1011_ _1019_ _1020_ VPWR VGND sg13g2_nor3_1
X_2449_ _1569_ net728 net765 _1868_ VPWR VGND sg13g2_nand3_1
XFILLER_29_503 VPWR VGND sg13g2_decap_8
X_4119_ net819 VGND VPWR _0083_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_25_764 VPWR VGND sg13g2_decap_8
XFILLER_40_723 VPWR VGND sg13g2_decap_8
XFILLER_33_77 VPWR VGND sg13g2_fill_1
XFILLER_21_970 VPWR VGND sg13g2_decap_8
XFILLER_32_1014 VPWR VGND sg13g2_decap_8
XFILLER_4_613 VPWR VGND sg13g2_decap_8
XFILLER_48_801 VPWR VGND sg13g2_decap_8
XFILLER_0_885 VPWR VGND sg13g2_decap_8
Xhold7 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\] VPWR VGND net56 sg13g2_dlygate4sd3_1
XFILLER_48_878 VPWR VGND sg13g2_decap_8
XFILLER_47_333 VPWR VGND sg13g2_decap_8
XFILLER_35_528 VPWR VGND sg13g2_decap_8
XFILLER_16_731 VPWR VGND sg13g2_decap_8
XFILLER_31_745 VPWR VGND sg13g2_decap_8
XFILLER_30_244 VPWR VGND sg13g2_fill_1
XFILLER_8_985 VPWR VGND sg13g2_decap_8
XFILLER_7_495 VPWR VGND sg13g2_decap_8
X_3421_ _0946_ _0945_ _0944_ VPWR VGND sg13g2_nand2b_1
X_3352_ _0879_ net655 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] net674
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2303_ _1673_ _1722_ _1538_ _1723_ VPWR VGND sg13g2_nand3_1
X_3283_ _0810_ _0809_ _0670_ _0811_ VPWR VGND sg13g2_a21o_1
X_2234_ _1654_ _1642_ net758 net746 net755 VPWR VGND sg13g2_a22oi_1
XFILLER_39_845 VPWR VGND sg13g2_decap_8
X_2165_ _1563_ _1584_ _1585_ VPWR VGND sg13g2_nor2_1
XFILLER_26_506 VPWR VGND sg13g2_decap_8
X_2096_ net766 _1515_ _1516_ VPWR VGND sg13g2_nor2_2
XFILLER_19_591 VPWR VGND sg13g2_decap_8
XFILLER_22_734 VPWR VGND sg13g2_decap_8
XFILLER_10_907 VPWR VGND sg13g2_decap_8
X_2998_ _0552_ _0549_ _0551_ VPWR VGND sg13g2_xnor2_1
X_3619_ _1046_ _1047_ _1121_ _1123_ VPWR VGND sg13g2_nor3_1
XFILLER_1_605 VPWR VGND sg13g2_decap_8
XFILLER_0_137 VPWR VGND sg13g2_fill_1
XFILLER_29_311 VPWR VGND sg13g2_decap_4
XFILLER_45_837 VPWR VGND sg13g2_decap_8
XFILLER_44_358 VPWR VGND sg13g2_decap_8
XFILLER_25_561 VPWR VGND sg13g2_decap_8
XFILLER_40_520 VPWR VGND sg13g2_decap_8
XFILLER_13_767 VPWR VGND sg13g2_decap_8
XFILLER_40_597 VPWR VGND sg13g2_decap_8
XFILLER_9_749 VPWR VGND sg13g2_decap_8
XFILLER_5_966 VPWR VGND sg13g2_decap_8
XFILLER_4_487 VPWR VGND sg13g2_decap_8
XFILLER_0_682 VPWR VGND sg13g2_decap_8
XFILLER_48_675 VPWR VGND sg13g2_decap_8
XFILLER_47_152 VPWR VGND sg13g2_fill_1
XFILLER_36_815 VPWR VGND sg13g2_decap_8
X_3970_ _1386_ VPWR _0176_ VGND _1196_ _1387_ sg13g2_o21ai_1
X_2921_ VGND VPWR net796 net720 _0477_ _0448_ sg13g2_a21oi_1
XFILLER_31_542 VPWR VGND sg13g2_decap_8
X_2852_ VPWR VGND _0410_ net580 _0409_ _2008_ _0411_ net626 sg13g2_a221oi_1
X_2783_ net775 _1951_ _1956_ _0344_ VPWR VGND sg13g2_nor3_2
XFILLER_8_782 VPWR VGND sg13g2_decap_8
XFILLER_7_292 VPWR VGND sg13g2_fill_2
X_3404_ _0929_ _0926_ _0927_ _0928_ VPWR VGND sg13g2_and3_1
Xfanout706 _0619_ net706 VPWR VGND sg13g2_buf_2
Xfanout728 _1677_ net728 VPWR VGND sg13g2_buf_8
Xfanout717 net719 net717 VPWR VGND sg13g2_buf_8
Xfanout739 _1533_ net739 VPWR VGND sg13g2_buf_8
X_3335_ _0862_ net597 net621 _0863_ VPWR VGND sg13g2_a21o_1
X_3266_ net703 net697 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] _0794_
+ VPWR VGND net691 sg13g2_nand4_1
X_2217_ VPWR VGND _1581_ _1635_ _1636_ _1607_ _1637_ _1622_ sg13g2_a221oi_1
XFILLER_39_642 VPWR VGND sg13g2_decap_8
X_3197_ _0725_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] net674 VPWR
+ VGND sg13g2_nand2_1
XFILLER_27_826 VPWR VGND sg13g2_decap_8
X_2148_ net782 net785 _1568_ VPWR VGND sg13g2_nor2b_2
X_2079_ VPWR _1501_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_42_807 VPWR VGND sg13g2_decap_8
XFILLER_35_892 VPWR VGND sg13g2_decap_8
XFILLER_22_531 VPWR VGND sg13g2_decap_8
XFILLER_10_704 VPWR VGND sg13g2_decap_8
XFILLER_6_719 VPWR VGND sg13g2_decap_8
XFILLER_5_207 VPWR VGND sg13g2_fill_1
XFILLER_2_903 VPWR VGND sg13g2_decap_8
X_4040__5 VPWR net41 clknet_leaf_0_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_30_67 VPWR VGND sg13g2_fill_1
XFILLER_49_428 VPWR VGND sg13g2_decap_8
XFILLER_1_479 VPWR VGND sg13g2_decap_8
XFILLER_39_87 VPWR VGND sg13g2_fill_1
XFILLER_18_826 VPWR VGND sg13g2_decap_8
XFILLER_45_634 VPWR VGND sg13g2_decap_8
XFILLER_26_870 VPWR VGND sg13g2_decap_8
XFILLER_41_840 VPWR VGND sg13g2_decap_8
XFILLER_13_564 VPWR VGND sg13g2_decap_8
XFILLER_9_546 VPWR VGND sg13g2_decap_8
XFILLER_5_763 VPWR VGND sg13g2_decap_8
XFILLER_4_262 VPWR VGND sg13g2_fill_2
X_3120_ net745 _1514_ net778 _0648_ VPWR VGND net764 sg13g2_nand4_1
XFILLER_49_995 VPWR VGND sg13g2_decap_8
XFILLER_48_472 VPWR VGND sg13g2_decap_8
X_3051_ sap_3_inst.alu.tmp\[1\] net715 _0594_ VPWR VGND sg13g2_nor2_1
XFILLER_36_612 VPWR VGND sg13g2_decap_8
XFILLER_24_818 VPWR VGND sg13g2_decap_8
XFILLER_36_689 VPWR VGND sg13g2_decap_8
X_3953_ _1376_ _1377_ _1374_ _1379_ VPWR VGND _1378_ sg13g2_nand4_1
X_2904_ VGND VPWR net798 _1472_ _0461_ _0433_ sg13g2_a21oi_1
XFILLER_32_895 VPWR VGND sg13g2_decap_8
X_3884_ net815 net816 _1299_ _1317_ VPWR VGND sg13g2_nor3_2
X_2835_ VGND VPWR net805 _0364_ _0394_ _0363_ sg13g2_a21oi_1
X_2766_ VGND VPWR _0327_ _1958_ _1950_ sg13g2_or2_1
X_2697_ _0280_ _1517_ net756 VPWR VGND sg13g2_nand2_1
X_3318_ net591 _0842_ _0846_ VPWR VGND sg13g2_nor2_2
X_3249_ _0776_ VPWR _0777_ VGND _1470_ _0690_ sg13g2_o21ai_1
XFILLER_27_623 VPWR VGND sg13g2_decap_8
XFILLER_42_604 VPWR VGND sg13g2_decap_8
XFILLER_26_155 VPWR VGND sg13g2_fill_1
XFILLER_10_501 VPWR VGND sg13g2_decap_8
XFILLER_23_862 VPWR VGND sg13g2_decap_8
XFILLER_22_394 VPWR VGND sg13g2_fill_2
XFILLER_6_516 VPWR VGND sg13g2_decap_8
XFILLER_10_578 VPWR VGND sg13g2_decap_8
XFILLER_2_700 VPWR VGND sg13g2_decap_8
XFILLER_2_777 VPWR VGND sg13g2_decap_8
XFILLER_2_38 VPWR VGND sg13g2_decap_8
XFILLER_46_954 VPWR VGND sg13g2_decap_8
XFILLER_18_623 VPWR VGND sg13g2_decap_8
XFILLER_45_431 VPWR VGND sg13g2_decap_8
XFILLER_33_637 VPWR VGND sg13g2_decap_8
XFILLER_17_199 VPWR VGND sg13g2_fill_2
XFILLER_32_125 VPWR VGND sg13g2_fill_2
XFILLER_32_147 VPWR VGND sg13g2_fill_1
XFILLER_14_884 VPWR VGND sg13g2_decap_8
XFILLER_12_1001 VPWR VGND sg13g2_decap_8
X_2620_ _0209_ net630 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] net639
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2551_ _1963_ net644 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] net646
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2482_ _1895_ _1897_ _1898_ VPWR VGND sg13g2_nor2_1
XFILLER_5_560 VPWR VGND sg13g2_decap_8
X_4221_ net837 VGND VPWR _0184_ sap_3_inst.alu.act\[7\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_4152_ net842 VGND VPWR _0116_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\]
+ clknet_5_29__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3103_ VPWR VGND _1611_ _0610_ _0627_ net775 _0631_ _1823_ sg13g2_a221oi_1
X_4083_ net837 VGND VPWR _0047_ sap_3_inst.out\[6\] clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_49_792 VPWR VGND sg13g2_decap_8
X_3034_ _0327_ _0497_ _0515_ _0552_ _0579_ VPWR VGND sg13g2_nor4_1
XFILLER_37_954 VPWR VGND sg13g2_decap_8
XFILLER_24_615 VPWR VGND sg13g2_decap_8
X_3936_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] _1363_
+ _1306_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] _1364_ _1301_ sg13g2_a221oi_1
XFILLER_20_843 VPWR VGND sg13g2_decap_8
XFILLER_32_692 VPWR VGND sg13g2_decap_8
X_3867_ _1298_ _1299_ _1300_ VPWR VGND sg13g2_nor2_2
XFILLER_31_191 VPWR VGND sg13g2_fill_2
X_2818_ VGND VPWR net574 _0371_ _0378_ net708 sg13g2_a21oi_1
X_3798_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] net661 _1252_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_3_519 VPWR VGND sg13g2_decap_8
X_2749_ _0310_ _1517_ _0307_ VPWR VGND sg13g2_nand2_1
XFILLER_47_718 VPWR VGND sg13g2_decap_8
XFILLER_28_910 VPWR VGND sg13g2_decap_8
XFILLER_43_924 VPWR VGND sg13g2_decap_8
XFILLER_42_401 VPWR VGND sg13g2_decap_8
XFILLER_28_987 VPWR VGND sg13g2_decap_8
XFILLER_15_637 VPWR VGND sg13g2_decap_8
XFILLER_27_497 VPWR VGND sg13g2_decap_8
XFILLER_42_478 VPWR VGND sg13g2_decap_8
XFILLER_30_618 VPWR VGND sg13g2_decap_8
XFILLER_11_832 VPWR VGND sg13g2_decap_8
XFILLER_7_803 VPWR VGND sg13g2_decap_8
Xclkbuf_5_31__f_sap_3_inst.alu.clk_regs clknet_4_15_0_sap_3_inst.alu.clk_regs clknet_5_31__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_2_574 VPWR VGND sg13g2_decap_8
XFILLER_46_751 VPWR VGND sg13g2_decap_8
XFILLER_19_976 VPWR VGND sg13g2_decap_8
XFILLER_34_913 VPWR VGND sg13g2_decap_8
XFILLER_18_497 VPWR VGND sg13g2_decap_8
XFILLER_14_681 VPWR VGND sg13g2_decap_8
XFILLER_20_106 VPWR VGND sg13g2_fill_2
XFILLER_9_151 VPWR VGND sg13g2_fill_1
XFILLER_9_140 VPWR VGND sg13g2_fill_2
X_3721_ net18 net617 _1200_ VPWR VGND sg13g2_nor2_1
XFILLER_9_184 VPWR VGND sg13g2_fill_1
X_3652_ net599 _0909_ _1146_ VPWR VGND sg13g2_nor2_1
X_2603_ net805 net803 _2012_ VPWR VGND sg13g2_xor2_1
X_3583_ net605 _0914_ _1093_ VPWR VGND sg13g2_nor2_1
XFILLER_6_880 VPWR VGND sg13g2_decap_8
X_2534_ _1946_ _1868_ _1945_ VPWR VGND sg13g2_nand2_2
X_2465_ _1883_ net637 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] net638
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2396_ _1816_ net638 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] net640
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4204_ net848 VGND VPWR _0168_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[7\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_3_81 VPWR VGND sg13g2_fill_1
X_4135_ net819 VGND VPWR _0099_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4066_ net838 VGND VPWR _0030_ sap_3_inst.alu.flags\[5\] net47 sg13g2_dfrbpq_1
XFILLER_37_751 VPWR VGND sg13g2_decap_8
X_3017_ _0570_ sap_3_inst.out\[0\] net717 VPWR VGND sg13g2_nand2_1
XFILLER_24_412 VPWR VGND sg13g2_decap_8
XFILLER_19_1018 VPWR VGND sg13g2_decap_8
XFILLER_25_946 VPWR VGND sg13g2_decap_8
XFILLER_40_905 VPWR VGND sg13g2_decap_8
XFILLER_24_489 VPWR VGND sg13g2_decap_8
XFILLER_20_640 VPWR VGND sg13g2_decap_8
X_3919_ VPWR VGND _1348_ net812 _1344_ _1446_ _1349_ net807 sg13g2_a221oi_1
XFILLER_47_515 VPWR VGND sg13g2_decap_8
XFILLER_16_913 VPWR VGND sg13g2_decap_8
XFILLER_28_784 VPWR VGND sg13g2_decap_8
XFILLER_43_721 VPWR VGND sg13g2_decap_8
XFILLER_31_927 VPWR VGND sg13g2_decap_8
XFILLER_43_798 VPWR VGND sg13g2_decap_8
XFILLER_7_600 VPWR VGND sg13g2_decap_8
XFILLER_6_110 VPWR VGND sg13g2_fill_2
XFILLER_10_194 VPWR VGND sg13g2_fill_2
XFILLER_7_677 VPWR VGND sg13g2_decap_8
XFILLER_6_165 VPWR VGND sg13g2_fill_1
XFILLER_3_883 VPWR VGND sg13g2_decap_8
X_2250_ VGND VPWR _1567_ _1669_ _1670_ _1556_ sg13g2_a21oi_1
X_2181_ _1598_ net749 net751 _1601_ VPWR VGND sg13g2_nand3_1
XFILLER_38_548 VPWR VGND sg13g2_decap_8
XFILLER_19_773 VPWR VGND sg13g2_decap_8
XFILLER_34_710 VPWR VGND sg13g2_decap_8
XFILLER_22_916 VPWR VGND sg13g2_decap_8
XFILLER_34_787 VPWR VGND sg13g2_decap_8
XFILLER_30_982 VPWR VGND sg13g2_decap_8
X_3704_ net598 _0958_ _1188_ VPWR VGND sg13g2_nor2_1
X_3635_ _1121_ _1132_ _1133_ VPWR VGND sg13g2_nor2_1
X_3566_ VGND VPWR _0829_ _1076_ _1078_ _1077_ sg13g2_a21oi_1
X_2517_ _1929_ _1930_ _1928_ _1931_ VPWR VGND sg13g2_nand3_1
X_3497_ net15 net33 net595 _1019_ VPWR VGND sg13g2_mux2_1
X_2448_ net763 _1570_ _1678_ _1867_ VPWR VGND sg13g2_nor3_2
X_2379_ _1799_ _1795_ _1797_ VPWR VGND sg13g2_nand2_2
XFILLER_29_559 VPWR VGND sg13g2_decap_8
X_4118_ net843 VGND VPWR _0082_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4049_ net831 VGND VPWR _0017_ u_ser.shadow_reg\[0\] clknet_3_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_25_743 VPWR VGND sg13g2_decap_8
XFILLER_40_702 VPWR VGND sg13g2_decap_8
XFILLER_12_404 VPWR VGND sg13g2_fill_2
XFILLER_13_949 VPWR VGND sg13g2_decap_8
XFILLER_24_264 VPWR VGND sg13g2_fill_1
XFILLER_40_779 VPWR VGND sg13g2_decap_8
XFILLER_3_113 VPWR VGND sg13g2_fill_1
XFILLER_4_669 VPWR VGND sg13g2_decap_8
XFILLER_3_146 VPWR VGND sg13g2_fill_2
XFILLER_0_864 VPWR VGND sg13g2_decap_8
XFILLER_47_312 VPWR VGND sg13g2_decap_8
Xhold8 _0157_ VPWR VGND net57 sg13g2_dlygate4sd3_1
XFILLER_48_857 VPWR VGND sg13g2_decap_8
XFILLER_47_389 VPWR VGND sg13g2_decap_8
XFILLER_16_710 VPWR VGND sg13g2_decap_8
XFILLER_35_507 VPWR VGND sg13g2_decap_8
XFILLER_28_581 VPWR VGND sg13g2_decap_8
XFILLER_43_595 VPWR VGND sg13g2_decap_8
XFILLER_16_787 VPWR VGND sg13g2_decap_8
XFILLER_31_724 VPWR VGND sg13g2_decap_8
XFILLER_8_964 VPWR VGND sg13g2_decap_8
XFILLER_48_1011 VPWR VGND sg13g2_decap_8
X_3420_ _0766_ VPWR _0945_ VGND net592 _0835_ sg13g2_o21ai_1
Xclkbuf_5_28__f_sap_3_inst.alu.clk_regs clknet_4_14_0_sap_3_inst.alu.clk_regs clknet_5_28__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3351_ _0878_ net665 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] net680
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_3_680 VPWR VGND sg13g2_decap_8
X_2302_ net757 VPWR _1722_ VGND _1679_ _1721_ sg13g2_o21ai_1
X_3282_ net735 VPWR _0810_ VGND _1586_ _1613_ sg13g2_o21ai_1
X_2233_ _1653_ _1639_ _1573_ net753 _1587_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_824 VPWR VGND sg13g2_decap_8
X_2164_ _1584_ net786 net783 VPWR VGND sg13g2_nand2_2
X_2095_ _1515_ net771 VPWR VGND net769 sg13g2_nand2b_2
XFILLER_19_570 VPWR VGND sg13g2_decap_8
XFILLER_22_713 VPWR VGND sg13g2_decap_8
XFILLER_34_584 VPWR VGND sg13g2_decap_8
XFILLER_21_223 VPWR VGND sg13g2_decap_8
X_2997_ VGND VPWR _0511_ _0514_ _0551_ _0550_ sg13g2_a21oi_1
XFILLER_21_278 VPWR VGND sg13g2_fill_1
X_3618_ _1122_ _0690_ _1076_ VPWR VGND sg13g2_nand2_2
X_3549_ _0079_ _1061_ _1063_ net584 _1483_ VPWR VGND sg13g2_a22oi_1
XFILLER_28_56 VPWR VGND sg13g2_fill_1
XFILLER_45_816 VPWR VGND sg13g2_decap_8
XFILLER_17_529 VPWR VGND sg13g2_decap_8
XFILLER_25_540 VPWR VGND sg13g2_decap_8
XFILLER_13_746 VPWR VGND sg13g2_decap_8
XFILLER_40_576 VPWR VGND sg13g2_decap_8
XFILLER_8_227 VPWR VGND sg13g2_fill_2
XFILLER_9_728 VPWR VGND sg13g2_decap_8
XFILLER_5_945 VPWR VGND sg13g2_decap_8
XFILLER_5_38 VPWR VGND sg13g2_decap_8
XFILLER_0_661 VPWR VGND sg13g2_decap_8
XFILLER_48_654 VPWR VGND sg13g2_decap_8
XFILLER_10_8 VPWR VGND sg13g2_fill_2
XFILLER_16_584 VPWR VGND sg13g2_decap_8
X_2920_ net573 net627 _0476_ VPWR VGND sg13g2_nor2b_1
XFILLER_43_392 VPWR VGND sg13g2_decap_8
XFILLER_31_521 VPWR VGND sg13g2_decap_8
X_2851_ VGND VPWR sap_3_inst.alu.act\[2\] net708 _0410_ net626 sg13g2_a21oi_1
X_2782_ _0342_ VPWR _0343_ VGND net806 sap_3_inst.alu.tmp\[0\] sg13g2_o21ai_1
XFILLER_31_598 VPWR VGND sg13g2_decap_8
XFILLER_8_761 VPWR VGND sg13g2_decap_8
X_3403_ _0928_ net675 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] net680
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] VPWR VGND sg13g2_a22oi_1
Xfanout718 net719 net718 VPWR VGND sg13g2_buf_2
Xfanout729 _1677_ net729 VPWR VGND sg13g2_buf_8
Xfanout707 _0314_ net707 VPWR VGND sg13g2_buf_8
X_3334_ _0862_ _0861_ VPWR VGND _0641_ sg13g2_nand2b_2
X_3265_ net703 net690 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] _0793_
+ VPWR VGND sg13g2_nand3_1
X_2216_ _1636_ _1573_ net730 VPWR VGND sg13g2_nand2_1
XFILLER_22_1014 VPWR VGND sg13g2_decap_8
XFILLER_39_621 VPWR VGND sg13g2_decap_8
X_3196_ _0723_ VPWR _0724_ VGND _1491_ net619 sg13g2_o21ai_1
XFILLER_26_304 VPWR VGND sg13g2_fill_1
XFILLER_27_805 VPWR VGND sg13g2_decap_8
X_2147_ VPWR VGND _1561_ net736 _1566_ net744 _1567_ _1565_ sg13g2_a221oi_1
XFILLER_39_698 VPWR VGND sg13g2_decap_8
X_2078_ VPWR _1500_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_22_510 VPWR VGND sg13g2_decap_8
XFILLER_34_370 VPWR VGND sg13g2_fill_1
XFILLER_35_871 VPWR VGND sg13g2_decap_8
XFILLER_22_587 VPWR VGND sg13g2_decap_8
XFILLER_2_959 VPWR VGND sg13g2_decap_8
XFILLER_49_407 VPWR VGND sg13g2_decap_8
XFILLER_45_613 VPWR VGND sg13g2_decap_8
XFILLER_18_805 VPWR VGND sg13g2_decap_8
XFILLER_33_819 VPWR VGND sg13g2_decap_8
XFILLER_38_1010 VPWR VGND sg13g2_decap_8
XFILLER_13_543 VPWR VGND sg13g2_decap_8
XFILLER_9_525 VPWR VGND sg13g2_decap_8
XFILLER_41_896 VPWR VGND sg13g2_decap_8
XFILLER_5_742 VPWR VGND sg13g2_decap_8
X_3050_ sap_3_inst.alu.tmp\[0\] net31 net715 _0050_ VPWR VGND sg13g2_mux2_1
XFILLER_49_974 VPWR VGND sg13g2_decap_8
XFILLER_48_451 VPWR VGND sg13g2_decap_8
XFILLER_35_123 VPWR VGND sg13g2_fill_1
XFILLER_36_668 VPWR VGND sg13g2_decap_8
XFILLER_17_893 VPWR VGND sg13g2_decap_8
X_3952_ _1378_ _1307_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] _1301_
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3883_ _1298_ _1302_ _1316_ VPWR VGND sg13g2_nor2_2
X_2903_ _0460_ _0427_ _0458_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_874 VPWR VGND sg13g2_decap_8
X_2834_ _0393_ net801 net721 VPWR VGND sg13g2_xnor2_1
X_2765_ _1950_ _1958_ _0326_ VPWR VGND sg13g2_nor2_2
X_2696_ _0279_ _1940_ _0278_ VPWR VGND sg13g2_nand2_1
X_3317_ net591 _0839_ _0845_ VPWR VGND sg13g2_nor2_1
XFILLER_27_602 VPWR VGND sg13g2_decap_8
X_3248_ net704 net702 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] _0776_
+ VPWR VGND net694 sg13g2_nand4_1
XFILLER_39_495 VPWR VGND sg13g2_decap_8
X_3179_ _0707_ net657 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] net681
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_15_819 VPWR VGND sg13g2_decap_8
XFILLER_27_679 VPWR VGND sg13g2_decap_8
XFILLER_23_841 VPWR VGND sg13g2_decap_8
XFILLER_10_557 VPWR VGND sg13g2_decap_8
XFILLER_2_756 VPWR VGND sg13g2_decap_8
XFILLER_18_602 VPWR VGND sg13g2_decap_8
XFILLER_46_933 VPWR VGND sg13g2_decap_8
XFILLER_45_410 VPWR VGND sg13g2_decap_8
XFILLER_45_487 VPWR VGND sg13g2_decap_8
XFILLER_18_679 VPWR VGND sg13g2_decap_8
XFILLER_33_616 VPWR VGND sg13g2_decap_8
XFILLER_14_863 VPWR VGND sg13g2_decap_8
XFILLER_41_693 VPWR VGND sg13g2_decap_8
X_2550_ _1962_ sap_3_inst.alu.flags\[3\] _1961_ VPWR VGND sg13g2_nand2_1
X_2481_ _1891_ _1892_ net648 _1897_ VPWR VGND _1896_ sg13g2_nand4_1
X_4220_ net837 VGND VPWR _0183_ sap_3_inst.alu.act\[6\] clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_4151_ net819 VGND VPWR _0115_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\]
+ clknet_5_5__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3102_ _0629_ _0628_ _1442_ _0630_ VPWR VGND sg13g2_a21o_1
X_4082_ net837 VGND VPWR _0046_ sap_3_inst.out\[5\] clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_49_771 VPWR VGND sg13g2_decap_8
X_3033_ VGND VPWR _0328_ _0574_ _0578_ _0577_ sg13g2_a21oi_1
XFILLER_37_933 VPWR VGND sg13g2_decap_8
XFILLER_17_690 VPWR VGND sg13g2_decap_8
X_3935_ _1360_ _1361_ _1358_ _1363_ VPWR VGND _1362_ sg13g2_nand4_1
XFILLER_20_822 VPWR VGND sg13g2_decap_8
XFILLER_32_671 VPWR VGND sg13g2_decap_8
X_3866_ _1299_ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\] VPWR VGND
+ sap_3_inst.reg_file.array_serializer_inst.word_index\[1\] sg13g2_nand2b_2
X_2817_ _0373_ _0374_ _0368_ _0377_ VPWR VGND _0376_ sg13g2_nand4_1
XFILLER_20_899 VPWR VGND sg13g2_decap_8
X_3797_ _1251_ VPWR _0139_ VGND net611 _1176_ sg13g2_o21ai_1
X_2748_ _1713_ _1856_ _0308_ _0309_ VPWR VGND sg13g2_nor3_1
X_2679_ _1613_ VPWR _0262_ VGND net744 _1638_ sg13g2_o21ai_1
Xclkbuf_5_2__f_sap_3_inst.alu.clk_regs clknet_4_1_0_sap_3_inst.alu.clk_regs clknet_5_2__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_36_12 VPWR VGND sg13g2_fill_2
XFILLER_43_903 VPWR VGND sg13g2_decap_8
XFILLER_28_966 VPWR VGND sg13g2_decap_8
XFILLER_15_616 VPWR VGND sg13g2_decap_8
XFILLER_27_476 VPWR VGND sg13g2_decap_8
XFILLER_42_457 VPWR VGND sg13g2_decap_8
XFILLER_11_811 VPWR VGND sg13g2_decap_8
XFILLER_7_859 VPWR VGND sg13g2_decap_8
XFILLER_11_888 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_fill_2
XFILLER_2_553 VPWR VGND sg13g2_decap_8
XFILLER_42_1017 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_730 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_sap_3_inst.alu.clk clknet_1_0__leaf_sap_3_inst.alu.clk clknet_leaf_0_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_19_955 VPWR VGND sg13g2_decap_8
XFILLER_18_454 VPWR VGND sg13g2_fill_2
XFILLER_34_969 VPWR VGND sg13g2_decap_8
X_3720_ net616 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] _1199_ _0114_
+ VPWR VGND sg13g2_a21o_1
XFILLER_14_660 VPWR VGND sg13g2_decap_8
XFILLER_41_490 VPWR VGND sg13g2_decap_8
X_3651_ _0099_ _1085_ _1145_ net623 _1464_ VPWR VGND sg13g2_a22oi_1
X_2602_ _2011_ _2009_ _2010_ VPWR VGND sg13g2_xnor2_1
X_3582_ net600 _0922_ _1091_ _1092_ VPWR VGND sg13g2_nor3_1
X_2533_ VGND VPWR net714 _1945_ _1943_ _1933_ sg13g2_a21oi_2
X_2464_ _1882_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\] net650
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] VPWR VGND sg13g2_a22oi_1
X_4203_ net848 VGND VPWR _0167_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[6\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
X_2395_ _1810_ _1814_ _1815_ VPWR VGND sg13g2_and2_1
XFILLER_3_71 VPWR VGND sg13g2_fill_2
X_4134_ net843 VGND VPWR _0098_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4065_ net834 VGND VPWR _0029_ sap_3_inst.alu.flags\[4\] net46 sg13g2_dfrbpq_1
XFILLER_37_730 VPWR VGND sg13g2_decap_8
X_3016_ _0540_ VPWR _0040_ VGND net581 _0569_ sg13g2_o21ai_1
XFILLER_25_925 VPWR VGND sg13g2_decap_8
XFILLER_36_262 VPWR VGND sg13g2_fill_2
XFILLER_24_468 VPWR VGND sg13g2_decap_8
XFILLER_33_980 VPWR VGND sg13g2_decap_8
X_3918_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] _1347_
+ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] _1348_ _1308_ sg13g2_a221oi_1
X_3849_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\] _1285_ _1286_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_20_696 VPWR VGND sg13g2_decap_8
XFILLER_3_306 VPWR VGND sg13g2_fill_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_43_700 VPWR VGND sg13g2_decap_8
XFILLER_28_763 VPWR VGND sg13g2_decap_8
XFILLER_43_777 VPWR VGND sg13g2_decap_8
XFILLER_16_969 VPWR VGND sg13g2_decap_8
XFILLER_31_906 VPWR VGND sg13g2_decap_8
XFILLER_11_685 VPWR VGND sg13g2_decap_8
XFILLER_7_656 VPWR VGND sg13g2_decap_8
XFILLER_3_862 VPWR VGND sg13g2_decap_8
XFILLER_2_350 VPWR VGND sg13g2_fill_2
X_2180_ _1527_ _1564_ _1580_ _1600_ VPWR VGND sg13g2_or3_1
XFILLER_38_527 VPWR VGND sg13g2_decap_8
XFILLER_19_752 VPWR VGND sg13g2_decap_8
XFILLER_18_262 VPWR VGND sg13g2_fill_2
XFILLER_33_210 VPWR VGND sg13g2_fill_2
XFILLER_34_766 VPWR VGND sg13g2_decap_8
XFILLER_15_980 VPWR VGND sg13g2_decap_8
XFILLER_30_961 VPWR VGND sg13g2_decap_8
X_3703_ _0963_ net607 net32 _1187_ VPWR VGND sg13g2_a21o_1
X_3634_ _1132_ _1064_ _1113_ VPWR VGND sg13g2_nand2_1
X_3565_ net9 _0828_ _1077_ VPWR VGND sg13g2_nor2_1
X_2516_ _1930_ net630 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] net649
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3496_ _1017_ VPWR _1018_ VGND net621 _1014_ sg13g2_o21ai_1
X_2447_ _1820_ _1841_ _1859_ _1866_ net24 VPWR VGND sg13g2_or4_1
XFILLER_25_1023 VPWR VGND sg13g2_decap_4
X_2378_ _1795_ _1797_ _1798_ VPWR VGND sg13g2_and2_1
X_4117_ net828 VGND VPWR _0081_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\]
+ clknet_5_14__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_538 VPWR VGND sg13g2_decap_8
XFILLER_44_519 VPWR VGND sg13g2_decap_8
XFILLER_25_722 VPWR VGND sg13g2_decap_8
XFILLER_13_928 VPWR VGND sg13g2_decap_8
XFILLER_25_799 VPWR VGND sg13g2_decap_8
XFILLER_40_758 VPWR VGND sg13g2_decap_8
XFILLER_4_648 VPWR VGND sg13g2_decap_8
XFILLER_0_843 VPWR VGND sg13g2_decap_8
XFILLER_48_836 VPWR VGND sg13g2_decap_8
Xhold9 u_ser.shadow_reg\[3\] VPWR VGND net58 sg13g2_dlygate4sd3_1
XFILLER_47_368 VPWR VGND sg13g2_decap_8
XFILLER_28_560 VPWR VGND sg13g2_decap_8
XFILLER_16_766 VPWR VGND sg13g2_decap_8
XFILLER_31_703 VPWR VGND sg13g2_decap_8
XFILLER_43_574 VPWR VGND sg13g2_decap_8
XFILLER_15_276 VPWR VGND sg13g2_fill_1
XFILLER_8_943 VPWR VGND sg13g2_decap_8
XFILLER_11_471 VPWR VGND sg13g2_fill_1
XFILLER_12_994 VPWR VGND sg13g2_decap_8
X_3350_ _0876_ VPWR _0877_ VGND _1467_ _0700_ sg13g2_o21ai_1
X_2301_ _1544_ _1719_ _1720_ _1721_ VPWR VGND sg13g2_nor3_1
X_3281_ _0809_ _1608_ _1630_ VPWR VGND sg13g2_nand2_1
XFILLER_39_803 VPWR VGND sg13g2_decap_8
X_2232_ VGND VPWR _1630_ _1650_ _1652_ _1609_ sg13g2_a21oi_1
XFILLER_38_313 VPWR VGND sg13g2_fill_1
X_2163_ net785 net782 _1583_ VPWR VGND sg13g2_and2_1
XFILLER_0_1025 VPWR VGND sg13g2_decap_4
X_2094_ net768 net770 _1514_ VPWR VGND sg13g2_nor2b_2
XFILLER_34_563 VPWR VGND sg13g2_decap_8
XFILLER_22_769 VPWR VGND sg13g2_decap_8
X_2996_ sap_3_inst.alu.tmp\[6\] net791 _0550_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_1_1__f_clk_div_out clknet_0_clk_div_out clknet_1_1__leaf_clk_div_out VPWR
+ VGND sg13g2_buf_8
X_3617_ net674 _1075_ _1121_ VPWR VGND sg13g2_nor2_2
X_3548_ net584 _1062_ _1063_ VPWR VGND sg13g2_nor2_1
X_3479_ _1001_ net621 _1000_ VPWR VGND sg13g2_nand2_1
XFILLER_17_508 VPWR VGND sg13g2_decap_8
XFILLER_38_891 VPWR VGND sg13g2_decap_8
XFILLER_13_725 VPWR VGND sg13g2_decap_8
XFILLER_9_707 VPWR VGND sg13g2_decap_8
XFILLER_25_596 VPWR VGND sg13g2_decap_8
XFILLER_40_555 VPWR VGND sg13g2_decap_8
XFILLER_8_239 VPWR VGND sg13g2_fill_2
XFILLER_5_924 VPWR VGND sg13g2_decap_8
XFILLER_0_640 VPWR VGND sg13g2_decap_8
XFILLER_48_633 VPWR VGND sg13g2_decap_8
XFILLER_44_883 VPWR VGND sg13g2_decap_8
XFILLER_43_371 VPWR VGND sg13g2_decap_8
XFILLER_16_563 VPWR VGND sg13g2_decap_8
XFILLER_31_500 VPWR VGND sg13g2_decap_8
X_2850_ net708 _0407_ _0408_ _0409_ VPWR VGND sg13g2_or3_1
XFILLER_15_1022 VPWR VGND sg13g2_decap_8
XFILLER_31_577 VPWR VGND sg13g2_decap_8
XFILLER_8_740 VPWR VGND sg13g2_decap_8
XFILLER_12_791 VPWR VGND sg13g2_decap_8
X_2781_ _1951_ _0331_ _0342_ VPWR VGND sg13g2_nor2_2
X_3402_ _0927_ net667 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] net678
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] VPWR VGND sg13g2_a22oi_1
Xfanout708 _0314_ net708 VPWR VGND sg13g2_buf_8
Xfanout719 _0267_ net719 VPWR VGND sg13g2_buf_8
X_3333_ _0851_ VPWR _0861_ VGND _0280_ _0860_ sg13g2_o21ai_1
X_3264_ net690 net687 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] _0792_
+ VPWR VGND sg13g2_nand3_1
XFILLER_39_600 VPWR VGND sg13g2_decap_8
X_2215_ VGND VPWR _1630_ _1634_ _1635_ _1619_ sg13g2_a21oi_1
X_3195_ _0723_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] net680 VPWR
+ VGND sg13g2_nand2_1
XFILLER_39_677 VPWR VGND sg13g2_decap_8
X_2146_ net777 net767 net763 _1566_ VGND VPWR _1524_ sg13g2_nor4_2
X_2077_ VPWR _1499_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_35_850 VPWR VGND sg13g2_decap_8
XFILLER_22_566 VPWR VGND sg13g2_decap_8
X_2979_ VGND VPWR _0534_ _0532_ _0530_ sg13g2_or2_1
XFILLER_10_739 VPWR VGND sg13g2_decap_8
XFILLER_2_938 VPWR VGND sg13g2_decap_8
XFILLER_29_154 VPWR VGND sg13g2_fill_2
XFILLER_45_669 VPWR VGND sg13g2_decap_8
XFILLER_13_522 VPWR VGND sg13g2_decap_8
XFILLER_25_393 VPWR VGND sg13g2_decap_8
XFILLER_41_875 VPWR VGND sg13g2_decap_8
XFILLER_9_504 VPWR VGND sg13g2_decap_8
XFILLER_13_599 VPWR VGND sg13g2_decap_8
XFILLER_5_721 VPWR VGND sg13g2_decap_8
XFILLER_5_798 VPWR VGND sg13g2_decap_8
XFILLER_45_1026 VPWR VGND sg13g2_fill_2
XFILLER_49_953 VPWR VGND sg13g2_decap_8
XFILLER_48_430 VPWR VGND sg13g2_decap_8
XFILLER_36_647 VPWR VGND sg13g2_decap_8
XFILLER_17_872 VPWR VGND sg13g2_decap_8
X_3951_ _1377_ _1308_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] _1306_
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_44_680 VPWR VGND sg13g2_decap_8
X_2902_ _0427_ _0458_ _0459_ VPWR VGND sg13g2_nor2_1
XFILLER_32_853 VPWR VGND sg13g2_decap_8
X_3882_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] _1314_
+ _1315_ net808 sg13g2_a21oi_1
X_2833_ _0392_ _0344_ _0382_ VPWR VGND sg13g2_nand2_1
X_2764_ net714 _0324_ _0325_ VPWR VGND sg13g2_nor2b_1
X_2695_ VGND VPWR net737 _1559_ _0278_ _0277_ sg13g2_a21oi_1
X_3316_ _0844_ net590 _0837_ VPWR VGND sg13g2_nand2_1
XFILLER_6_1020 VPWR VGND sg13g2_decap_8
X_3247_ _0771_ _0772_ _0773_ _0774_ _0775_ VPWR VGND sg13g2_and4_1
X_3178_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] net671
+ net662 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] _0706_ net676 sg13g2_a221oi_1
XFILLER_39_474 VPWR VGND sg13g2_decap_8
X_2129_ _1444_ net784 _1524_ _1549_ VPWR VGND sg13g2_nor3_2
XFILLER_27_658 VPWR VGND sg13g2_decap_8
XFILLER_25_36 VPWR VGND sg13g2_fill_1
XFILLER_26_168 VPWR VGND sg13g2_fill_1
XFILLER_42_639 VPWR VGND sg13g2_decap_8
XFILLER_23_820 VPWR VGND sg13g2_decap_8
XFILLER_23_897 VPWR VGND sg13g2_decap_8
XFILLER_10_536 VPWR VGND sg13g2_decap_8
XFILLER_22_396 VPWR VGND sg13g2_fill_1
XFILLER_2_735 VPWR VGND sg13g2_decap_8
XFILLER_46_912 VPWR VGND sg13g2_decap_8
XFILLER_18_658 VPWR VGND sg13g2_decap_8
XFILLER_46_989 VPWR VGND sg13g2_decap_8
XFILLER_45_466 VPWR VGND sg13g2_decap_8
XFILLER_14_842 VPWR VGND sg13g2_decap_8
XFILLER_41_672 VPWR VGND sg13g2_decap_8
XFILLER_40_171 VPWR VGND sg13g2_fill_2
XFILLER_9_378 VPWR VGND sg13g2_fill_2
X_2480_ _1896_ net637 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] net638
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_595 VPWR VGND sg13g2_decap_8
X_4150_ net843 VGND VPWR _0114_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\]
+ clknet_5_26__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3101_ _0629_ _1716_ _1851_ VPWR VGND sg13g2_nand2_1
XFILLER_49_750 VPWR VGND sg13g2_decap_8
X_4081_ net837 VGND VPWR _0045_ sap_3_inst.out\[4\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3032_ VGND VPWR _0485_ _0576_ _0577_ _0575_ sg13g2_a21oi_1
XFILLER_37_912 VPWR VGND sg13g2_decap_8
XFILLER_37_989 VPWR VGND sg13g2_decap_8
X_3934_ _1362_ _1309_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] _1300_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_801 VPWR VGND sg13g2_decap_8
XFILLER_32_650 VPWR VGND sg13g2_decap_8
X_3865_ _1298_ net815 VPWR VGND net816 sg13g2_nand2b_2
X_2816_ VGND VPWR _0326_ _0361_ _0376_ _0375_ sg13g2_a21oi_1
XFILLER_20_878 VPWR VGND sg13g2_decap_8
X_3796_ _1251_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] net611 VPWR
+ VGND sg13g2_nand2_1
X_2747_ net741 _1515_ _1716_ _0308_ VPWR VGND sg13g2_nor3_1
X_2678_ _1618_ VPWR _0261_ VGND net744 _1632_ sg13g2_o21ai_1
XFILLER_28_945 VPWR VGND sg13g2_decap_8
XFILLER_27_455 VPWR VGND sg13g2_decap_8
XFILLER_43_959 VPWR VGND sg13g2_decap_8
XFILLER_42_436 VPWR VGND sg13g2_decap_8
XFILLER_23_694 VPWR VGND sg13g2_decap_8
XFILLER_35_1025 VPWR VGND sg13g2_decap_4
XFILLER_11_867 VPWR VGND sg13g2_decap_8
XFILLER_7_838 VPWR VGND sg13g2_decap_8
XFILLER_2_532 VPWR VGND sg13g2_decap_8
XFILLER_38_709 VPWR VGND sg13g2_decap_8
XFILLER_19_934 VPWR VGND sg13g2_decap_8
XFILLER_46_786 VPWR VGND sg13g2_decap_8
XFILLER_34_948 VPWR VGND sg13g2_decap_8
XFILLER_9_120 VPWR VGND sg13g2_fill_2
X_3650_ net623 _1086_ _1144_ _1145_ VPWR VGND sg13g2_nor3_1
XFILLER_9_197 VPWR VGND sg13g2_fill_1
X_2601_ net797 net795 _2010_ VPWR VGND sg13g2_xor2_1
X_3581_ net19 net11 _1075_ _1091_ VPWR VGND sg13g2_mux2_1
X_2532_ _1933_ _1941_ _1944_ VPWR VGND sg13g2_and2_1
X_2463_ _1881_ _1878_ _1880_ _1858_ net7 VPWR VGND sg13g2_a22oi_1
X_4202_ net848 VGND VPWR _0166_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[5\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
X_2394_ _1814_ net642 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] _1730_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4133_ net829 VGND VPWR _0097_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\]
+ clknet_5_15__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4064_ net821 VGND VPWR _0004_ sap_3_inst.controller.stage\[3\] net45 sg13g2_dfrbpq_2
XFILLER_3_1023 VPWR VGND sg13g2_decap_4
X_3015_ _0569_ _0541_ _0568_ VPWR VGND sg13g2_nand2_1
XFILLER_25_904 VPWR VGND sg13g2_decap_8
XFILLER_37_786 VPWR VGND sg13g2_decap_8
XFILLER_12_609 VPWR VGND sg13g2_decap_8
XFILLER_24_447 VPWR VGND sg13g2_decap_8
X_3917_ _1343_ _1345_ _1342_ _1347_ VPWR VGND _1346_ sg13g2_nand4_1
XFILLER_20_675 VPWR VGND sg13g2_decap_8
X_3848_ _1285_ _1278_ _1279_ VPWR VGND sg13g2_nand2_1
X_3779_ net13 net613 _1238_ _1239_ VPWR VGND sg13g2_nor3_1
XFILLER_28_742 VPWR VGND sg13g2_decap_8
XFILLER_16_948 VPWR VGND sg13g2_decap_8
XFILLER_43_756 VPWR VGND sg13g2_decap_8
XFILLER_23_491 VPWR VGND sg13g2_decap_8
XFILLER_11_664 VPWR VGND sg13g2_decap_8
XFILLER_7_635 VPWR VGND sg13g2_decap_8
XFILLER_10_196 VPWR VGND sg13g2_fill_1
XFILLER_3_841 VPWR VGND sg13g2_decap_8
XFILLER_2_340 VPWR VGND sg13g2_fill_1
XFILLER_38_506 VPWR VGND sg13g2_decap_8
XFILLER_19_731 VPWR VGND sg13g2_decap_8
XFILLER_46_583 VPWR VGND sg13g2_decap_8
XFILLER_34_745 VPWR VGND sg13g2_decap_8
XFILLER_30_940 VPWR VGND sg13g2_decap_8
X_3702_ _1181_ VPWR _0109_ VGND net579 _1186_ sg13g2_o21ai_1
X_3633_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] _1131_ _1122_ _0095_
+ VPWR VGND sg13g2_mux2_1
X_2081__1 VPWR net37 clknet_1_1__leaf_clk_div_out VGND sg13g2_inv_1
X_3564_ _1076_ net667 VPWR VGND net685 sg13g2_nand2b_2
X_3495_ VPWR _1017_ _1016_ VGND sg13g2_inv_1
X_2515_ _1929_ net636 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] net644
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] VPWR VGND sg13g2_a22oi_1
X_2446_ VGND VPWR _1805_ _1865_ _1866_ _1673_ sg13g2_a21oi_1
XFILLER_25_1002 VPWR VGND sg13g2_decap_8
X_4116_ net827 VGND VPWR _0080_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\]
+ clknet_5_9__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2377_ _1797_ _1520_ _1796_ VPWR VGND sg13g2_nand2_1
XFILLER_29_517 VPWR VGND sg13g2_decap_8
XFILLER_25_701 VPWR VGND sg13g2_decap_8
XFILLER_37_583 VPWR VGND sg13g2_decap_8
XFILLER_13_907 VPWR VGND sg13g2_decap_8
XFILLER_40_737 VPWR VGND sg13g2_decap_8
XFILLER_25_778 VPWR VGND sg13g2_decap_8
XFILLER_12_439 VPWR VGND sg13g2_fill_2
XFILLER_21_984 VPWR VGND sg13g2_decap_8
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
XFILLER_4_627 VPWR VGND sg13g2_decap_8
XFILLER_3_148 VPWR VGND sg13g2_fill_1
XFILLER_0_822 VPWR VGND sg13g2_decap_8
XFILLER_48_815 VPWR VGND sg13g2_decap_8
XFILLER_0_899 VPWR VGND sg13g2_decap_8
XFILLER_47_347 VPWR VGND sg13g2_decap_8
XFILLER_43_553 VPWR VGND sg13g2_decap_8
XFILLER_16_745 VPWR VGND sg13g2_decap_8
XFILLER_31_759 VPWR VGND sg13g2_decap_8
XFILLER_8_922 VPWR VGND sg13g2_decap_8
XFILLER_12_973 VPWR VGND sg13g2_decap_8
XFILLER_8_999 VPWR VGND sg13g2_decap_8
X_2300_ net741 _1515_ _1675_ _1720_ VPWR VGND sg13g2_nor3_1
X_3280_ _0808_ _0711_ _0806_ VPWR VGND sg13g2_xnor2_1
X_2231_ _1644_ _1648_ _1651_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_4 VPWR VGND sg13g2_fill_1
X_2162_ net780 _1527_ _1563_ _1580_ _1582_ VPWR VGND sg13g2_or4_1
XFILLER_39_859 VPWR VGND sg13g2_decap_8
X_2093_ net783 net781 _1513_ VPWR VGND net786 sg13g2_nand3b_1
XFILLER_0_1004 VPWR VGND sg13g2_decap_8
XFILLER_46_380 VPWR VGND sg13g2_decap_8
XFILLER_34_542 VPWR VGND sg13g2_decap_8
XFILLER_22_748 VPWR VGND sg13g2_decap_8
X_2995_ _0549_ _0546_ _0548_ VPWR VGND sg13g2_nand2_2
X_3616_ _0089_ _1117_ _1120_ net619 _1500_ VPWR VGND sg13g2_a22oi_1
X_3547_ net599 _0981_ _1062_ VPWR VGND sg13g2_nor2_1
XFILLER_0_107 VPWR VGND sg13g2_fill_2
XFILLER_1_619 VPWR VGND sg13g2_decap_8
X_3478_ _1000_ net664 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] net677
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2429_ _1849_ _1565_ net728 VPWR VGND sg13g2_nand2_1
XFILLER_38_870 VPWR VGND sg13g2_decap_8
XFILLER_13_704 VPWR VGND sg13g2_decap_8
XFILLER_25_575 VPWR VGND sg13g2_decap_8
XFILLER_40_534 VPWR VGND sg13g2_decap_8
XFILLER_12_236 VPWR VGND sg13g2_fill_2
XFILLER_8_229 VPWR VGND sg13g2_fill_1
XFILLER_21_781 VPWR VGND sg13g2_decap_8
XFILLER_5_903 VPWR VGND sg13g2_decap_8
XFILLER_48_612 VPWR VGND sg13g2_decap_8
XFILLER_0_696 VPWR VGND sg13g2_decap_8
XFILLER_48_689 VPWR VGND sg13g2_decap_8
XFILLER_29_881 VPWR VGND sg13g2_decap_8
XFILLER_36_829 VPWR VGND sg13g2_decap_8
XFILLER_16_542 VPWR VGND sg13g2_decap_8
XFILLER_44_862 VPWR VGND sg13g2_decap_8
XFILLER_15_1001 VPWR VGND sg13g2_decap_8
XFILLER_31_556 VPWR VGND sg13g2_decap_8
X_2780_ VGND VPWR net803 net682 _0341_ net708 sg13g2_a21oi_1
XFILLER_12_770 VPWR VGND sg13g2_decap_8
XFILLER_8_796 VPWR VGND sg13g2_decap_8
X_3401_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] net657
+ _0926_ net671 sg13g2_a21oi_1
X_3332_ VGND VPWR _0312_ _0859_ _0860_ _0637_ sg13g2_a21oi_1
Xfanout709 net710 net709 VPWR VGND sg13g2_buf_8
XFILLER_4_991 VPWR VGND sg13g2_decap_8
X_3263_ _0791_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] net663 VPWR
+ VGND sg13g2_nand2_1
X_3194_ _0715_ _0717_ _0718_ _0720_ _0722_ VPWR VGND sg13g2_or4_1
X_2214_ _1571_ _1632_ _1634_ VPWR VGND sg13g2_nor2_1
X_2145_ net767 _1563_ _1565_ VPWR VGND sg13g2_nor2_2
XFILLER_38_144 VPWR VGND sg13g2_fill_2
XFILLER_39_656 VPWR VGND sg13g2_decap_8
XFILLER_26_328 VPWR VGND sg13g2_fill_1
X_2076_ VPWR _1498_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] VGND
+ sg13g2_inv_1
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_10_718 VPWR VGND sg13g2_decap_8
XFILLER_22_545 VPWR VGND sg13g2_decap_8
X_2978_ _0533_ _0530_ _0532_ VPWR VGND sg13g2_nand2_1
XFILLER_2_917 VPWR VGND sg13g2_decap_8
XFILLER_45_648 VPWR VGND sg13g2_decap_8
XFILLER_13_501 VPWR VGND sg13g2_decap_8
XFILLER_26_884 VPWR VGND sg13g2_decap_8
XFILLER_41_854 VPWR VGND sg13g2_decap_8
XFILLER_13_578 VPWR VGND sg13g2_decap_8
XFILLER_5_700 VPWR VGND sg13g2_decap_8
XFILLER_5_777 VPWR VGND sg13g2_decap_8
XFILLER_45_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_932 VPWR VGND sg13g2_decap_8
XFILLER_1_983 VPWR VGND sg13g2_decap_8
XFILLER_0_493 VPWR VGND sg13g2_decap_8
XFILLER_48_486 VPWR VGND sg13g2_decap_8
XFILLER_36_626 VPWR VGND sg13g2_decap_8
X_3950_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] _1309_
+ _1376_ net808 sg13g2_a21oi_1
XFILLER_17_851 VPWR VGND sg13g2_decap_8
XFILLER_35_169 VPWR VGND sg13g2_fill_1
X_2901_ _0458_ _0452_ _0457_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_832 VPWR VGND sg13g2_decap_8
X_3881_ _1303_ _1305_ _1314_ VPWR VGND sg13g2_nor2_2
XFILLER_31_331 VPWR VGND sg13g2_decap_4
X_2832_ _0391_ net625 _0388_ VPWR VGND sg13g2_nand2_1
X_2763_ _0324_ _0317_ _0318_ VPWR VGND sg13g2_nand2_2
X_2694_ net736 _0274_ _0276_ _0277_ VPWR VGND sg13g2_nor3_1
XFILLER_8_593 VPWR VGND sg13g2_decap_8
X_3315_ _0843_ _0710_ _0841_ VPWR VGND sg13g2_nand2_1
X_3246_ _0767_ _0768_ _0769_ _0770_ _0774_ VPWR VGND sg13g2_and4_1
X_3177_ _0705_ net688 _0694_ VPWR VGND sg13g2_nand2_2
X_2128_ net767 _1547_ _1548_ VPWR VGND sg13g2_nor2_2
XFILLER_27_637 VPWR VGND sg13g2_decap_8
XFILLER_42_618 VPWR VGND sg13g2_decap_8
X_2059_ VPWR _1481_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] VGND
+ sg13g2_inv_1
XFILLER_25_48 VPWR VGND sg13g2_fill_2
XFILLER_23_876 VPWR VGND sg13g2_decap_8
XFILLER_10_515 VPWR VGND sg13g2_decap_8
XFILLER_2_714 VPWR VGND sg13g2_decap_8
XFILLER_1_235 VPWR VGND sg13g2_fill_2
XFILLER_46_968 VPWR VGND sg13g2_decap_8
XFILLER_45_445 VPWR VGND sg13g2_decap_8
XFILLER_18_637 VPWR VGND sg13g2_decap_8
XFILLER_14_821 VPWR VGND sg13g2_decap_8
XFILLER_26_681 VPWR VGND sg13g2_decap_8
XFILLER_41_651 VPWR VGND sg13g2_decap_8
XFILLER_14_898 VPWR VGND sg13g2_decap_8
XFILLER_12_1015 VPWR VGND sg13g2_decap_8
XFILLER_5_574 VPWR VGND sg13g2_decap_8
X_3100_ _0628_ _1638_ net753 VPWR VGND sg13g2_nand2b_1
XFILLER_1_780 VPWR VGND sg13g2_decap_8
X_4080_ net831 VGND VPWR _0044_ sap_3_inst.out\[3\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3031_ _0427_ _0451_ _0511_ _0549_ _0576_ VPWR VGND sg13g2_nor4_1
XFILLER_48_283 VPWR VGND sg13g2_decap_8
XFILLER_37_968 VPWR VGND sg13g2_decap_8
XFILLER_24_629 VPWR VGND sg13g2_decap_8
X_3933_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] _1314_
+ _1361_ net807 sg13g2_a21oi_1
X_3864_ VGND VPWR _0155_ _1297_ _0160_ _1287_ sg13g2_a21oi_1
X_2815_ _0369_ VPWR _0375_ VGND net804 _0324_ sg13g2_o21ai_1
XFILLER_20_857 VPWR VGND sg13g2_decap_8
X_3795_ net614 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] _1250_ _0138_
+ VPWR VGND sg13g2_a21o_1
X_2746_ _1713_ VPWR _0307_ VGND _0301_ _0306_ sg13g2_o21ai_1
X_2677_ VGND VPWR _1822_ _0260_ mem_ram_we _1531_ sg13g2_a21oi_1
XFILLER_28_1022 VPWR VGND sg13g2_decap_8
X_3229_ net703 net697 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] _0757_
+ VPWR VGND net692 sg13g2_nand4_1
XFILLER_28_924 VPWR VGND sg13g2_decap_8
XFILLER_27_412 VPWR VGND sg13g2_fill_2
XFILLER_27_434 VPWR VGND sg13g2_decap_8
XFILLER_43_938 VPWR VGND sg13g2_decap_8
XFILLER_42_415 VPWR VGND sg13g2_decap_8
XFILLER_36_990 VPWR VGND sg13g2_decap_8
XFILLER_35_1004 VPWR VGND sg13g2_decap_8
XFILLER_23_673 VPWR VGND sg13g2_decap_8
XFILLER_11_846 VPWR VGND sg13g2_decap_8
XFILLER_7_817 VPWR VGND sg13g2_decap_8
Xclkbuf_4_8_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_8_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_2_511 VPWR VGND sg13g2_decap_8
XFILLER_7_2 VPWR VGND sg13g2_fill_1
XFILLER_2_588 VPWR VGND sg13g2_decap_8
XFILLER_19_913 VPWR VGND sg13g2_decap_8
XFILLER_46_765 VPWR VGND sg13g2_decap_8
XFILLER_34_927 VPWR VGND sg13g2_decap_8
XFILLER_42_982 VPWR VGND sg13g2_decap_8
XFILLER_14_695 VPWR VGND sg13g2_decap_8
X_2600_ _2009_ net789 net792 VPWR VGND sg13g2_xnor2_1
X_3580_ _0083_ _1085_ _1090_ net618 _1466_ VPWR VGND sg13g2_a22oi_1
X_2531_ _1942_ VPWR _1943_ VGND net737 _1938_ sg13g2_o21ai_1
XFILLER_6_894 VPWR VGND sg13g2_decap_8
X_2462_ _1880_ net628 _1879_ VPWR VGND sg13g2_nand2_1
X_4201_ net846 VGND VPWR _0165_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[4\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_1
X_2393_ _1813_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] net647
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4132_ net826 VGND VPWR _0096_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_3_1002 VPWR VGND sg13g2_decap_8
XFILLER_3_95 VPWR VGND sg13g2_fill_2
X_4063_ net821 VGND VPWR _0003_ sap_3_inst.controller.stage\[2\] net44 sg13g2_dfrbpq_1
X_3014_ _0567_ VPWR _0568_ VGND _0565_ _0566_ sg13g2_o21ai_1
XFILLER_37_765 VPWR VGND sg13g2_decap_8
XFILLER_24_426 VPWR VGND sg13g2_decap_8
XFILLER_40_919 VPWR VGND sg13g2_decap_8
Xclkbuf_5_7__f_sap_3_inst.alu.clk_regs clknet_4_3_0_sap_3_inst.alu.clk_regs clknet_5_7__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3916_ _1346_ net809 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] _1307_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_654 VPWR VGND sg13g2_decap_8
X_3847_ VGND VPWR net817 _0155_ _1284_ net56 sg13g2_a21oi_1
X_3778_ _1236_ _1237_ _1238_ VPWR VGND sg13g2_nor2_1
XFILLER_4_809 VPWR VGND sg13g2_decap_8
X_2729_ VPWR mem_mar_we _0299_ VGND sg13g2_inv_1
XFILLER_47_529 VPWR VGND sg13g2_decap_8
XFILLER_28_721 VPWR VGND sg13g2_decap_8
XFILLER_27_220 VPWR VGND sg13g2_fill_2
XFILLER_43_735 VPWR VGND sg13g2_decap_8
XFILLER_16_927 VPWR VGND sg13g2_decap_8
XFILLER_28_798 VPWR VGND sg13g2_decap_8
XFILLER_23_470 VPWR VGND sg13g2_decap_8
XFILLER_24_993 VPWR VGND sg13g2_decap_8
XFILLER_7_614 VPWR VGND sg13g2_decap_8
XFILLER_11_643 VPWR VGND sg13g2_decap_8
XFILLER_3_820 VPWR VGND sg13g2_decap_8
XFILLER_3_897 VPWR VGND sg13g2_decap_8
XFILLER_19_710 VPWR VGND sg13g2_decap_8
XFILLER_46_562 VPWR VGND sg13g2_decap_8
XFILLER_19_787 VPWR VGND sg13g2_decap_8
XFILLER_34_724 VPWR VGND sg13g2_decap_8
Xclkbuf_5_14__f_sap_3_inst.alu.clk_regs clknet_4_7_0_sap_3_inst.alu.clk_regs clknet_5_14__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3701_ _1185_ VPWR _1186_ VGND net713 _1184_ sg13g2_o21ai_1
X_3632_ _1131_ _1061_ _1062_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_996 VPWR VGND sg13g2_decap_8
X_3563_ net618 net684 _1075_ VPWR VGND sg13g2_nor2_2
XFILLER_45_0 VPWR VGND sg13g2_fill_1
X_3494_ net602 VPWR _1016_ VGND net669 _1015_ sg13g2_o21ai_1
XFILLER_6_691 VPWR VGND sg13g2_decap_8
X_2514_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] net642
+ net633 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] _1928_ net722 sg13g2_a221oi_1
X_2445_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] _1864_
+ _1811_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] _1865_ _1806_ sg13g2_a221oi_1
X_4115_ net828 VGND VPWR _0079_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\]
+ clknet_5_13__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2376_ _1503_ _1557_ net786 _1796_ VPWR VGND _1676_ sg13g2_nand4_1
XFILLER_37_562 VPWR VGND sg13g2_decap_8
XFILLER_25_757 VPWR VGND sg13g2_decap_8
XFILLER_40_716 VPWR VGND sg13g2_decap_8
XFILLER_33_59 VPWR VGND sg13g2_fill_2
X_4043__8 VPWR net44 clknet_leaf_2_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_21_963 VPWR VGND sg13g2_decap_8
XFILLER_32_1007 VPWR VGND sg13g2_decap_8
XFILLER_4_606 VPWR VGND sg13g2_decap_8
XFILLER_0_801 VPWR VGND sg13g2_decap_8
XFILLER_47_304 VPWR VGND sg13g2_fill_2
XFILLER_0_878 VPWR VGND sg13g2_decap_8
XFILLER_47_326 VPWR VGND sg13g2_decap_8
XFILLER_16_724 VPWR VGND sg13g2_decap_8
XFILLER_43_532 VPWR VGND sg13g2_decap_8
XFILLER_28_595 VPWR VGND sg13g2_decap_8
XFILLER_24_790 VPWR VGND sg13g2_decap_8
XFILLER_31_738 VPWR VGND sg13g2_decap_8
XFILLER_8_901 VPWR VGND sg13g2_decap_8
XFILLER_12_952 VPWR VGND sg13g2_decap_8
XFILLER_8_978 VPWR VGND sg13g2_decap_8
XFILLER_7_466 VPWR VGND sg13g2_fill_2
XFILLER_48_1025 VPWR VGND sg13g2_decap_4
XFILLER_3_694 VPWR VGND sg13g2_decap_8
X_2230_ _1644_ _1649_ _1650_ VPWR VGND sg13g2_nor2_1
XFILLER_2_160 VPWR VGND sg13g2_fill_2
X_2161_ net780 _1527_ _1563_ _1581_ VGND VPWR _1580_ sg13g2_nor4_2
XFILLER_17_4 VPWR VGND sg13g2_fill_1
XFILLER_39_838 VPWR VGND sg13g2_decap_8
X_2092_ _1512_ net782 VPWR VGND net785 sg13g2_nand2b_2
XFILLER_47_893 VPWR VGND sg13g2_decap_8
XFILLER_0_52 VPWR VGND sg13g2_decap_8
XFILLER_19_584 VPWR VGND sg13g2_decap_8
XFILLER_34_521 VPWR VGND sg13g2_decap_8
XFILLER_22_727 VPWR VGND sg13g2_decap_8
X_2994_ _0548_ net787 sap_3_inst.alu.tmp\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_34_598 VPWR VGND sg13g2_decap_8
XFILLER_30_793 VPWR VGND sg13g2_decap_8
X_3615_ VPWR VGND _1119_ net618 _1118_ net607 _1120_ _1030_ sg13g2_a221oi_1
X_3546_ VGND VPWR _0828_ _0987_ _1061_ net22 sg13g2_a21oi_1
X_3477_ _0999_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] net674 VPWR
+ VGND sg13g2_nand2_1
X_2428_ _1602_ _1685_ net777 _1848_ VPWR VGND sg13g2_nand3_1
X_2359_ VGND VPWR net783 _1720_ _1779_ _1520_ sg13g2_a21oi_1
XFILLER_29_304 VPWR VGND sg13g2_decap_8
X_4029_ VPWR _0191_ _1432_ VGND sg13g2_inv_1
XFILLER_44_36 VPWR VGND sg13g2_fill_1
XFILLER_25_554 VPWR VGND sg13g2_decap_8
XFILLER_40_513 VPWR VGND sg13g2_decap_8
XFILLER_21_760 VPWR VGND sg13g2_decap_8
XFILLER_5_959 VPWR VGND sg13g2_decap_8
XFILLER_0_675 VPWR VGND sg13g2_decap_8
XFILLER_48_668 VPWR VGND sg13g2_decap_8
XFILLER_36_808 VPWR VGND sg13g2_decap_8
XFILLER_29_860 VPWR VGND sg13g2_decap_8
XFILLER_44_841 VPWR VGND sg13g2_decap_8
XFILLER_16_521 VPWR VGND sg13g2_decap_8
XFILLER_16_598 VPWR VGND sg13g2_decap_8
XFILLER_31_535 VPWR VGND sg13g2_decap_8
XFILLER_8_775 VPWR VGND sg13g2_decap_8
X_3400_ _0923_ _0924_ _0925_ VPWR VGND sg13g2_and2_1
X_3331_ _0857_ _0858_ _0856_ _0859_ VPWR VGND sg13g2_nand3_1
XFILLER_4_970 VPWR VGND sg13g2_decap_8
XFILLER_3_491 VPWR VGND sg13g2_decap_8
X_3262_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] net697 net692 net687
+ _0790_ VPWR VGND sg13g2_and4_1
X_3193_ _0715_ _0717_ _0718_ _0721_ VGND VPWR _0720_ sg13g2_nor4_2
X_2213_ _1633_ net755 net747 VPWR VGND sg13g2_nand2_2
XFILLER_39_635 VPWR VGND sg13g2_decap_8
X_2144_ net780 net770 net768 _1564_ VPWR VGND sg13g2_nand3_1
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_819 VPWR VGND sg13g2_decap_8
XFILLER_47_690 VPWR VGND sg13g2_decap_8
X_2075_ VPWR _1497_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_35_885 VPWR VGND sg13g2_decap_8
XFILLER_22_524 VPWR VGND sg13g2_decap_8
X_2977_ _0531_ VPWR _0532_ VGND net793 net721 sg13g2_o21ai_1
XFILLER_30_590 VPWR VGND sg13g2_decap_8
X_3529_ net585 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] _1048_ _0074_
+ VPWR VGND sg13g2_a21o_1
XFILLER_29_101 VPWR VGND sg13g2_fill_2
XFILLER_45_627 VPWR VGND sg13g2_decap_8
XFILLER_18_819 VPWR VGND sg13g2_decap_8
XFILLER_26_863 VPWR VGND sg13g2_decap_8
XFILLER_41_833 VPWR VGND sg13g2_decap_8
XFILLER_38_1024 VPWR VGND sg13g2_decap_4
XFILLER_40_310 VPWR VGND sg13g2_fill_1
XFILLER_13_557 VPWR VGND sg13g2_decap_8
XFILLER_9_539 VPWR VGND sg13g2_decap_8
XFILLER_5_756 VPWR VGND sg13g2_decap_8
XFILLER_4_277 VPWR VGND sg13g2_fill_2
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_962 VPWR VGND sg13g2_decap_8
XFILLER_49_911 VPWR VGND sg13g2_decap_8
XFILLER_49_988 VPWR VGND sg13g2_decap_8
XFILLER_48_465 VPWR VGND sg13g2_decap_8
XFILLER_36_605 VPWR VGND sg13g2_decap_8
XFILLER_17_830 VPWR VGND sg13g2_decap_8
X_2900_ VGND VPWR _0418_ _0424_ _0457_ _0421_ sg13g2_a21oi_1
XFILLER_32_811 VPWR VGND sg13g2_decap_8
X_3880_ net816 net815 _1311_ _1313_ VPWR VGND sg13g2_a21o_1
X_2831_ _0388_ _0360_ _0390_ VPWR VGND sg13g2_xor2_1
XFILLER_32_888 VPWR VGND sg13g2_decap_8
X_2762_ sap_3_inst.alu.tmp\[0\] net806 _0323_ VPWR VGND sg13g2_xor2_1
XFILLER_8_572 VPWR VGND sg13g2_decap_8
X_2693_ _1935_ _0275_ _0276_ VPWR VGND sg13g2_nor2b_1
X_3314_ _0733_ _0742_ _0722_ _0842_ VPWR VGND _0837_ sg13g2_nand4_1
X_3245_ _0773_ net667 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] net671
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_421 VPWR VGND sg13g2_fill_1
XFILLER_27_616 VPWR VGND sg13g2_decap_8
X_3176_ _0704_ net701 net693 net688 VPWR VGND sg13g2_and3_1
XFILLER_39_454 VPWR VGND sg13g2_fill_1
X_2127_ _1547_ net769 net771 VPWR VGND sg13g2_nand2b_1
XFILLER_25_27 VPWR VGND sg13g2_fill_2
X_2058_ VPWR _1480_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[5\] VGND
+ sg13g2_inv_1
XFILLER_35_682 VPWR VGND sg13g2_decap_8
XFILLER_23_855 VPWR VGND sg13g2_decap_8
XFILLER_6_509 VPWR VGND sg13g2_decap_8
XFILLER_49_229 VPWR VGND sg13g2_decap_8
XFILLER_18_616 VPWR VGND sg13g2_decap_8
XFILLER_46_947 VPWR VGND sg13g2_decap_8
XFILLER_45_424 VPWR VGND sg13g2_decap_8
XFILLER_14_800 VPWR VGND sg13g2_decap_8
XFILLER_26_660 VPWR VGND sg13g2_decap_8
XFILLER_41_630 VPWR VGND sg13g2_decap_8
XFILLER_14_877 VPWR VGND sg13g2_decap_8
XFILLER_40_173 VPWR VGND sg13g2_fill_1
XFILLER_5_553 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_49_785 VPWR VGND sg13g2_decap_8
X_3030_ VGND VPWR _0548_ _0561_ _0575_ _0545_ sg13g2_a21oi_1
XFILLER_37_947 VPWR VGND sg13g2_decap_8
XFILLER_24_608 VPWR VGND sg13g2_decap_8
XFILLER_36_446 VPWR VGND sg13g2_fill_1
XFILLER_45_991 VPWR VGND sg13g2_decap_8
X_3932_ _1360_ _1308_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] net810
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_32_685 VPWR VGND sg13g2_decap_8
X_3863_ _1297_ _1296_ _1278_ _1281_ net54 VPWR VGND sg13g2_a22oi_1
X_2814_ VPWR VGND net625 _0362_ _0359_ _0335_ _0374_ _0356_ sg13g2_a221oi_1
XFILLER_20_836 VPWR VGND sg13g2_decap_8
X_3794_ net613 _1046_ _1047_ _1250_ VPWR VGND sg13g2_nor3_1
X_2745_ VGND VPWR _1685_ _0302_ _0306_ _0305_ sg13g2_a21oi_1
X_2676_ _1834_ VPWR _0260_ VGND _1731_ _0259_ sg13g2_o21ai_1
XFILLER_28_1001 VPWR VGND sg13g2_decap_8
XFILLER_28_903 VPWR VGND sg13g2_decap_8
X_3228_ _0748_ _0752_ _0753_ _0754_ _0756_ VPWR VGND sg13g2_or4_1
X_3159_ _0686_ _0685_ _0684_ _0687_ VPWR VGND sg13g2_a21o_2
XFILLER_39_273 VPWR VGND sg13g2_fill_1
XFILLER_43_917 VPWR VGND sg13g2_decap_8
XFILLER_11_825 VPWR VGND sg13g2_decap_8
XFILLER_23_652 VPWR VGND sg13g2_decap_8
XFILLER_6_328 VPWR VGND sg13g2_fill_2
XFILLER_2_567 VPWR VGND sg13g2_decap_8
XFILLER_46_744 VPWR VGND sg13g2_decap_8
XFILLER_19_969 VPWR VGND sg13g2_decap_8
XFILLER_34_906 VPWR VGND sg13g2_decap_8
XFILLER_27_980 VPWR VGND sg13g2_decap_8
XFILLER_42_961 VPWR VGND sg13g2_decap_8
XFILLER_14_674 VPWR VGND sg13g2_decap_8
X_2530_ _1942_ _1548_ net735 VPWR VGND sg13g2_nand2_1
XFILLER_6_873 VPWR VGND sg13g2_decap_8
X_2461_ _1879_ sap_3_inst.alu.flags\[6\] _1839_ VPWR VGND sg13g2_nand2_1
X_4200_ net841 VGND VPWR _0164_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[3\]
+ clknet_3_3__leaf_clk sg13g2_dfrbpq_1
X_2392_ _1738_ _1765_ _1783_ _1812_ VGND VPWR _1799_ sg13g2_nor4_2
X_4131_ net828 VGND VPWR _0095_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\]
+ clknet_5_13__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_3_41 VPWR VGND sg13g2_fill_2
X_4062_ net821 VGND VPWR _0002_ sap_3_inst.controller.stage\[1\] net43 sg13g2_dfrbpq_2
XFILLER_49_582 VPWR VGND sg13g2_decap_8
X_3013_ VGND VPWR sap_3_inst.alu.act\[7\] _0314_ _0567_ net627 sg13g2_a21oi_1
XFILLER_37_744 VPWR VGND sg13g2_decap_8
XFILLER_18_980 VPWR VGND sg13g2_decap_8
XFILLER_24_405 VPWR VGND sg13g2_decap_8
XFILLER_25_939 VPWR VGND sg13g2_decap_8
XFILLER_36_287 VPWR VGND sg13g2_decap_4
X_3915_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] _1306_
+ _1345_ net807 sg13g2_a21oi_1
XFILLER_20_633 VPWR VGND sg13g2_decap_8
XFILLER_33_994 VPWR VGND sg13g2_decap_8
X_3846_ VGND VPWR net817 _0155_ _0156_ _1283_ sg13g2_a21oi_1
X_3777_ _1237_ _0872_ _0955_ VPWR VGND sg13g2_nand2_1
X_2728_ _0299_ _1538_ _0298_ _1505_ net758 VPWR VGND sg13g2_a22oi_1
X_2659_ _0246_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] net722
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_47_508 VPWR VGND sg13g2_decap_8
XFILLER_28_700 VPWR VGND sg13g2_decap_8
XFILLER_16_906 VPWR VGND sg13g2_decap_8
XFILLER_28_777 VPWR VGND sg13g2_decap_8
XFILLER_43_714 VPWR VGND sg13g2_decap_8
XFILLER_24_972 VPWR VGND sg13g2_decap_8
XFILLER_11_622 VPWR VGND sg13g2_decap_8
XFILLER_11_699 VPWR VGND sg13g2_decap_8
XFILLER_6_136 VPWR VGND sg13g2_fill_1
XFILLER_3_876 VPWR VGND sg13g2_decap_8
Xfanout690 _0659_ net690 VPWR VGND sg13g2_buf_8
XFILLER_46_541 VPWR VGND sg13g2_decap_8
XFILLER_19_766 VPWR VGND sg13g2_decap_8
XFILLER_34_703 VPWR VGND sg13g2_decap_8
XFILLER_22_909 VPWR VGND sg13g2_decap_8
XFILLER_18_1022 VPWR VGND sg13g2_decap_8
XFILLER_33_268 VPWR VGND sg13g2_fill_1
XFILLER_15_994 VPWR VGND sg13g2_decap_8
X_3700_ _1185_ _0946_ net604 net597 net572 VPWR VGND sg13g2_a22oi_1
XFILLER_30_975 VPWR VGND sg13g2_decap_8
X_3631_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] _1060_ _1122_ _0094_
+ VPWR VGND sg13g2_mux2_1
X_3562_ _1074_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] net620 VPWR
+ VGND sg13g2_nand2_1
XFILLER_6_670 VPWR VGND sg13g2_decap_8
X_2513_ _1927_ _1925_ _1926_ VPWR VGND sg13g2_nand2_1
X_3493_ _1015_ _0732_ _0845_ VPWR VGND sg13g2_xnor2_1
X_2444_ _1861_ _1862_ _1860_ _1864_ VPWR VGND _1863_ sg13g2_nand4_1
X_2375_ _1789_ _1794_ _1785_ _1795_ VPWR VGND sg13g2_nand3_1
X_4114_ net841 VGND VPWR _0078_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\]
+ clknet_5_31__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_37_541 VPWR VGND sg13g2_decap_8
XFILLER_25_736 VPWR VGND sg13g2_decap_8
XFILLER_33_791 VPWR VGND sg13g2_decap_8
XFILLER_21_942 VPWR VGND sg13g2_decap_8
X_3829_ net15 net610 _1114_ _1271_ VPWR VGND sg13g2_nor3_1
XFILLER_0_857 VPWR VGND sg13g2_decap_8
XFILLER_43_511 VPWR VGND sg13g2_decap_8
XFILLER_16_703 VPWR VGND sg13g2_decap_8
XFILLER_28_574 VPWR VGND sg13g2_decap_8
XFILLER_31_717 VPWR VGND sg13g2_decap_8
XFILLER_43_588 VPWR VGND sg13g2_decap_8
XFILLER_12_931 VPWR VGND sg13g2_decap_8
XFILLER_8_957 VPWR VGND sg13g2_decap_8
XFILLER_11_496 VPWR VGND sg13g2_decap_8
XFILLER_48_1004 VPWR VGND sg13g2_decap_8
XFILLER_3_673 VPWR VGND sg13g2_decap_8
XFILLER_39_817 VPWR VGND sg13g2_decap_8
X_2160_ net785 net779 _1580_ VPWR VGND net782 sg13g2_nand3b_1
X_2091_ sap_3_inst.controller.opcode\[0\] net784 _1511_ VPWR VGND sg13g2_nor2b_2
XFILLER_47_872 VPWR VGND sg13g2_decap_8
XFILLER_0_31 VPWR VGND sg13g2_decap_8
XFILLER_19_563 VPWR VGND sg13g2_decap_8
XFILLER_34_500 VPWR VGND sg13g2_decap_8
XFILLER_22_706 VPWR VGND sg13g2_decap_8
XFILLER_34_577 VPWR VGND sg13g2_decap_8
X_2993_ net787 sap_3_inst.alu.tmp\[7\] _0547_ VPWR VGND sg13g2_and2_1
XFILLER_15_791 VPWR VGND sg13g2_decap_8
XFILLER_14_290 VPWR VGND sg13g2_fill_1
XFILLER_30_772 VPWR VGND sg13g2_decap_8
X_3614_ _1119_ _0289_ _1075_ VPWR VGND sg13g2_nand2_1
X_3545_ _1060_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] net585 _0078_
+ VPWR VGND sg13g2_mux2_1
XFILLER_0_109 VPWR VGND sg13g2_fill_1
X_3476_ _0970_ VPWR _0071_ VGND _0986_ _0998_ sg13g2_o21ai_1
X_2427_ net752 _1846_ _1847_ VPWR VGND sg13g2_and2_1
X_2358_ _1777_ VPWR _1778_ VGND _1773_ _1776_ sg13g2_o21ai_1
XFILLER_45_809 VPWR VGND sg13g2_decap_8
X_2289_ _1641_ _1708_ _1709_ VPWR VGND sg13g2_and2_1
X_4028_ _1432_ _1430_ net816 _1429_ net809 VPWR VGND sg13g2_a22oi_1
XFILLER_25_533 VPWR VGND sg13g2_decap_8
XFILLER_13_739 VPWR VGND sg13g2_decap_8
XFILLER_40_569 VPWR VGND sg13g2_decap_8
XFILLER_5_938 VPWR VGND sg13g2_decap_8
XFILLER_0_654 VPWR VGND sg13g2_decap_8
XFILLER_48_647 VPWR VGND sg13g2_decap_8
XFILLER_16_500 VPWR VGND sg13g2_decap_8
XFILLER_44_820 VPWR VGND sg13g2_decap_8
XFILLER_44_897 VPWR VGND sg13g2_decap_8
XFILLER_43_385 VPWR VGND sg13g2_decap_8
XFILLER_16_577 VPWR VGND sg13g2_decap_8
XFILLER_31_514 VPWR VGND sg13g2_decap_8
XFILLER_8_754 VPWR VGND sg13g2_decap_8
X_3330_ _1769_ _0625_ _0854_ _0855_ _0858_ VPWR VGND sg13g2_nor4_1
X_3261_ _0777_ _0785_ _0786_ _0787_ _0789_ VPWR VGND sg13g2_or4_1
X_3192_ _0720_ _0716_ _0719_ VPWR VGND sg13g2_nand2_1
X_2212_ net755 net746 _1632_ VPWR VGND sg13g2_and2_1
XFILLER_22_1007 VPWR VGND sg13g2_decap_8
XFILLER_39_614 VPWR VGND sg13g2_decap_8
X_2143_ _1563_ net768 net770 VPWR VGND sg13g2_nand2_2
X_2074_ VPWR _1496_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_35_864 VPWR VGND sg13g2_decap_8
XFILLER_22_503 VPWR VGND sg13g2_decap_8
X_2976_ _0531_ _0477_ _0478_ VPWR VGND sg13g2_nand2_1
XFILLER_30_39 VPWR VGND sg13g2_fill_1
X_3528_ net585 _1046_ _1047_ _1048_ VPWR VGND sg13g2_nor3_1
X_3459_ net602 VPWR _0982_ VGND net669 _0981_ sg13g2_o21ai_1
XFILLER_45_606 VPWR VGND sg13g2_decap_8
XFILLER_26_842 VPWR VGND sg13g2_decap_8
XFILLER_38_1003 VPWR VGND sg13g2_decap_8
XFILLER_41_812 VPWR VGND sg13g2_decap_8
XFILLER_13_536 VPWR VGND sg13g2_decap_8
XFILLER_41_889 VPWR VGND sg13g2_decap_8
XFILLER_9_518 VPWR VGND sg13g2_decap_8
XFILLER_5_735 VPWR VGND sg13g2_decap_8
XFILLER_1_941 VPWR VGND sg13g2_decap_8
XFILLER_49_967 VPWR VGND sg13g2_decap_8
XFILLER_48_444 VPWR VGND sg13g2_decap_8
XFILLER_44_694 VPWR VGND sg13g2_decap_8
XFILLER_17_886 VPWR VGND sg13g2_decap_8
X_2830_ _0389_ _0360_ _0388_ VPWR VGND sg13g2_nand2b_1
XFILLER_32_867 VPWR VGND sg13g2_decap_8
X_2761_ _0322_ net806 sap_3_inst.alu.tmp\[0\] VPWR VGND sg13g2_nand2_1
X_2692_ VPWR VGND _1685_ _1787_ _1566_ net735 _0275_ _1565_ sg13g2_a221oi_1
XFILLER_8_551 VPWR VGND sg13g2_decap_8
X_3313_ _0721_ _0732_ _0741_ _0838_ _0841_ VPWR VGND sg13g2_nor4_1
X_3244_ _0772_ net666 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] net674
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_0 VPWR VGND sg13g2_fill_1
X_3175_ _0703_ _0662_ net688 VPWR VGND sg13g2_nand2_1
X_2126_ _1443_ net771 _1546_ VPWR VGND sg13g2_nor2_1
XFILLER_39_488 VPWR VGND sg13g2_decap_8
X_2057_ VPWR _1479_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_23_834 VPWR VGND sg13g2_decap_8
XFILLER_35_661 VPWR VGND sg13g2_decap_8
X_2959_ _0513_ VPWR _0514_ VGND _0495_ _0512_ sg13g2_o21ai_1
XFILLER_2_749 VPWR VGND sg13g2_decap_8
XFILLER_46_926 VPWR VGND sg13g2_decap_8
XFILLER_45_403 VPWR VGND sg13g2_decap_8
XFILLER_33_609 VPWR VGND sg13g2_decap_8
XFILLER_14_856 VPWR VGND sg13g2_decap_8
XFILLER_41_686 VPWR VGND sg13g2_decap_8
XFILLER_5_532 VPWR VGND sg13g2_decap_8
XFILLER_49_764 VPWR VGND sg13g2_decap_8
XFILLER_37_926 VPWR VGND sg13g2_decap_8
XFILLER_36_436 VPWR VGND sg13g2_fill_1
XFILLER_45_970 VPWR VGND sg13g2_decap_8
XFILLER_17_683 VPWR VGND sg13g2_decap_8
XFILLER_44_491 VPWR VGND sg13g2_decap_8
X_3931_ _1359_ net809 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] _1307_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_815 VPWR VGND sg13g2_decap_8
X_3862_ VGND VPWR _1289_ _1291_ _1296_ _1295_ sg13g2_a21oi_1
XFILLER_32_664 VPWR VGND sg13g2_decap_8
X_2813_ _0370_ _0372_ _0329_ _0373_ VPWR VGND sg13g2_nand3_1
X_3793_ _1245_ VPWR _0137_ VGND _1248_ _1249_ sg13g2_o21ai_1
X_2744_ _1848_ _0303_ _1843_ _0305_ VPWR VGND _0304_ sg13g2_nand4_1
XFILLER_9_882 VPWR VGND sg13g2_decap_8
X_2675_ _1706_ _1752_ _1700_ _0259_ VPWR VGND _1826_ sg13g2_nand4_1
X_3227_ _0748_ _0752_ _0753_ _0755_ VGND VPWR _0754_ sg13g2_nor4_2
XFILLER_39_241 VPWR VGND sg13g2_fill_1
X_3158_ _0686_ net764 _1535_ VPWR VGND sg13g2_nand2_1
XFILLER_27_414 VPWR VGND sg13g2_fill_1
XFILLER_28_959 VPWR VGND sg13g2_decap_8
X_2109_ _1525_ _1526_ _1523_ _1529_ VPWR VGND _1528_ sg13g2_nand4_1
XFILLER_15_609 VPWR VGND sg13g2_decap_8
XFILLER_27_469 VPWR VGND sg13g2_decap_8
X_3089_ _0616_ VPWR _0617_ VGND net724 _0614_ sg13g2_o21ai_1
XFILLER_23_631 VPWR VGND sg13g2_decap_8
XFILLER_11_804 VPWR VGND sg13g2_decap_8
XFILLER_2_546 VPWR VGND sg13g2_decap_8
Xclkbuf_5_22__f_sap_3_inst.alu.clk_regs clknet_4_11_0_sap_3_inst.alu.clk_regs clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_46_723 VPWR VGND sg13g2_decap_8
XFILLER_19_948 VPWR VGND sg13g2_decap_8
XFILLER_42_940 VPWR VGND sg13g2_decap_8
XFILLER_14_653 VPWR VGND sg13g2_decap_8
XFILLER_41_483 VPWR VGND sg13g2_decap_8
XFILLER_6_852 VPWR VGND sg13g2_decap_8
X_2460_ VGND VPWR _1878_ net629 net792 sg13g2_or2_1
XFILLER_5_395 VPWR VGND sg13g2_fill_1
X_2391_ _1738_ _1765_ _1784_ _1811_ VGND VPWR _1798_ sg13g2_nor4_2
X_4130_ net841 VGND VPWR _0094_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\]
+ clknet_5_31__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_3_64 VPWR VGND sg13g2_decap_8
XFILLER_49_561 VPWR VGND sg13g2_decap_8
X_4061_ net821 VGND VPWR _0001_ sap_3_inst.controller.stage\[0\] net42 sg13g2_dfrbpq_1
X_3012_ _0562_ net575 net707 _0566_ VPWR VGND sg13g2_a21o_1
XFILLER_37_723 VPWR VGND sg13g2_decap_8
XFILLER_25_918 VPWR VGND sg13g2_decap_8
XFILLER_36_277 VPWR VGND sg13g2_fill_2
X_3914_ _1344_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] _1309_
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_973 VPWR VGND sg13g2_decap_8
XFILLER_20_612 VPWR VGND sg13g2_decap_8
X_3845_ net817 _1278_ _1283_ VPWR VGND sg13g2_nor2_1
XFILLER_20_689 VPWR VGND sg13g2_decap_8
X_3776_ VGND VPWR _0908_ _0930_ _1236_ _0953_ sg13g2_a21oi_1
X_2727_ _0298_ net757 _0297_ VPWR VGND sg13g2_nand2_1
X_2658_ _0245_ net637 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] net640
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2589_ _1999_ _1996_ _1998_ _1858_ net3 VPWR VGND sg13g2_a22oi_1
XFILLER_28_756 VPWR VGND sg13g2_decap_8
XFILLER_24_951 VPWR VGND sg13g2_decap_8
XFILLER_10_100 VPWR VGND sg13g2_fill_2
XFILLER_11_601 VPWR VGND sg13g2_decap_8
XFILLER_10_122 VPWR VGND sg13g2_fill_1
XFILLER_7_649 VPWR VGND sg13g2_decap_8
XFILLER_11_678 VPWR VGND sg13g2_decap_8
XFILLER_3_855 VPWR VGND sg13g2_decap_8
Xfanout691 _0658_ net691 VPWR VGND sg13g2_buf_8
Xfanout680 _0660_ net680 VPWR VGND sg13g2_buf_8
XFILLER_46_520 VPWR VGND sg13g2_decap_8
XFILLER_18_233 VPWR VGND sg13g2_fill_2
XFILLER_19_745 VPWR VGND sg13g2_decap_8
XFILLER_46_597 VPWR VGND sg13g2_decap_8
XFILLER_34_759 VPWR VGND sg13g2_decap_8
XFILLER_15_973 VPWR VGND sg13g2_decap_8
XFILLER_18_1001 VPWR VGND sg13g2_decap_8
XFILLER_30_954 VPWR VGND sg13g2_decap_8
X_3630_ VGND VPWR _1451_ _1121_ _0093_ _1130_ sg13g2_a21oi_1
X_3561_ VGND VPWR _1501_ net585 _0081_ _1073_ sg13g2_a21oi_1
X_2512_ _1926_ net638 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] net646
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3492_ VGND VPWR _1013_ _1014_ _1007_ _0979_ sg13g2_a21oi_2
X_2443_ _1863_ _1807_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] net650
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2374_ _1682_ net723 _1791_ _1793_ _1794_ VPWR VGND sg13g2_nor4_1
XFILLER_25_1016 VPWR VGND sg13g2_decap_8
X_4113_ net822 VGND VPWR _0077_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\]
+ clknet_5_6__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_25_1027 VPWR VGND sg13g2_fill_2
XFILLER_37_520 VPWR VGND sg13g2_decap_8
XFILLER_25_715 VPWR VGND sg13g2_decap_8
XFILLER_37_597 VPWR VGND sg13g2_decap_8
XFILLER_21_921 VPWR VGND sg13g2_decap_8
XFILLER_33_770 VPWR VGND sg13g2_decap_8
XFILLER_21_998 VPWR VGND sg13g2_decap_8
X_3828_ _0151_ _1270_ _0288_ net610 _1481_ VPWR VGND sg13g2_a22oi_1
X_3759_ _1222_ _1221_ _0896_ _1219_ _0893_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_836 VPWR VGND sg13g2_decap_8
XFILLER_48_829 VPWR VGND sg13g2_decap_8
XFILLER_47_306 VPWR VGND sg13g2_fill_1
XFILLER_28_553 VPWR VGND sg13g2_decap_8
XFILLER_16_759 VPWR VGND sg13g2_decap_8
XFILLER_43_567 VPWR VGND sg13g2_decap_8
XFILLER_12_910 VPWR VGND sg13g2_decap_8
XFILLER_8_936 VPWR VGND sg13g2_decap_8
XFILLER_12_987 VPWR VGND sg13g2_decap_8
Xclkbuf_4_1_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_1_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_3_652 VPWR VGND sg13g2_decap_8
XFILLER_2_162 VPWR VGND sg13g2_fill_1
Xclkbuf_5_19__f_sap_3_inst.alu.clk_regs clknet_4_9_0_sap_3_inst.alu.clk_regs clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_47_851 VPWR VGND sg13g2_decap_8
X_2090_ _1510_ _1505_ _1507_ VPWR VGND sg13g2_nand2_1
XFILLER_19_542 VPWR VGND sg13g2_decap_8
XFILLER_0_1018 VPWR VGND sg13g2_decap_8
XFILLER_46_394 VPWR VGND sg13g2_decap_8
XFILLER_0_87 VPWR VGND sg13g2_fill_2
X_4047__12 VPWR net48 clknet_leaf_0_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_34_556 VPWR VGND sg13g2_decap_8
X_2992_ VGND VPWR _0546_ sap_3_inst.alu.tmp\[7\] net787 sg13g2_or2_1
XFILLER_15_770 VPWR VGND sg13g2_decap_8
XFILLER_9_41 VPWR VGND sg13g2_fill_2
XFILLER_30_751 VPWR VGND sg13g2_decap_8
X_3613_ _1118_ _1076_ net34 VPWR VGND sg13g2_nand2b_1
X_3544_ _1057_ _1059_ _1060_ VPWR VGND sg13g2_nor2_2
X_3475_ VGND VPWR net669 _0995_ _0998_ _0997_ sg13g2_a21oi_1
X_2426_ net731 VPWR _1846_ VGND _1441_ _1648_ sg13g2_o21ai_1
X_2357_ _1555_ net725 _1777_ VPWR VGND sg13g2_nor2_1
X_2288_ _1635_ _1696_ _1699_ _1707_ _1708_ VPWR VGND sg13g2_nor4_1
X_4027_ _1430_ _1431_ _0190_ VPWR VGND sg13g2_and2_1
XFILLER_38_884 VPWR VGND sg13g2_decap_8
XFILLER_25_512 VPWR VGND sg13g2_decap_8
XFILLER_13_718 VPWR VGND sg13g2_decap_8
XFILLER_25_589 VPWR VGND sg13g2_decap_8
XFILLER_40_548 VPWR VGND sg13g2_decap_8
XFILLER_21_795 VPWR VGND sg13g2_decap_8
XFILLER_5_917 VPWR VGND sg13g2_decap_8
XFILLER_0_633 VPWR VGND sg13g2_decap_8
XFILLER_48_626 VPWR VGND sg13g2_decap_8
XFILLER_18_83 VPWR VGND sg13g2_fill_1
XFILLER_29_895 VPWR VGND sg13g2_decap_8
XFILLER_44_876 VPWR VGND sg13g2_decap_8
XFILLER_16_556 VPWR VGND sg13g2_decap_8
XFILLER_34_71 VPWR VGND sg13g2_fill_2
XFILLER_15_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_733 VPWR VGND sg13g2_decap_8
XFILLER_12_784 VPWR VGND sg13g2_decap_8
X_3260_ _0777_ _0785_ _0786_ _0787_ _0788_ VPWR VGND sg13g2_nor4_1
X_3191_ _0719_ net658 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] net680
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2211_ net759 sap_3_inst.controller.stage\[3\] _1631_ VPWR VGND sg13g2_nor2b_1
X_2142_ net768 net770 _1562_ VPWR VGND sg13g2_and2_1
X_2073_ VPWR _1495_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_35_843 VPWR VGND sg13g2_decap_8
XFILLER_22_559 VPWR VGND sg13g2_decap_8
X_2975_ _0530_ net790 net721 VPWR VGND sg13g2_xnor2_1
X_3527_ net592 net598 _1047_ VPWR VGND sg13g2_nor2_2
XFILLER_1_408 VPWR VGND sg13g2_fill_2
X_3458_ _0981_ _0741_ _0844_ VPWR VGND sg13g2_xnor2_1
X_2409_ net763 _1560_ _1575_ _1829_ VPWR VGND sg13g2_nor3_1
X_3389_ _0915_ net19 net595 VPWR VGND sg13g2_nand2_1
XFILLER_26_821 VPWR VGND sg13g2_decap_8
XFILLER_38_681 VPWR VGND sg13g2_decap_8
XFILLER_13_515 VPWR VGND sg13g2_decap_8
XFILLER_26_898 VPWR VGND sg13g2_decap_8
XFILLER_41_868 VPWR VGND sg13g2_decap_8
XFILLER_25_386 VPWR VGND sg13g2_decap_8
XFILLER_21_592 VPWR VGND sg13g2_decap_8
XFILLER_5_714 VPWR VGND sg13g2_decap_8
XFILLER_1_920 VPWR VGND sg13g2_decap_8
XFILLER_45_1019 VPWR VGND sg13g2_decap_8
XFILLER_1_997 VPWR VGND sg13g2_decap_8
XFILLER_49_946 VPWR VGND sg13g2_decap_8
XFILLER_48_423 VPWR VGND sg13g2_decap_8
XFILLER_29_692 VPWR VGND sg13g2_decap_8
XFILLER_17_865 VPWR VGND sg13g2_decap_8
XFILLER_44_673 VPWR VGND sg13g2_decap_8
XFILLER_43_150 VPWR VGND sg13g2_fill_1
XFILLER_32_846 VPWR VGND sg13g2_decap_8
XFILLER_8_530 VPWR VGND sg13g2_decap_8
X_2760_ _0320_ VPWR _0321_ VGND net626 _0315_ sg13g2_o21ai_1
XFILLER_12_581 VPWR VGND sg13g2_decap_8
X_2691_ VGND VPWR _1630_ _0264_ _0274_ _0273_ sg13g2_a21oi_1
X_3312_ _0742_ _0837_ _0733_ _0840_ VPWR VGND sg13g2_nand3_1
X_3243_ _0771_ net663 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] net676
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_1013 VPWR VGND sg13g2_decap_8
X_3174_ _0702_ net700 net693 net688 VPWR VGND sg13g2_and3_2
XFILLER_39_467 VPWR VGND sg13g2_decap_8
XFILLER_48_990 VPWR VGND sg13g2_decap_8
X_2125_ _1443_ net766 _1545_ VPWR VGND sg13g2_nor2_1
XFILLER_26_117 VPWR VGND sg13g2_decap_4
X_2056_ VPWR _1478_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_35_640 VPWR VGND sg13g2_decap_8
XFILLER_23_813 VPWR VGND sg13g2_decap_8
XFILLER_10_529 VPWR VGND sg13g2_decap_8
X_2958_ _0513_ net794 sap_3_inst.alu.tmp\[5\] VPWR VGND sg13g2_nand2b_1
X_2889_ VPWR _0446_ _0445_ VGND sg13g2_inv_1
XFILLER_2_728 VPWR VGND sg13g2_decap_8
XFILLER_46_905 VPWR VGND sg13g2_decap_8
XFILLER_45_459 VPWR VGND sg13g2_decap_8
XFILLER_14_835 VPWR VGND sg13g2_decap_8
XFILLER_26_695 VPWR VGND sg13g2_decap_8
XFILLER_41_665 VPWR VGND sg13g2_decap_8
XFILLER_15_62 VPWR VGND sg13g2_fill_2
XFILLER_5_511 VPWR VGND sg13g2_decap_8
XFILLER_5_588 VPWR VGND sg13g2_decap_8
XFILLER_49_743 VPWR VGND sg13g2_decap_8
XFILLER_0_260 VPWR VGND sg13g2_fill_1
XFILLER_1_794 VPWR VGND sg13g2_decap_8
XFILLER_37_905 VPWR VGND sg13g2_decap_8
XFILLER_48_297 VPWR VGND sg13g2_decap_8
X_3930_ _1358_ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] _1316_
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_17_662 VPWR VGND sg13g2_decap_8
XFILLER_44_470 VPWR VGND sg13g2_decap_8
XFILLER_32_643 VPWR VGND sg13g2_decap_8
X_3861_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[7\] _1290_
+ _1295_ _1294_ sg13g2_a21oi_1
X_2812_ _0372_ _0347_ _0371_ VPWR VGND sg13g2_nand2_1
X_3792_ net662 VPWR _1249_ VGND _0834_ _1040_ sg13g2_o21ai_1
X_2743_ net728 _1715_ _1616_ _0304_ VPWR VGND sg13g2_nand3_1
XFILLER_9_861 VPWR VGND sg13g2_decap_8
XFILLER_8_393 VPWR VGND sg13g2_fill_2
X_2674_ net741 net766 _1521_ sap_3_inst.clock.hlt VPWR VGND sg13g2_nor3_1
X_3226_ _0749_ _0751_ _0743_ _0754_ VPWR VGND sg13g2_nand3_1
X_3157_ _0685_ _1535_ _0636_ VPWR VGND sg13g2_nand2_2
XFILLER_27_426 VPWR VGND sg13g2_fill_2
XFILLER_28_938 VPWR VGND sg13g2_decap_8
X_2108_ net776 net781 _1528_ VPWR VGND sg13g2_nor2_2
XFILLER_27_448 VPWR VGND sg13g2_decap_8
X_3088_ VGND VPWR net725 _0615_ _0616_ _1516_ sg13g2_a21oi_1
XFILLER_42_429 VPWR VGND sg13g2_decap_8
XFILLER_23_610 VPWR VGND sg13g2_decap_8
X_2039_ VPWR _1461_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[1\] VGND
+ sg13g2_inv_1
XFILLER_35_1018 VPWR VGND sg13g2_decap_8
XFILLER_23_687 VPWR VGND sg13g2_decap_8
XFILLER_10_359 VPWR VGND sg13g2_fill_2
XFILLER_2_525 VPWR VGND sg13g2_decap_8
Xfanout840 net849 net840 VPWR VGND sg13g2_buf_8
XFILLER_46_702 VPWR VGND sg13g2_decap_8
XFILLER_19_927 VPWR VGND sg13g2_decap_8
XFILLER_46_779 VPWR VGND sg13g2_decap_8
XFILLER_14_632 VPWR VGND sg13g2_decap_8
XFILLER_26_492 VPWR VGND sg13g2_decap_8
XFILLER_42_996 VPWR VGND sg13g2_decap_8
XFILLER_41_462 VPWR VGND sg13g2_decap_8
XFILLER_13_175 VPWR VGND sg13g2_fill_2
XFILLER_6_831 VPWR VGND sg13g2_decap_8
XFILLER_10_893 VPWR VGND sg13g2_decap_8
X_2390_ _1810_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] net637
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_49_540 VPWR VGND sg13g2_decap_8
XFILLER_1_591 VPWR VGND sg13g2_decap_8
X_4060_ net833 VGND VPWR _0028_ sap_3_inst.alu.flags\[3\] net41 sg13g2_dfrbpq_1
XFILLER_3_1027 VPWR VGND sg13g2_fill_2
XFILLER_3_1016 VPWR VGND sg13g2_decap_8
X_3011_ VPWR VGND _0329_ _0564_ _0563_ _1944_ _0565_ _0544_ sg13g2_a221oi_1
XFILLER_37_702 VPWR VGND sg13g2_decap_8
XFILLER_36_234 VPWR VGND sg13g2_fill_2
XFILLER_37_779 VPWR VGND sg13g2_decap_8
X_3913_ _1343_ _1314_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] _1301_
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_952 VPWR VGND sg13g2_decap_8
X_3844_ _1280_ _1278_ _1282_ _0155_ VPWR VGND sg13g2_a21o_2
XFILLER_20_668 VPWR VGND sg13g2_decap_8
X_3775_ _1235_ VPWR _0133_ VGND _1448_ net661 sg13g2_o21ai_1
X_2726_ _1539_ VPWR _0297_ VGND _1544_ _0296_ sg13g2_o21ai_1
X_2657_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] net643
+ net631 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] _0244_ net650 sg13g2_a221oi_1
X_2588_ _1998_ net629 _1997_ VPWR VGND sg13g2_nand2_1
X_3209_ _0737_ net668 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] net670
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_41_1022 VPWR VGND sg13g2_decap_8
X_4189_ net827 VGND VPWR _0153_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_27_234 VPWR VGND sg13g2_fill_1
XFILLER_28_735 VPWR VGND sg13g2_decap_8
XFILLER_43_749 VPWR VGND sg13g2_decap_8
XFILLER_24_930 VPWR VGND sg13g2_decap_8
XFILLER_23_484 VPWR VGND sg13g2_decap_8
XFILLER_11_657 VPWR VGND sg13g2_decap_8
XFILLER_7_628 VPWR VGND sg13g2_decap_8
XFILLER_6_105 VPWR VGND sg13g2_fill_1
XFILLER_3_834 VPWR VGND sg13g2_decap_8
XFILLER_19_724 VPWR VGND sg13g2_decap_8
Xfanout692 net696 net692 VPWR VGND sg13g2_buf_8
Xfanout681 _0660_ net681 VPWR VGND sg13g2_buf_2
Xfanout670 net673 net670 VPWR VGND sg13g2_buf_8
XFILLER_46_576 VPWR VGND sg13g2_decap_8
XFILLER_34_738 VPWR VGND sg13g2_decap_8
XFILLER_15_952 VPWR VGND sg13g2_decap_8
XFILLER_30_933 VPWR VGND sg13g2_decap_8
XFILLER_42_793 VPWR VGND sg13g2_decap_8
X_3560_ net585 _1071_ _1072_ _1073_ VPWR VGND sg13g2_nor3_1
XFILLER_10_690 VPWR VGND sg13g2_decap_8
X_2511_ _1925_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] net640
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3491_ net591 _0978_ _1007_ _1013_ VPWR VGND sg13g2_nor3_1
X_2442_ _1862_ net647 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] _1730_
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2373_ net776 _1792_ _1793_ VPWR VGND sg13g2_nor2_1
X_4112_ net842 VGND VPWR _0076_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\]
+ clknet_5_30__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_37_576 VPWR VGND sg13g2_decap_8
XFILLER_21_900 VPWR VGND sg13g2_decap_8
XFILLER_21_977 VPWR VGND sg13g2_decap_8
X_3827_ VPWR VGND net711 net610 _0995_ net602 _1270_ _0980_ sg13g2_a221oi_1
X_3758_ net653 _1220_ _1221_ VPWR VGND sg13g2_nor2_1
X_2709_ net576 _0213_ net10 VPWR VGND sg13g2_and2_1
X_3689_ VPWR VGND net601 net18 _0898_ net588 _1176_ _0872_ sg13g2_a221oi_1
XFILLER_0_815 VPWR VGND sg13g2_decap_8
XFILLER_48_808 VPWR VGND sg13g2_decap_8
XFILLER_28_532 VPWR VGND sg13g2_decap_8
XFILLER_15_226 VPWR VGND sg13g2_fill_1
XFILLER_16_738 VPWR VGND sg13g2_decap_8
XFILLER_43_546 VPWR VGND sg13g2_decap_8
XFILLER_23_281 VPWR VGND sg13g2_fill_2
XFILLER_8_915 VPWR VGND sg13g2_decap_8
XFILLER_7_403 VPWR VGND sg13g2_fill_1
XFILLER_12_966 VPWR VGND sg13g2_decap_8
XFILLER_3_631 VPWR VGND sg13g2_decap_8
XFILLER_47_830 VPWR VGND sg13g2_decap_8
XFILLER_19_521 VPWR VGND sg13g2_decap_8
XFILLER_46_373 VPWR VGND sg13g2_decap_8
XFILLER_19_598 VPWR VGND sg13g2_decap_8
XFILLER_34_535 VPWR VGND sg13g2_decap_8
X_2991_ net787 sap_3_inst.alu.tmp\[7\] _0545_ VPWR VGND sg13g2_nor2_1
XFILLER_42_590 VPWR VGND sg13g2_decap_8
XFILLER_9_53 VPWR VGND sg13g2_fill_2
XFILLER_30_730 VPWR VGND sg13g2_decap_8
XFILLER_9_64 VPWR VGND sg13g2_fill_2
X_3612_ _1040_ _1116_ net602 _1117_ VPWR VGND sg13g2_nand3_1
XFILLER_7_992 VPWR VGND sg13g2_decap_8
X_3543_ _1058_ VPWR _1059_ VGND net605 _0963_ sg13g2_o21ai_1
X_3474_ net711 VPWR _0997_ VGND net669 _0990_ sg13g2_o21ai_1
X_2425_ _1844_ VPWR _1845_ VGND _1724_ _1727_ sg13g2_o21ai_1
XFILLER_9_1022 VPWR VGND sg13g2_decap_8
X_2356_ _1774_ _1775_ _1700_ _1776_ VPWR VGND sg13g2_nand3_1
X_2287_ _1701_ VPWR _1707_ VGND net765 _1706_ sg13g2_o21ai_1
X_4026_ _1429_ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\] sap_3_inst.reg_file.array_serializer_inst.word_index\[1\]
+ _1431_ VPWR VGND sg13g2_a21o_1
XFILLER_38_863 VPWR VGND sg13g2_decap_8
XFILLER_25_568 VPWR VGND sg13g2_decap_8
XFILLER_40_527 VPWR VGND sg13g2_decap_8
XFILLER_21_774 VPWR VGND sg13g2_decap_8
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_612 VPWR VGND sg13g2_decap_8
XFILLER_48_605 VPWR VGND sg13g2_decap_8
XFILLER_0_689 VPWR VGND sg13g2_decap_8
XFILLER_29_874 VPWR VGND sg13g2_decap_8
XFILLER_44_855 VPWR VGND sg13g2_decap_8
XFILLER_16_535 VPWR VGND sg13g2_decap_8
XFILLER_31_549 VPWR VGND sg13g2_decap_8
XFILLER_8_712 VPWR VGND sg13g2_decap_8
XFILLER_12_763 VPWR VGND sg13g2_decap_8
XFILLER_34_83 VPWR VGND sg13g2_fill_1
XFILLER_8_789 VPWR VGND sg13g2_decap_8
XFILLER_7_244 VPWR VGND sg13g2_fill_2
XFILLER_4_984 VPWR VGND sg13g2_decap_8
X_2210_ _1630_ net743 _1629_ VPWR VGND sg13g2_nand2_2
X_3190_ _0713_ VPWR _0718_ VGND _1495_ net613 sg13g2_o21ai_1
X_2141_ _1561_ net742 net734 VPWR VGND sg13g2_nand2_1
XFILLER_39_649 VPWR VGND sg13g2_decap_8
X_2072_ _1494_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[7\] VPWR VGND
+ sg13g2_inv_2
XFILLER_35_822 VPWR VGND sg13g2_decap_8
XFILLER_35_899 VPWR VGND sg13g2_decap_8
X_2974_ _0529_ net790 net720 VPWR VGND sg13g2_nand2_1
XFILLER_22_538 VPWR VGND sg13g2_decap_8
X_3526_ net31 _0874_ _1045_ _1046_ VPWR VGND sg13g2_nor3_2
X_3457_ _0980_ _0956_ _0977_ VPWR VGND sg13g2_xnor2_1
X_2408_ VGND VPWR net733 _1647_ _1828_ _1605_ sg13g2_a21oi_1
X_3388_ _0907_ _0885_ _0914_ VPWR VGND sg13g2_xor2_1
X_2339_ _1741_ VPWR _1759_ VGND _1756_ _1758_ sg13g2_o21ai_1
X_4009_ _1415_ VPWR _1418_ VGND _1439_ _1416_ sg13g2_o21ai_1
XFILLER_26_800 VPWR VGND sg13g2_decap_8
XFILLER_38_660 VPWR VGND sg13g2_decap_8
XFILLER_25_310 VPWR VGND sg13g2_fill_1
XFILLER_26_877 VPWR VGND sg13g2_decap_8
XFILLER_41_847 VPWR VGND sg13g2_decap_8
XFILLER_21_571 VPWR VGND sg13g2_decap_8
XFILLER_49_925 VPWR VGND sg13g2_decap_8
XFILLER_48_402 VPWR VGND sg13g2_decap_8
XFILLER_1_976 VPWR VGND sg13g2_decap_8
XFILLER_0_486 VPWR VGND sg13g2_decap_8
XFILLER_36_619 VPWR VGND sg13g2_decap_8
XFILLER_48_479 VPWR VGND sg13g2_decap_8
XFILLER_29_671 VPWR VGND sg13g2_decap_8
XFILLER_16_310 VPWR VGND sg13g2_fill_1
XFILLER_17_844 VPWR VGND sg13g2_decap_8
XFILLER_44_652 VPWR VGND sg13g2_decap_8
XFILLER_32_825 VPWR VGND sg13g2_decap_8
XFILLER_31_335 VPWR VGND sg13g2_fill_2
XFILLER_40_891 VPWR VGND sg13g2_decap_8
XFILLER_12_560 VPWR VGND sg13g2_decap_8
X_2690_ _0265_ _0269_ _1825_ _0273_ VPWR VGND _0272_ sg13g2_nand4_1
XFILLER_8_586 VPWR VGND sg13g2_decap_8
X_3311_ _0839_ _0742_ _0837_ VPWR VGND sg13g2_nand2_1
XFILLER_4_781 VPWR VGND sg13g2_decap_8
X_3242_ net703 net700 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] _0770_
+ VPWR VGND net693 sg13g2_nand4_1
X_3173_ _0701_ net664 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] net665
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2124_ net756 VPWR _1544_ VGND net740 _1541_ sg13g2_o21ai_1
Xclkbuf_5_30__f_sap_3_inst.alu.clk_regs clknet_4_15_0_sap_3_inst.alu.clk_regs clknet_5_30__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2055_ VPWR _1477_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_35_696 VPWR VGND sg13g2_decap_8
XFILLER_10_508 VPWR VGND sg13g2_decap_8
XFILLER_23_869 VPWR VGND sg13g2_decap_8
X_2957_ net794 sap_3_inst.alu.tmp\[5\] _0512_ VPWR VGND sg13g2_nor2b_1
X_2888_ _0445_ net796 net720 VPWR VGND sg13g2_xnor2_1
XFILLER_2_707 VPWR VGND sg13g2_decap_8
X_3509_ _1028_ _1029_ _1030_ VPWR VGND sg13g2_nor2_1
XFILLER_17_118 VPWR VGND sg13g2_fill_1
XFILLER_45_438 VPWR VGND sg13g2_decap_8
XFILLER_14_814 VPWR VGND sg13g2_decap_8
XFILLER_26_674 VPWR VGND sg13g2_decap_8
XFILLER_41_644 VPWR VGND sg13g2_decap_8
XFILLER_13_346 VPWR VGND sg13g2_fill_2
XFILLER_12_1008 VPWR VGND sg13g2_decap_8
XFILLER_5_567 VPWR VGND sg13g2_decap_8
XFILLER_49_722 VPWR VGND sg13g2_decap_8
XFILLER_1_773 VPWR VGND sg13g2_decap_8
XFILLER_49_799 VPWR VGND sg13g2_decap_8
XFILLER_48_276 VPWR VGND sg13g2_decap_8
XFILLER_17_641 VPWR VGND sg13g2_decap_8
XFILLER_32_622 VPWR VGND sg13g2_decap_8
X_3860_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\] VPWR _1294_ VGND sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\]
+ _1293_ sg13g2_o21ai_1
X_2811_ _0371_ _0322_ _0357_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_165 VPWR VGND sg13g2_decap_4
XFILLER_32_699 VPWR VGND sg13g2_decap_8
X_3791_ VPWR VGND net713 _1068_ _1247_ _0872_ _1248_ _1246_ sg13g2_a221oi_1
XFILLER_9_840 VPWR VGND sg13g2_decap_8
X_2742_ _1551_ _1742_ _0303_ VPWR VGND sg13g2_and2_1
X_2673_ _0231_ VPWR _0025_ VGND _0230_ _0258_ sg13g2_o21ai_1
XFILLER_28_1015 VPWR VGND sg13g2_decap_8
X_3225_ _0745_ VPWR _0753_ VGND _1477_ _0661_ sg13g2_o21ai_1
XFILLER_39_221 VPWR VGND sg13g2_fill_1
X_3156_ VPWR VGND _0683_ _0275_ _0675_ _1623_ _0684_ _0668_ sg13g2_a221oi_1
XFILLER_27_405 VPWR VGND sg13g2_decap_8
XFILLER_28_917 VPWR VGND sg13g2_decap_8
X_2107_ VGND VPWR _1527_ net772 net774 sg13g2_or2_1
X_3087_ net741 _1594_ _0615_ VPWR VGND sg13g2_nor2_1
XFILLER_42_408 VPWR VGND sg13g2_decap_8
X_2038_ _1460_ net796 VPWR VGND sg13g2_inv_2
XFILLER_36_983 VPWR VGND sg13g2_decap_8
XFILLER_35_493 VPWR VGND sg13g2_decap_8
XFILLER_23_666 VPWR VGND sg13g2_decap_8
XFILLER_11_839 VPWR VGND sg13g2_decap_8
X_3989_ _1402_ VPWR _0180_ VGND net582 _1401_ sg13g2_o21ai_1
XFILLER_2_504 VPWR VGND sg13g2_decap_8
Xfanout830 rst_n net830 VPWR VGND sg13g2_buf_8
Xfanout841 net842 net841 VPWR VGND sg13g2_buf_8
XFILLER_19_906 VPWR VGND sg13g2_decap_8
XFILLER_46_758 VPWR VGND sg13g2_decap_8
XFILLER_14_611 VPWR VGND sg13g2_decap_8
XFILLER_26_471 VPWR VGND sg13g2_decap_8
XFILLER_27_994 VPWR VGND sg13g2_decap_8
XFILLER_42_975 VPWR VGND sg13g2_decap_8
XFILLER_41_441 VPWR VGND sg13g2_decap_8
XFILLER_14_688 VPWR VGND sg13g2_decap_8
XFILLER_6_810 VPWR VGND sg13g2_decap_8
XFILLER_10_872 VPWR VGND sg13g2_decap_8
XFILLER_5_320 VPWR VGND sg13g2_fill_1
XFILLER_6_887 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_3_55 VPWR VGND sg13g2_decap_4
XFILLER_1_570 VPWR VGND sg13g2_decap_8
X_3010_ _0560_ VPWR _0564_ VGND _0327_ _0553_ sg13g2_o21ai_1
XFILLER_49_596 VPWR VGND sg13g2_decap_8
XFILLER_37_758 VPWR VGND sg13g2_decap_8
XFILLER_18_994 VPWR VGND sg13g2_decap_8
XFILLER_24_419 VPWR VGND sg13g2_decap_8
XFILLER_33_931 VPWR VGND sg13g2_decap_8
X_3912_ _1342_ net810 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] _1300_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\] VPWR VGND sg13g2_a22oi_1
X_3843_ net75 sap_3_inst.reg_file.array_serializer_inst.state\[0\] _1282_ VPWR VGND
+ sg13g2_nor2b_1
XFILLER_20_647 VPWR VGND sg13g2_decap_8
XFILLER_32_496 VPWR VGND sg13g2_decap_8
X_3774_ _1231_ VPWR _1235_ VGND _1233_ _1234_ sg13g2_o21ai_1
X_2725_ VGND VPWR _0292_ _0295_ _0296_ _1556_ sg13g2_a21oi_1
X_2656_ _0243_ _0240_ _0242_ _1858_ net1 VPWR VGND sg13g2_a22oi_1
X_2587_ _1997_ sap_3_inst.alu.flags\[2\] _1839_ VPWR VGND sg13g2_nand2_1
XFILLER_41_1001 VPWR VGND sg13g2_decap_8
X_4188_ net825 VGND VPWR _0152_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\]
+ clknet_5_11__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3208_ _0736_ net656 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] net663
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_28_714 VPWR VGND sg13g2_decap_8
X_3139_ _1787_ net719 _0667_ VPWR VGND _0621_ sg13g2_nand3b_1
Xclkbuf_5_27__f_sap_3_inst.alu.clk_regs clknet_4_13_0_sap_3_inst.alu.clk_regs clknet_5_27__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_43_728 VPWR VGND sg13g2_decap_8
XFILLER_36_780 VPWR VGND sg13g2_decap_8
XFILLER_23_463 VPWR VGND sg13g2_decap_8
XFILLER_24_986 VPWR VGND sg13g2_decap_8
XFILLER_7_607 VPWR VGND sg13g2_decap_8
XFILLER_11_636 VPWR VGND sg13g2_decap_8
XFILLER_3_813 VPWR VGND sg13g2_decap_8
Xfanout660 _0702_ net660 VPWR VGND sg13g2_buf_8
Xfanout682 _0340_ net682 VPWR VGND sg13g2_buf_8
XFILLER_19_703 VPWR VGND sg13g2_decap_8
Xfanout671 net673 net671 VPWR VGND sg13g2_buf_8
Xfanout693 net696 net693 VPWR VGND sg13g2_buf_1
XFILLER_46_555 VPWR VGND sg13g2_decap_8
XFILLER_34_717 VPWR VGND sg13g2_decap_8
XFILLER_15_931 VPWR VGND sg13g2_decap_8
XFILLER_27_791 VPWR VGND sg13g2_decap_8
XFILLER_42_772 VPWR VGND sg13g2_decap_8
XFILLER_30_912 VPWR VGND sg13g2_decap_8
XFILLER_30_989 VPWR VGND sg13g2_decap_8
X_2510_ _1923_ VPWR _1924_ VGND net797 net628 sg13g2_o21ai_1
X_3490_ _0978_ _1007_ _1012_ VPWR VGND sg13g2_nor2_1
X_2441_ _1861_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] net645
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_684 VPWR VGND sg13g2_decap_8
X_2372_ net752 _1642_ net755 _1792_ VPWR VGND sg13g2_nand3_1
X_4111_ net820 VGND VPWR _0075_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\]
+ clknet_5_1__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_49_393 VPWR VGND sg13g2_decap_8
XFILLER_37_555 VPWR VGND sg13g2_decap_8
XFILLER_40_709 VPWR VGND sg13g2_decap_8
XFILLER_18_791 VPWR VGND sg13g2_decap_8
XFILLER_21_956 VPWR VGND sg13g2_decap_8
X_3826_ _0150_ _1154_ _1269_ net608 _1475_ VPWR VGND sg13g2_a22oi_1
X_3757_ net660 net588 _1220_ VPWR VGND sg13g2_nor2_1
X_2708_ VPWR VGND _0238_ _1673_ _0235_ _1468_ net9 net650 sg13g2_a221oi_1
X_3688_ net579 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] _1175_ _0106_
+ VPWR VGND sg13g2_a21o_1
X_2639_ net18 _0227_ VPWR VGND sg13g2_inv_4
XFILLER_47_319 VPWR VGND sg13g2_decap_8
XFILLER_28_511 VPWR VGND sg13g2_decap_8
XFILLER_43_525 VPWR VGND sg13g2_decap_8
XFILLER_16_717 VPWR VGND sg13g2_decap_8
XFILLER_28_588 VPWR VGND sg13g2_decap_8
XFILLER_12_945 VPWR VGND sg13g2_decap_8
XFILLER_24_783 VPWR VGND sg13g2_decap_8
XFILLER_48_1018 VPWR VGND sg13g2_decap_8
XFILLER_3_610 VPWR VGND sg13g2_decap_8
XFILLER_3_687 VPWR VGND sg13g2_decap_8
XFILLER_46_352 VPWR VGND sg13g2_decap_8
XFILLER_47_886 VPWR VGND sg13g2_decap_8
XFILLER_0_45 VPWR VGND sg13g2_fill_2
XFILLER_19_577 VPWR VGND sg13g2_decap_8
XFILLER_34_514 VPWR VGND sg13g2_decap_8
X_2990_ _0544_ _0542_ _0543_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_208 VPWR VGND sg13g2_fill_2
XFILLER_9_43 VPWR VGND sg13g2_fill_1
X_3611_ _1116_ net619 _1042_ VPWR VGND sg13g2_nand2_1
XFILLER_30_786 VPWR VGND sg13g2_decap_8
XFILLER_31_1011 VPWR VGND sg13g2_decap_8
XFILLER_7_971 VPWR VGND sg13g2_decap_8
X_3542_ net601 VPWR _1058_ VGND net663 _0958_ sg13g2_o21ai_1
X_3473_ net712 _0995_ _0996_ VPWR VGND sg13g2_nor2_1
X_2424_ _1844_ net731 _1843_ VPWR VGND sg13g2_nand2_1
XFILLER_9_1001 VPWR VGND sg13g2_decap_8
X_2355_ _1553_ _1676_ net783 _1775_ VPWR VGND sg13g2_nand3_1
X_2286_ _1706_ net749 _1705_ VPWR VGND sg13g2_nand2_1
X_4025_ _1430_ _1429_ _1302_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_842 VPWR VGND sg13g2_decap_8
XFILLER_25_547 VPWR VGND sg13g2_decap_8
XFILLER_40_506 VPWR VGND sg13g2_decap_8
XFILLER_21_753 VPWR VGND sg13g2_decap_8
X_3809_ net613 _1071_ _1072_ _1258_ VPWR VGND sg13g2_nor3_1
XFILLER_0_668 VPWR VGND sg13g2_decap_8
XFILLER_29_853 VPWR VGND sg13g2_decap_8
XFILLER_44_834 VPWR VGND sg13g2_decap_8
XFILLER_16_514 VPWR VGND sg13g2_decap_8
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_24_580 VPWR VGND sg13g2_decap_8
XFILLER_31_528 VPWR VGND sg13g2_decap_8
XFILLER_34_73 VPWR VGND sg13g2_fill_1
XFILLER_12_742 VPWR VGND sg13g2_decap_8
XFILLER_7_201 VPWR VGND sg13g2_fill_2
XFILLER_8_768 VPWR VGND sg13g2_decap_8
XFILLER_4_963 VPWR VGND sg13g2_decap_8
XFILLER_3_484 VPWR VGND sg13g2_decap_8
X_2140_ _1560_ net755 net754 VPWR VGND sg13g2_nand2_1
XFILLER_39_628 VPWR VGND sg13g2_decap_8
X_2071_ VPWR _1493_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_47_683 VPWR VGND sg13g2_decap_8
XFILLER_35_801 VPWR VGND sg13g2_decap_8
XFILLER_22_517 VPWR VGND sg13g2_decap_8
XFILLER_35_878 VPWR VGND sg13g2_decap_8
X_2973_ VPWR VGND _0527_ net575 _0526_ _0326_ _0528_ _0516_ sg13g2_a221oi_1
XFILLER_30_583 VPWR VGND sg13g2_decap_8
X_3525_ net590 net605 _1045_ VPWR VGND sg13g2_nor2_1
X_3456_ _0979_ _0977_ _0956_ VPWR VGND sg13g2_nand2b_1
X_2407_ net748 _1647_ _1827_ VPWR VGND sg13g2_nor2_1
X_3387_ _0913_ _0885_ _0907_ VPWR VGND sg13g2_nand2_1
X_2338_ _1752_ _1754_ _1751_ _1758_ VPWR VGND _1757_ sg13g2_nand4_1
X_2269_ _1688_ VPWR _1689_ VGND _1604_ _1659_ sg13g2_o21ai_1
X_4008_ _1417_ _1415_ _1416_ VPWR VGND sg13g2_nand2_1
XFILLER_26_856 VPWR VGND sg13g2_decap_8
XFILLER_38_1017 VPWR VGND sg13g2_decap_8
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_826 VPWR VGND sg13g2_decap_8
XFILLER_21_550 VPWR VGND sg13g2_decap_8
XFILLER_5_749 VPWR VGND sg13g2_decap_8
XFILLER_49_904 VPWR VGND sg13g2_decap_8
XFILLER_1_955 VPWR VGND sg13g2_decap_8
XFILLER_48_458 VPWR VGND sg13g2_decap_8
XFILLER_17_823 VPWR VGND sg13g2_decap_8
XFILLER_29_650 VPWR VGND sg13g2_decap_8
XFILLER_44_631 VPWR VGND sg13g2_decap_8
XFILLER_32_804 VPWR VGND sg13g2_decap_8
XFILLER_40_870 VPWR VGND sg13g2_decap_8
Xclkbuf_5_1__f_sap_3_inst.alu.clk_regs clknet_4_0_0_sap_3_inst.alu.clk_regs clknet_5_1__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_8_565 VPWR VGND sg13g2_decap_8
XFILLER_4_760 VPWR VGND sg13g2_decap_8
X_3310_ _0755_ _0766_ _0775_ net588 _0838_ VPWR VGND sg13g2_or4_1
X_3241_ net701 net692 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] _0769_
+ VPWR VGND net688 sg13g2_nand4_1
X_3172_ net691 net687 net697 _0700_ VPWR VGND sg13g2_nand3_1
X_2123_ _1523_ _1542_ net765 _1543_ VPWR VGND sg13g2_nand3_1
XFILLER_27_609 VPWR VGND sg13g2_decap_8
XFILLER_47_480 VPWR VGND sg13g2_decap_8
X_2054_ VPWR _1476_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_35_675 VPWR VGND sg13g2_decap_8
XFILLER_23_848 VPWR VGND sg13g2_decap_8
X_2956_ _0511_ net791 sap_3_inst.alu.tmp\[6\] VPWR VGND sg13g2_xnor2_1
X_2887_ net32 net627 _0444_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_892 VPWR VGND sg13g2_decap_8
Xclkbuf_0_sap_3_inst.alu.clk_regs sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3508_ VGND VPWR _0992_ _1007_ _1029_ _1027_ sg13g2_a21oi_1
X_3439_ _0963_ _0755_ _0802_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_609 VPWR VGND sg13g2_decap_8
XFILLER_45_417 VPWR VGND sg13g2_decap_8
XFILLER_39_992 VPWR VGND sg13g2_decap_8
XFILLER_26_653 VPWR VGND sg13g2_decap_8
XFILLER_41_623 VPWR VGND sg13g2_decap_8
XFILLER_22_881 VPWR VGND sg13g2_decap_8
XFILLER_40_188 VPWR VGND sg13g2_fill_2
XFILLER_5_546 VPWR VGND sg13g2_decap_8
Xoutput30 net30 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_752 VPWR VGND sg13g2_decap_8
XFILLER_49_701 VPWR VGND sg13g2_decap_8
XFILLER_49_778 VPWR VGND sg13g2_decap_8
XFILLER_17_620 VPWR VGND sg13g2_decap_8
XFILLER_45_984 VPWR VGND sg13g2_decap_8
XFILLER_16_163 VPWR VGND sg13g2_fill_2
XFILLER_17_697 VPWR VGND sg13g2_decap_8
XFILLER_32_601 VPWR VGND sg13g2_decap_8
X_2810_ _0323_ _0356_ net762 _0370_ VPWR VGND sg13g2_nand3_1
XFILLER_20_829 VPWR VGND sg13g2_decap_8
XFILLER_32_678 VPWR VGND sg13g2_decap_8
X_3790_ _0702_ net654 _0289_ _1247_ VPWR VGND sg13g2_nand3_1
X_2741_ net748 VPWR _0302_ VGND net763 _1570_ sg13g2_o21ai_1
XFILLER_9_896 VPWR VGND sg13g2_decap_8
X_2672_ _0257_ VPWR _0258_ VGND _1868_ net31 sg13g2_o21ai_1
X_3224_ _0746_ _0747_ _0744_ _0752_ VPWR VGND _0750_ sg13g2_nand4_1
.ends

