module heichips25_template (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net38;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire \sap_3_inst.alu.clk_regs ;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire clk_div_out;
 wire mem_mar_we;
 wire mem_ram_we;
 wire regFile_serial;
 wire regFile_serial_start;
 wire \sap_3_inst.alu.acc[0] ;
 wire \sap_3_inst.alu.acc[1] ;
 wire \sap_3_inst.alu.acc[2] ;
 wire \sap_3_inst.alu.acc[3] ;
 wire \sap_3_inst.alu.acc[4] ;
 wire \sap_3_inst.alu.acc[5] ;
 wire \sap_3_inst.alu.acc[6] ;
 wire \sap_3_inst.alu.acc[7] ;
 wire \sap_3_inst.alu.act[0] ;
 wire \sap_3_inst.alu.act[1] ;
 wire \sap_3_inst.alu.act[2] ;
 wire \sap_3_inst.alu.act[3] ;
 wire \sap_3_inst.alu.act[4] ;
 wire \sap_3_inst.alu.act[5] ;
 wire \sap_3_inst.alu.act[6] ;
 wire \sap_3_inst.alu.act[7] ;
 wire \sap_3_inst.alu.carry ;
 wire \sap_3_inst.alu.clk ;
 wire \sap_3_inst.alu.flags[0] ;
 wire \sap_3_inst.alu.flags[1] ;
 wire \sap_3_inst.alu.flags[2] ;
 wire \sap_3_inst.alu.flags[3] ;
 wire \sap_3_inst.alu.flags[4] ;
 wire \sap_3_inst.alu.flags[5] ;
 wire \sap_3_inst.alu.flags[6] ;
 wire \sap_3_inst.alu.flags[7] ;
 wire \sap_3_inst.alu.tmp[0] ;
 wire \sap_3_inst.alu.tmp[1] ;
 wire \sap_3_inst.alu.tmp[2] ;
 wire \sap_3_inst.alu.tmp[3] ;
 wire \sap_3_inst.alu.tmp[4] ;
 wire \sap_3_inst.alu.tmp[5] ;
 wire \sap_3_inst.alu.tmp[6] ;
 wire \sap_3_inst.alu.tmp[7] ;
 wire \sap_3_inst.clock.hlt ;
 wire \sap_3_inst.controller.opcode[0] ;
 wire \sap_3_inst.controller.opcode[1] ;
 wire \sap_3_inst.controller.opcode[2] ;
 wire \sap_3_inst.controller.opcode[3] ;
 wire \sap_3_inst.controller.opcode[4] ;
 wire \sap_3_inst.controller.opcode[5] ;
 wire \sap_3_inst.controller.opcode[6] ;
 wire \sap_3_inst.controller.opcode[7] ;
 wire \sap_3_inst.controller.stage[0] ;
 wire \sap_3_inst.controller.stage[1] ;
 wire \sap_3_inst.controller.stage[2] ;
 wire \sap_3_inst.controller.stage[3] ;
 wire \sap_3_inst.out[0] ;
 wire \sap_3_inst.out[1] ;
 wire \sap_3_inst.out[2] ;
 wire \sap_3_inst.out[3] ;
 wire \sap_3_inst.out[4] ;
 wire \sap_3_inst.out[5] ;
 wire \sap_3_inst.out[6] ;
 wire \sap_3_inst.out[7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.bit_pos[0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.state[0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.state[1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.word_index[0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.word_index[1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.word_index[2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.word_index[3] ;
 wire sap_3_outputReg_serial;
 wire sap_3_outputReg_start_sync;
 wire \u_ser.bit_pos[0] ;
 wire \u_ser.bit_pos[1] ;
 wire \u_ser.bit_pos[2] ;
 wire \u_ser.shadow_reg[0] ;
 wire \u_ser.shadow_reg[1] ;
 wire \u_ser.shadow_reg[2] ;
 wire \u_ser.shadow_reg[3] ;
 wire \u_ser.shadow_reg[4] ;
 wire \u_ser.shadow_reg[5] ;
 wire \u_ser.shadow_reg[6] ;
 wire \u_ser.shadow_reg[7] ;
 wire \u_ser.state[0] ;
 wire \u_ser.state[1] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net36;
 wire net37;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_0_clk_div_out;
 wire clknet_1_0__leaf_clk_div_out;
 wire clknet_1_1__leaf_clk_div_out;
 wire \clknet_leaf_0_sap_3_inst.alu.clk ;
 wire \clknet_leaf_1_sap_3_inst.alu.clk ;
 wire \clknet_leaf_2_sap_3_inst.alu.clk ;
 wire \clknet_0_sap_3_inst.alu.clk ;
 wire \clknet_1_0__leaf_sap_3_inst.alu.clk ;
 wire \clknet_1_1__leaf_sap_3_inst.alu.clk ;
 wire \clknet_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_0_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_1_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_2_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_3_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_4_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_5_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_6_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_7_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_8_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_9_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_10_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_11_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_12_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_13_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_14_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_15_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_0__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_1__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_2__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_3__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_4__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_5__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_6__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_7__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_8__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_9__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_10__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_11__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_12__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_13__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_14__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_15__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_16__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_17__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_18__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_19__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_20__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_21__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_22__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_23__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_24__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_25__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_26__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_27__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_28__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_29__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_30__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_31__leaf_sap_3_inst.alu.clk_regs ;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;

 sg13g2_inv_1 _2015_ (.VDD(VPWR),
    .Y(_1437_),
    .A(\u_ser.state[1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2016_ (.VDD(VPWR),
    .Y(_1438_),
    .A(\u_ser.state[0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2017_ (.VDD(VPWR),
    .Y(_1439_),
    .A(\u_ser.bit_pos[2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2018_ (.VDD(VPWR),
    .Y(_1440_),
    .A(net77),
    .VSS(VGND));
 sg13g2_inv_4 _2019_ (.A(net777),
    .Y(_1441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2020_ (.A(\sap_3_inst.controller.opcode[4] ),
    .Y(_1442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2021_ (.Y(_1443_),
    .A(net768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2022_ (.A(net780),
    .Y(_1444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2023_ (.Y(_1445_),
    .A(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2024_ (.Y(_1446_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2025_ (.VDD(VPWR),
    .Y(_1447_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2026_ (.VDD(VPWR),
    .Y(_1448_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2027_ (.VDD(VPWR),
    .Y(_1449_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2028_ (.VDD(VPWR),
    .Y(_1450_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2029_ (.VDD(VPWR),
    .Y(_1451_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2030_ (.VDD(VPWR),
    .Y(_1452_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2031_ (.VDD(VPWR),
    .Y(_1453_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2032_ (.VDD(VPWR),
    .Y(_1454_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2033_ (.VDD(VPWR),
    .Y(_1455_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2034_ (.VDD(VPWR),
    .Y(_1456_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2035_ (.VDD(VPWR),
    .Y(_1457_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .VSS(VGND));
 sg13g2_inv_2 _2036_ (.Y(_1458_),
    .A(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2037_ (.VDD(VPWR),
    .Y(_1459_),
    .A(net805),
    .VSS(VGND));
 sg13g2_inv_2 _2038_ (.Y(_1460_),
    .A(net796),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2039_ (.VDD(VPWR),
    .Y(_1461_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2040_ (.VDD(VPWR),
    .Y(_1462_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2041_ (.VDD(VPWR),
    .Y(_1463_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2042_ (.VDD(VPWR),
    .Y(_1464_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2043_ (.VDD(VPWR),
    .Y(_1465_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2044_ (.VDD(VPWR),
    .Y(_1466_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2045_ (.VDD(VPWR),
    .Y(_1467_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .VSS(VGND));
 sg13g2_inv_4 _2046_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[0][0] ),
    .Y(_1468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2047_ (.VDD(VPWR),
    .Y(_1469_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2048_ (.VDD(VPWR),
    .Y(_1470_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2049_ (.VDD(VPWR),
    .Y(_1471_),
    .A(\sap_3_inst.alu.tmp[2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2050_ (.VDD(VPWR),
    .Y(_1472_),
    .A(\sap_3_inst.alu.tmp[3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2051_ (.VDD(VPWR),
    .Y(_1473_),
    .A(\sap_3_inst.alu.tmp[4] ),
    .VSS(VGND));
 sg13g2_inv_2 _2052_ (.Y(_1474_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2053_ (.VDD(VPWR),
    .Y(_1475_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2054_ (.VDD(VPWR),
    .Y(_1476_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2055_ (.VDD(VPWR),
    .Y(_1477_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2056_ (.VDD(VPWR),
    .Y(_1478_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2057_ (.VDD(VPWR),
    .Y(_1479_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2058_ (.VDD(VPWR),
    .Y(_1480_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2059_ (.VDD(VPWR),
    .Y(_1481_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2060_ (.VDD(VPWR),
    .Y(_1482_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2061_ (.VDD(VPWR),
    .Y(_1483_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .VSS(VGND));
 sg13g2_inv_2 _2062_ (.Y(_1484_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2063_ (.VDD(VPWR),
    .Y(_1485_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2064_ (.VDD(VPWR),
    .Y(_1486_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2065_ (.VDD(VPWR),
    .Y(_1487_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2066_ (.VDD(VPWR),
    .Y(_1488_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2067_ (.VDD(VPWR),
    .Y(_1489_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2068_ (.VDD(VPWR),
    .Y(_1490_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2069_ (.VDD(VPWR),
    .Y(_1491_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2070_ (.VDD(VPWR),
    .Y(_1492_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2071_ (.VDD(VPWR),
    .Y(_1493_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .VSS(VGND));
 sg13g2_inv_2 _2072_ (.Y(_1494_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2073_ (.VDD(VPWR),
    .Y(_1495_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2074_ (.VDD(VPWR),
    .Y(_1496_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2075_ (.VDD(VPWR),
    .Y(_1497_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2076_ (.VDD(VPWR),
    .Y(_1498_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2077_ (.VDD(VPWR),
    .Y(_1499_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2078_ (.VDD(VPWR),
    .Y(_1500_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2079_ (.VDD(VPWR),
    .Y(_1501_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2080_ (.VDD(VPWR),
    .Y(_1502_),
    .A(net60),
    .VSS(VGND));
 sg13g2_inv_1 _2082__2 (.VDD(VPWR),
    .Y(net38),
    .A(\clknet_leaf_0_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4038__3 (.VDD(VPWR),
    .Y(net39),
    .A(\clknet_leaf_1_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_nor2_2 _2083_ (.A(net760),
    .B(net761),
    .Y(_1503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2084_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1504_),
    .B(net761),
    .A(net760));
 sg13g2_nor2_2 _2085_ (.A(\sap_3_inst.controller.stage[3] ),
    .B(net759),
    .Y(_1505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2086_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1506_),
    .B(net759),
    .A(\sap_3_inst.controller.stage[3] ));
 sg13g2_and2_1 _2087_ (.A(net760),
    .B(net761),
    .X(_1507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2088_ (.Y(_1508_),
    .A(\sap_3_inst.controller.stage[1] ),
    .B(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2089_ (.A(_1506_),
    .B(_1508_),
    .Y(_1509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2090_ (.Y(_1510_),
    .A(_1505_),
    .B(_1507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2091_ (.A(\sap_3_inst.controller.opcode[0] ),
    .B_N(net784),
    .Y(_1511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2092_ (.Y(_1512_),
    .B(net782),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net785));
 sg13g2_nand3b_1 _2093_ (.B(net783),
    .C(net781),
    .Y(_1513_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net786));
 sg13g2_nor2b_2 _2094_ (.A(net768),
    .B_N(net770),
    .Y(_1514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2095_ (.Y(_1515_),
    .B(net771),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net769));
 sg13g2_nor2_2 _2096_ (.A(net766),
    .B(_1515_),
    .Y(_1516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2097_ (.Y(_1517_),
    .B(_1514_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net766));
 sg13g2_and2_1 _2098_ (.A(net774),
    .B(net772),
    .X(_1518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2099_ (.Y(_1519_),
    .A(net774),
    .B(net772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2100_ (.A(net778),
    .B(_1515_),
    .C(net763),
    .Y(_1520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2101_ (.B(_1514_),
    .C(_1518_),
    .A(_1441_),
    .Y(_1521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2102_ (.A(net766),
    .B(net756),
    .Y(_1522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2103_ (.A(net768),
    .B(net770),
    .Y(_1523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2104_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1524_),
    .B(net770),
    .A(net769));
 sg13g2_nor2_2 _2105_ (.A(net785),
    .B(net782),
    .Y(_1525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2106_ (.A(net774),
    .B(net772),
    .Y(_1526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2107_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1527_),
    .B(net772),
    .A(net774));
 sg13g2_nor2_2 _2108_ (.A(net776),
    .B(net781),
    .Y(_1528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2109_ (.B(_1525_),
    .C(_1526_),
    .A(_1523_),
    .Y(_1529_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1528_));
 sg13g2_nor2b_2 _2110_ (.A(_1522_),
    .B_N(_1529_),
    .Y(_1530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2111_ (.B1(_1529_),
    .VDD(VPWR),
    .Y(_1531_),
    .VSS(VGND),
    .A1(net767),
    .A2(net756));
 sg13g2_nor2b_2 _2112_ (.A(net760),
    .B_N(net761),
    .Y(_1532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2113_ (.Y(_1533_),
    .A(_1505_),
    .B(_1532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2114_ (.A(net761),
    .B_N(net760),
    .Y(_1534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2115_ (.Y(_1535_),
    .A(_1505_),
    .B(_1534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2116_ (.Y(_1536_),
    .A(net760),
    .B(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2117_ (.B(_1533_),
    .C(_1535_),
    .A(_1530_),
    .Y(_1537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2118_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net740),
    .A2(_1516_),
    .Y(_1538_),
    .B1(_1537_));
 sg13g2_nand2_1 _2119_ (.Y(_1539_),
    .A(net740),
    .B(_1520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2120_ (.A(net776),
    .B_N(net781),
    .Y(_1540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2121_ (.B(_1523_),
    .C(_1525_),
    .A(net765),
    .Y(_1541_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1540_));
 sg13g2_nor4_1 _2122_ (.A(net779),
    .B(_1444_),
    .C(net786),
    .D(net783),
    .Y(_1542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2123_ (.B(_1523_),
    .C(_1542_),
    .A(net765),
    .Y(_1543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2124_ (.B1(net756),
    .VDD(VPWR),
    .Y(_1544_),
    .VSS(VGND),
    .A1(net740),
    .A2(_1541_));
 sg13g2_nor2_1 _2125_ (.A(_1443_),
    .B(net766),
    .Y(_1545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2126_ (.A(_1443_),
    .B(net771),
    .Y(_1546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2127_ (.Y(_1547_),
    .B(net769),
    .A_N(net771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2128_ (.A(net767),
    .B(_1547_),
    .Y(_1548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2129_ (.A(_1444_),
    .B(net784),
    .C(_1524_),
    .Y(_1549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2130_ (.B(_1523_),
    .C(net781),
    .Y(_1550_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net783));
 sg13g2_nor2_2 _2131_ (.A(_1548_),
    .B(_1549_),
    .Y(_1551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2132_ (.Y(_1552_),
    .B(_1550_),
    .A_N(_1548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2133_ (.A(net740),
    .B(_1547_),
    .Y(_1553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2134_ (.Y(_1554_),
    .A(net745),
    .B(_1546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2135_ (.A(net767),
    .B(_1554_),
    .Y(_1555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2136_ (.A(_1551_),
    .B(_1555_),
    .Y(_1556_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2137_ (.A(\sap_3_inst.controller.stage[3] ),
    .B_N(net759),
    .Y(_1557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2138_ (.Y(_1558_),
    .B(net759),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\sap_3_inst.controller.stage[3] ));
 sg13g2_and2_1 _2139_ (.A(net755),
    .B(net754),
    .X(_1559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2140_ (.Y(_1560_),
    .A(net755),
    .B(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2141_ (.Y(_1561_),
    .A(net742),
    .B(net734),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2142_ (.A(net768),
    .B(net770),
    .X(_1562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2143_ (.Y(_1563_),
    .A(net768),
    .B(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2144_ (.B(net780),
    .C(net770),
    .A(net768),
    .Y(_1564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2145_ (.A(net767),
    .B(_1563_),
    .Y(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2146_ (.A(net777),
    .B(net767),
    .C(net763),
    .Y(_1566_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1524_));
 sg13g2_a221oi_1 _2147_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1561_),
    .C1(net736),
    .B1(_1566_),
    .A1(net744),
    .Y(_1567_),
    .A2(_1565_));
 sg13g2_nor2b_2 _2148_ (.A(net782),
    .B_N(net785),
    .Y(_1568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _2149_ (.X(_1569_),
    .A(_1528_),
    .B(_1562_),
    .C(_1568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2150_ (.B(_1562_),
    .C(_1568_),
    .A(_1528_),
    .Y(_1570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2151_ (.A(_1534_),
    .B(net754),
    .X(_1571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2152_ (.Y(_1572_),
    .A(_1534_),
    .B(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2153_ (.Y(_1573_),
    .B1(_1534_),
    .B2(net754),
    .A2(_1507_),
    .A1(_1505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2154_ (.Y(_1574_),
    .A(net742),
    .B(net732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2155_ (.Y(_1575_),
    .B(_1568_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1564_));
 sg13g2_and2_1 _2156_ (.A(_1536_),
    .B(_1557_),
    .X(_1576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2157_ (.Y(_1577_),
    .A(_1536_),
    .B(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2158_ (.A(_1575_),
    .B(net731),
    .Y(_1578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2159_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1569_),
    .A2(_1574_),
    .Y(_1579_),
    .B1(_1578_));
 sg13g2_nand3b_1 _2160_ (.B(net785),
    .C(net779),
    .Y(_1580_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net782));
 sg13g2_nor4_2 _2161_ (.A(net780),
    .B(_1527_),
    .C(_1563_),
    .Y(_1581_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1580_));
 sg13g2_or4_1 _2162_ (.A(net780),
    .B(_1527_),
    .C(_1563_),
    .D(_1580_),
    .X(_1582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2163_ (.A(net785),
    .B(net782),
    .X(_1583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2164_ (.Y(_1584_),
    .A(net786),
    .B(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2165_ (.A(_1563_),
    .B(_1584_),
    .Y(_1585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2166_ (.A(_1526_),
    .B(_1528_),
    .C(_1562_),
    .D(_1583_),
    .X(_1586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2167_ (.B(_1528_),
    .C(_1562_),
    .A(_1526_),
    .Y(_1587_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1583_));
 sg13g2_nand3_1 _2168_ (.B(_1528_),
    .C(_1568_),
    .A(_1523_),
    .Y(_1588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2169_ (.X(_1589_),
    .A(_1582_),
    .B(_1587_),
    .C(net753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2170_ (.A(net768),
    .B(\sap_3_inst.controller.opcode[2] ),
    .C(net771),
    .Y(_1590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2171_ (.A(net768),
    .B(net780),
    .C(net770),
    .X(_1591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2172_ (.A(_1512_),
    .B(_1591_),
    .Y(_1592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2173_ (.A(net774),
    .B_N(net772),
    .Y(_1593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2174_ (.Y(_1594_),
    .B(net773),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net774));
 sg13g2_nor3_2 _2175_ (.A(_1512_),
    .B(_1591_),
    .C(_1594_),
    .Y(_1595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2176_ (.B(_1590_),
    .C(_1593_),
    .A(_1511_),
    .Y(_1596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2177_ (.A(_1512_),
    .B(net764),
    .C(_1591_),
    .Y(_1597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2178_ (.B(net765),
    .C(_1590_),
    .A(_1511_),
    .Y(_1598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2179_ (.A(_1527_),
    .B(_1564_),
    .C(_1580_),
    .Y(_1599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2180_ (.A(_1527_),
    .B(_1564_),
    .C(_1580_),
    .X(_1600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2181_ (.B(_1598_),
    .C(net749),
    .A(net751),
    .Y(_1601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2182_ (.A(net773),
    .B(_1512_),
    .C(_1591_),
    .Y(_1602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2183_ (.B(_1511_),
    .C(_1590_),
    .Y(_1603_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net772));
 sg13g2_nor2_2 _2184_ (.A(_1580_),
    .B(_1591_),
    .Y(_1604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2185_ (.Y(_1605_),
    .B(_1590_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1580_));
 sg13g2_nor3_1 _2186_ (.A(_1592_),
    .B(net750),
    .C(_1604_),
    .Y(_1606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2187_ (.A(_1589_),
    .B(_1606_),
    .X(_1607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2188_ (.A(net785),
    .B(net782),
    .C(_1564_),
    .Y(_1608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2189_ (.B(_1525_),
    .C(_1562_),
    .A(net781),
    .Y(_1609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2190_ (.A(net750),
    .B(_1608_),
    .Y(_1610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2191_ (.Y(_1611_),
    .A(_1600_),
    .B(_1609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2192_ (.A(net780),
    .B(net786),
    .C(_1563_),
    .Y(_1612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2193_ (.A(net780),
    .B(_1512_),
    .C(_1563_),
    .Y(_1613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2194_ (.B(_1511_),
    .C(_1562_),
    .A(_1444_),
    .Y(_1614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2195_ (.A(_1586_),
    .B(_1599_),
    .C(_1608_),
    .Y(_1615_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1613_));
 sg13g2_nor2_1 _2196_ (.A(net766),
    .B(_1524_),
    .Y(_1616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2197_ (.Y(_1617_),
    .B(_1523_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net767));
 sg13g2_nor4_2 _2198_ (.A(net780),
    .B(net785),
    .C(net782),
    .Y(_1618_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1563_));
 sg13g2_nand3_1 _2199_ (.B(_1525_),
    .C(_1562_),
    .A(_1444_),
    .Y(_1619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2200_ (.A(_1581_),
    .B(_1618_),
    .Y(_1620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2201_ (.Y(_1621_),
    .A(_1582_),
    .B(_1619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2202_ (.A(net751),
    .B(_1615_),
    .C(_1617_),
    .D(_1620_),
    .X(_1622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2203_ (.A(_1607_),
    .B(_1622_),
    .X(_1623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2204_ (.Y(_1624_),
    .A(_1607_),
    .B(_1622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2205_ (.X(_1625_),
    .A(_1579_),
    .B(_1607_),
    .C(_1622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2206_ (.Y(_1626_),
    .A(_1579_),
    .B(_1623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2207_ (.A(_1442_),
    .B(net772),
    .Y(_1627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2208_ (.S0(net775),
    .A0(\sap_3_inst.alu.flags[0] ),
    .A1(net762),
    .A2(\sap_3_inst.alu.flags[2] ),
    .A3(\sap_3_inst.alu.flags[3] ),
    .S1(net773),
    .X(_1628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2209_ (.Y(_1629_),
    .A(net778),
    .B(_1628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2210_ (.Y(_1630_),
    .A(net743),
    .B(_1629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2211_ (.A(net759),
    .B_N(\sap_3_inst.controller.stage[3] ),
    .Y(_1631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2212_ (.A(net755),
    .B(net746),
    .X(_1632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2213_ (.Y(_1633_),
    .A(net755),
    .B(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2214_ (.A(_1571_),
    .B(_1632_),
    .Y(_1634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2215_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1630_),
    .A2(_1634_),
    .Y(_1635_),
    .B1(_1619_));
 sg13g2_nand2_1 _2216_ (.Y(_1636_),
    .A(_1573_),
    .B(net730),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2217_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1581_),
    .C1(_1635_),
    .B1(_1636_),
    .A1(_1607_),
    .Y(_1637_),
    .A2(_1622_));
 sg13g2_and2_1 _2218_ (.A(net758),
    .B(net746),
    .X(_1638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2219_ (.Y(_1639_),
    .A(net758),
    .B(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2220_ (.Y(_1640_),
    .A(net732),
    .B(_1630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2221_ (.B1(_1613_),
    .VDD(VPWR),
    .Y(_1641_),
    .VSS(VGND),
    .A1(_1638_),
    .A2(_1640_));
 sg13g2_and2_1 _2222_ (.A(\sap_3_inst.controller.stage[3] ),
    .B(net759),
    .X(_1642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2223_ (.Y(_1643_),
    .A(net759),
    .B(_1507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2224_ (.A(_1507_),
    .B(_1642_),
    .X(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2225_ (.Y(_1645_),
    .A(net760),
    .B(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2226_ (.A(net761),
    .B(_1645_),
    .Y(_1646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2227_ (.Y(_1647_),
    .A(_1534_),
    .B(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2228_ (.Y(_1648_),
    .B1(_1642_),
    .B2(net755),
    .A2(net746),
    .A1(_1534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2229_ (.Y(_1649_),
    .A(net732),
    .B(_1648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2230_ (.A(_1644_),
    .B(_1649_),
    .Y(_1650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2231_ (.A(_1644_),
    .B_N(_1648_),
    .Y(_1651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2232_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1630_),
    .A2(_1650_),
    .Y(_1652_),
    .B1(_1609_));
 sg13g2_a22oi_1 _2233_ (.Y(_1653_),
    .B1(_1639_),
    .B2(_1573_),
    .A2(net753),
    .A1(_1587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2234_ (.Y(_1654_),
    .B1(_1642_),
    .B2(net758),
    .A2(net746),
    .A1(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2235_ (.VDD(VPWR),
    .Y(_1655_),
    .A(_1654_),
    .VSS(VGND));
 sg13g2_and2_1 _2236_ (.A(_1507_),
    .B(net746),
    .X(_1656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2237_ (.Y(_1657_),
    .A(_1507_),
    .B(net746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2238_ (.A(net748),
    .B(_1657_),
    .Y(_1658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2239_ (.A(net734),
    .B(_1603_),
    .Y(_1659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2240_ (.A(net742),
    .B(_1617_),
    .Y(_1660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2241_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1661_),
    .B(_1660_),
    .A(_1659_));
 sg13g2_a21oi_1 _2242_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net732),
    .A2(_1648_),
    .Y(_1662_),
    .B1(net749));
 sg13g2_a21oi_1 _2243_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1573_),
    .A2(_1654_),
    .Y(_1663_),
    .B1(net751));
 sg13g2_a21oi_1 _2244_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1573_),
    .A2(net730),
    .Y(_1664_),
    .B1(_1598_));
 sg13g2_nor2_1 _2245_ (.A(_1658_),
    .B(_1663_),
    .Y(_1665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2246_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1573_),
    .A2(_1651_),
    .Y(_1666_),
    .B1(net749));
 sg13g2_nor4_1 _2247_ (.A(_1653_),
    .B(_1661_),
    .C(_1664_),
    .D(_1666_),
    .Y(_1667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2248_ (.B(_1641_),
    .C(_1665_),
    .A(_1637_),
    .Y(_1668_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1667_));
 sg13g2_o21ai_1 _2249_ (.B1(_1626_),
    .VDD(VPWR),
    .Y(_1669_),
    .VSS(VGND),
    .A1(_1652_),
    .A2(_1668_));
 sg13g2_a21oi_1 _2250_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1567_),
    .A2(_1669_),
    .Y(_1670_),
    .B1(_1556_));
 sg13g2_o21ai_1 _2251_ (.B1(_1539_),
    .VDD(VPWR),
    .Y(_1671_),
    .VSS(VGND),
    .A1(_1544_),
    .A2(_1670_));
 sg13g2_nand2_1 _2252_ (.Y(_1672_),
    .A(net757),
    .B(_1671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2253_ (.Y(_1673_),
    .B1(_1538_),
    .B2(_1672_),
    .A2(_1505_),
    .A1(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2254_ (.VDD(VPWR),
    .Y(_1674_),
    .A(_1673_),
    .VSS(VGND));
 sg13g2_nor2_1 _2255_ (.A(_1444_),
    .B(_1584_),
    .Y(_1675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2256_ (.B(net786),
    .C(net783),
    .A(net781),
    .Y(_1676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2257_ (.A(_1504_),
    .B(_1558_),
    .Y(_1677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2258_ (.Y(_1678_),
    .A(net758),
    .B(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2259_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1676_),
    .A2(net729),
    .Y(_1679_),
    .B1(_1539_));
 sg13g2_a21oi_1 _2260_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net732),
    .A2(_1639_),
    .Y(_1680_),
    .B1(_1581_));
 sg13g2_a21oi_1 _2261_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1582_),
    .A2(_1598_),
    .Y(_1681_),
    .B1(_1634_));
 sg13g2_a21oi_1 _2262_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1603_),
    .A2(net748),
    .Y(_1682_),
    .B1(net727));
 sg13g2_a21oi_1 _2263_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net732),
    .A2(_1654_),
    .Y(_1683_),
    .B1(net751));
 sg13g2_nor4_1 _2264_ (.A(net744),
    .B(_1681_),
    .C(_1682_),
    .D(_1683_),
    .Y(_1684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2265_ (.A(_1508_),
    .B(_1558_),
    .Y(_1685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2266_ (.VDD(VPWR),
    .Y(_1686_),
    .A(_1685_),
    .VSS(VGND));
 sg13g2_a21oi_1 _2267_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1536_),
    .A2(net746),
    .Y(_1687_),
    .B1(net735));
 sg13g2_a22oi_1 _2268_ (.Y(_1688_),
    .B1(_1686_),
    .B2(_1687_),
    .A2(_1604_),
    .A1(net735),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2269_ (.B1(_1688_),
    .VDD(VPWR),
    .Y(_1689_),
    .VSS(VGND),
    .A1(_1604_),
    .A2(_1659_));
 sg13g2_nand2_1 _2270_ (.Y(_1690_),
    .A(_1504_),
    .B(_1642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2271_ (.B(_1645_),
    .C(_1690_),
    .A(net733),
    .Y(_1691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2272_ (.A(net776),
    .B(net751),
    .C(_1648_),
    .Y(_1692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2273_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net750),
    .A2(_1691_),
    .Y(_1693_),
    .B1(_1692_));
 sg13g2_nand3_1 _2274_ (.B(_1689_),
    .C(_1693_),
    .A(_1684_),
    .Y(_1694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2275_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1606_),
    .A2(_1680_),
    .Y(_1695_),
    .B1(_1694_));
 sg13g2_o21ai_1 _2276_ (.B1(_1567_),
    .VDD(VPWR),
    .Y(_1696_),
    .VSS(VGND),
    .A1(_1579_),
    .A2(_1599_));
 sg13g2_nor2_2 _2277_ (.A(net742),
    .B(_1629_),
    .Y(_1697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2278_ (.A(net744),
    .B(_1691_),
    .Y(_1698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2279_ (.A(_1609_),
    .B(_1697_),
    .C(_1698_),
    .Y(_1699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2280_ (.Y(_1700_),
    .A(_1566_),
    .B(_1571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2281_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1553_),
    .C1(_1660_),
    .B1(_1676_),
    .A1(_1566_),
    .Y(_1701_),
    .A2(_1571_));
 sg13g2_a22oi_1 _2282_ (.Y(_1702_),
    .B1(net746),
    .B2(net758),
    .A2(net754),
    .A1(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2283_ (.VDD(VPWR),
    .Y(_1703_),
    .A(net726),
    .VSS(VGND));
 sg13g2_nor2_1 _2284_ (.A(_1575_),
    .B(_1639_),
    .Y(_1704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2285_ (.A(_1575_),
    .B(net726),
    .Y(_1705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2286_ (.Y(_1706_),
    .A(net749),
    .B(_1705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2287_ (.B1(_1701_),
    .VDD(VPWR),
    .Y(_1707_),
    .VSS(VGND),
    .A1(net765),
    .A2(_1706_));
 sg13g2_nor4_1 _2288_ (.A(_1635_),
    .B(_1696_),
    .C(_1699_),
    .D(_1707_),
    .Y(_1708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2289_ (.A(_1641_),
    .B(_1708_),
    .X(_1709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2290_ (.B1(_1709_),
    .VDD(VPWR),
    .Y(_1710_),
    .VSS(VGND),
    .A1(_1607_),
    .A2(_1695_));
 sg13g2_nor2_1 _2291_ (.A(_1584_),
    .B(_1591_),
    .Y(_1711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2292_ (.B1(_1515_),
    .VDD(VPWR),
    .Y(_1712_),
    .VSS(VGND),
    .A1(_1584_),
    .A2(_1591_));
 sg13g2_nor2b_2 _2293_ (.A(_1712_),
    .B_N(_1541_),
    .Y(_1713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2294_ (.Y(_1714_),
    .B(_1541_),
    .A_N(_1712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2295_ (.A(_1441_),
    .B(net763),
    .Y(_1715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2296_ (.Y(_1716_),
    .A(net778),
    .B(_1518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2297_ (.A(net741),
    .B(_1715_),
    .Y(_1717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2298_ (.Y(_1718_),
    .B(_1556_),
    .A_N(_1717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2299_ (.X(_1719_),
    .A(_1710_),
    .B(_1713_),
    .C(_1718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2300_ (.A(net741),
    .B(_1515_),
    .C(_1675_),
    .Y(_1720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2301_ (.A(_1544_),
    .B(_1719_),
    .C(_1720_),
    .Y(_1721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2302_ (.B1(net757),
    .VDD(VPWR),
    .Y(_1722_),
    .VSS(VGND),
    .A1(_1679_),
    .A2(_1721_));
 sg13g2_nand3_1 _2303_ (.B(_1673_),
    .C(_1722_),
    .A(_1538_),
    .Y(_1723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2304_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1724_),
    .B(_1612_),
    .A(_1608_));
 sg13g2_inv_1 _2305_ (.VDD(VPWR),
    .Y(_1725_),
    .A(_1724_),
    .VSS(VGND));
 sg13g2_nand2_1 _2306_ (.Y(_1726_),
    .A(_1640_),
    .B(_1724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2307_ (.B(_1598_),
    .C(net749),
    .A(_1589_),
    .Y(_1727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2308_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1600_),
    .A2(_1609_),
    .Y(_1728_),
    .B1(_1648_));
 sg13g2_nand2_1 _2309_ (.Y(_1729_),
    .A(_1534_),
    .B(_1642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2310_ (.A(_1610_),
    .B(_1657_),
    .Y(_1730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2311_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1657_),
    .A2(_1729_),
    .Y(_1731_),
    .B1(_1610_));
 sg13g2_a21oi_1 _2312_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1639_),
    .A2(net727),
    .Y(_1732_),
    .B1(net748));
 sg13g2_o21ai_1 _2313_ (.B1(_1574_),
    .VDD(VPWR),
    .Y(_1733_),
    .VSS(VGND),
    .A1(net752),
    .A2(_1727_));
 sg13g2_a21o_1 _2314_ (.A2(_1732_),
    .A1(net765),
    .B1(_1660_),
    .X(_1734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2315_ (.A(_1728_),
    .B(_1731_),
    .C(_1734_),
    .Y(_1735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2316_ (.A(_1624_),
    .B(_1726_),
    .C(_1733_),
    .D(_1735_),
    .X(_1736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2317_ (.Y(_1737_),
    .B1(net743),
    .B2(_1565_),
    .A2(_1505_),
    .A1(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2318_ (.B1(_1737_),
    .VDD(VPWR),
    .Y(_1738_),
    .VSS(VGND),
    .A1(_1625_),
    .A2(_1736_));
 sg13g2_inv_2 _2319_ (.Y(_1739_),
    .A(_1738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2320_ (.Y(_1740_),
    .A(net781),
    .B(_1584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2321_ (.B1(net725),
    .VDD(VPWR),
    .Y(_1741_),
    .VSS(VGND),
    .A1(net740),
    .A2(_1740_));
 sg13g2_nand2_1 _2322_ (.Y(_1742_),
    .A(net743),
    .B(_1604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2323_ (.B1(_1742_),
    .VDD(VPWR),
    .Y(_1743_),
    .VSS(VGND),
    .A1(_1554_),
    .A2(_1740_));
 sg13g2_nand2_1 _2324_ (.Y(_1744_),
    .A(net734),
    .B(net733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2325_ (.A(_1566_),
    .B(_1744_),
    .X(_1745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2326_ (.B1(net773),
    .VDD(VPWR),
    .Y(_1746_),
    .VSS(VGND),
    .A1(_1441_),
    .A2(_1442_));
 sg13g2_nor2_1 _2327_ (.A(net740),
    .B(_1746_),
    .Y(_1747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2328_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1593_),
    .A2(_1638_),
    .Y(_1748_),
    .B1(_1576_));
 sg13g2_nor3_1 _2329_ (.A(_1581_),
    .B(_1597_),
    .C(_1618_),
    .Y(_1749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2330_ (.A(net730),
    .B(_1749_),
    .Y(_1750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2331_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net752),
    .C1(_1659_),
    .B1(_1655_),
    .A1(_1611_),
    .Y(_1751_),
    .A2(_1644_));
 sg13g2_nor2_1 _2332_ (.A(_1692_),
    .B(net725),
    .Y(_1752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2333_ (.B(net753),
    .C(_1614_),
    .A(_1587_),
    .Y(_1753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2334_ (.Y(_1754_),
    .A(_1638_),
    .B(_1753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2335_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1657_),
    .C1(net748),
    .B1(_1748_),
    .A1(_1594_),
    .Y(_1755_),
    .A2(net728));
 sg13g2_or4_1 _2336_ (.A(_1743_),
    .B(_1745_),
    .C(_1750_),
    .D(_1755_),
    .X(_1756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2337_ (.Y(_1757_),
    .B1(_1747_),
    .B2(net736),
    .A2(_1705_),
    .A1(_1593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2338_ (.B(_1752_),
    .C(_1754_),
    .A(_1751_),
    .Y(_1758_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1757_));
 sg13g2_o21ai_1 _2339_ (.B1(_1741_),
    .VDD(VPWR),
    .Y(_1759_),
    .VSS(VGND),
    .A1(_1756_),
    .A2(_1758_));
 sg13g2_nor2_1 _2340_ (.A(net727),
    .B(_1740_),
    .Y(_1760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2341_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1761_),
    .B(_1760_),
    .A(_1539_));
 sg13g2_nand2_2 _2342_ (.Y(_1762_),
    .A(_1505_),
    .B(_1508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2343_ (.B(_1761_),
    .C(_1762_),
    .A(_1530_),
    .Y(_1763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2344_ (.B1(_1762_),
    .VDD(VPWR),
    .Y(_1764_),
    .VSS(VGND),
    .A1(net766),
    .A2(_1521_));
 sg13g2_a21oi_2 _2345_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1763_),
    .Y(_1765_),
    .A2(_1759_),
    .A1(net756));
 sg13g2_inv_2 _2346_ (.Y(_1766_),
    .A(_1765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2347_ (.Y(_1767_),
    .A(_1627_),
    .B(_1705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2348_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1604_),
    .C1(_1728_),
    .B1(_1656_),
    .A1(_1597_),
    .Y(_1768_),
    .A2(_1632_));
 sg13g2_a21oi_1 _2349_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net740),
    .A2(net727),
    .Y(_1769_),
    .B1(_1603_));
 sg13g2_o21ai_1 _2350_ (.B1(_1602_),
    .VDD(VPWR),
    .Y(_1770_),
    .VSS(VGND),
    .A1(net745),
    .A2(net728));
 sg13g2_o21ai_1 _2351_ (.B1(net775),
    .VDD(VPWR),
    .Y(_1771_),
    .VSS(VGND),
    .A1(_1732_),
    .A2(_1769_));
 sg13g2_and4_1 _2352_ (.A(_1751_),
    .B(_1754_),
    .C(_1768_),
    .D(_1771_),
    .X(_1772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2353_ (.Y(_1773_),
    .B1(_1772_),
    .B2(_1637_),
    .A2(_1767_),
    .A1(_1625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2354_ (.B(net736),
    .C(_1717_),
    .A(net774),
    .Y(_1774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2355_ (.B(_1553_),
    .C(_1676_),
    .A(net783),
    .Y(_1775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2356_ (.B(_1774_),
    .C(_1775_),
    .A(_1700_),
    .Y(_1776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2357_ (.A(_1555_),
    .B(net725),
    .Y(_1777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2358_ (.B1(_1777_),
    .VDD(VPWR),
    .Y(_1778_),
    .VSS(VGND),
    .A1(_1773_),
    .A2(_1776_));
 sg13g2_a21oi_1 _2359_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net783),
    .A2(_1720_),
    .Y(_1779_),
    .B1(_1520_));
 sg13g2_nand3_1 _2360_ (.B(_1676_),
    .C(net729),
    .A(net783),
    .Y(_1780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2361_ (.Y(_1781_),
    .A(_1520_),
    .B(_1780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2362_ (.B(_1762_),
    .C(_1781_),
    .A(net757),
    .Y(_1782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2363_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1782_),
    .Y(_1783_),
    .A2(_1779_),
    .A1(_1778_));
 sg13g2_a21o_2 _2364_ (.A2(_1779_),
    .A1(_1778_),
    .B1(_1782_),
    .X(_1784_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2365_ (.B(_1623_),
    .C(_1704_),
    .A(net764),
    .Y(_1785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2366_ (.A(_1524_),
    .B(_1676_),
    .Y(_1786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2367_ (.A(_1546_),
    .B(_1565_),
    .C(_1566_),
    .Y(_1787_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1786_));
 sg13g2_nand2_1 _2368_ (.Y(_1788_),
    .A(_1515_),
    .B(_1787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2369_ (.B(net743),
    .C(_1676_),
    .A(net786),
    .Y(_1789_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1788_));
 sg13g2_nand4_1 _2370_ (.B(net745),
    .C(net763),
    .A(net777),
    .Y(_1790_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1549_));
 sg13g2_nand3_1 _2371_ (.B(_1742_),
    .C(_1790_),
    .A(net756),
    .Y(_1791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2372_ (.B(net752),
    .C(_1642_),
    .A(net755),
    .Y(_1792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2373_ (.A(net776),
    .B(_1792_),
    .Y(_1793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2374_ (.A(_1682_),
    .B(net723),
    .C(_1791_),
    .D(_1793_),
    .Y(_1794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2375_ (.B(_1789_),
    .C(_1794_),
    .A(_1785_),
    .Y(_1795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2376_ (.B(_1503_),
    .C(_1557_),
    .A(net786),
    .Y(_1796_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1676_));
 sg13g2_nand2_1 _2377_ (.Y(_1797_),
    .A(_1520_),
    .B(_1796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2378_ (.A(_1795_),
    .B(_1797_),
    .X(_1798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2379_ (.Y(_1799_),
    .A(_1795_),
    .B(_1797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2380_ (.A(_1738_),
    .B(_1765_),
    .C(_1783_),
    .Y(_1800_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1798_));
 sg13g2_nand4_1 _2381_ (.B(_1766_),
    .C(_1784_),
    .A(_1739_),
    .Y(_1801_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1799_));
 sg13g2_nor3_2 _2382_ (.A(_1739_),
    .B(_1784_),
    .C(_1798_),
    .Y(_1802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2383_ (.A(_1738_),
    .B(_1765_),
    .C(_1784_),
    .Y(_1803_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1799_));
 sg13g2_nor3_2 _2384_ (.A(_1739_),
    .B(_1784_),
    .C(_1799_),
    .Y(_1804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2385_ (.VDD(VPWR),
    .Y(_1805_),
    .A(net642),
    .VSS(VGND));
 sg13g2_nor3_2 _2386_ (.A(_1766_),
    .B(_1783_),
    .C(_1798_),
    .Y(_1806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2387_ (.A(_1766_),
    .B(_1784_),
    .C(_1798_),
    .Y(_1807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2388_ (.A(_1766_),
    .B(_1783_),
    .C(_1799_),
    .Y(_1808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2389_ (.A(_1739_),
    .B(_1783_),
    .C(_1798_),
    .Y(_1809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2390_ (.Y(_1810_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .A2(net637),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2391_ (.A(_1738_),
    .B(_1765_),
    .C(_1784_),
    .Y(_1811_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1798_));
 sg13g2_nor4_2 _2392_ (.A(_1738_),
    .B(_1765_),
    .C(_1783_),
    .Y(_1812_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1799_));
 sg13g2_a22oi_1 _2393_ (.Y(_1813_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .A2(net647),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2394_ (.Y(_1814_),
    .B1(net642),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .A2(_1730_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2395_ (.A(_1810_),
    .B(_1814_),
    .X(_1815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2396_ (.Y(_1816_),
    .B1(net638),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .A2(net640),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2397_ (.Y(_1817_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .A2(net645),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2398_ (.A(net648),
    .B(_1813_),
    .C(_1816_),
    .D(_1817_),
    .X(_1818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2399_ (.Y(_1819_),
    .B1(_1815_),
    .B2(_1818_),
    .A2(net650),
    .A1(_1494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2400_ (.A(_1723_),
    .B_N(_1819_),
    .Y(_1820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2401_ (.A(net756),
    .B(_1678_),
    .Y(_1821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2402_ (.Y(_1822_),
    .A(_1520_),
    .B(net728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2403_ (.A(_1550_),
    .B(net734),
    .Y(_1823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2404_ (.VDD(VPWR),
    .Y(_1824_),
    .A(_1823_),
    .VSS(VGND));
 sg13g2_a22oi_1 _2405_ (.Y(_1825_),
    .B1(_1685_),
    .B2(_1602_),
    .A2(_1646_),
    .A1(_1597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2406_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1826_),
    .B(_1825_),
    .A(net777));
 sg13g2_nor2_1 _2407_ (.A(net748),
    .B(_1647_),
    .Y(_1827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2408_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net733),
    .A2(_1647_),
    .Y(_1828_),
    .B1(_1605_));
 sg13g2_nor3_1 _2409_ (.A(net763),
    .B(_1560_),
    .C(_1575_),
    .Y(_1829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2410_ (.A(net737),
    .B(_1828_),
    .C(_1829_),
    .Y(_1830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2411_ (.Y(_1831_),
    .A(_1826_),
    .B(_1830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2412_ (.B1(_1831_),
    .VDD(VPWR),
    .Y(_1832_),
    .VSS(VGND),
    .A1(_1551_),
    .A2(_1823_));
 sg13g2_nor2_1 _2413_ (.A(net740),
    .B(_1676_),
    .Y(_1833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2414_ (.B1(net724),
    .VDD(VPWR),
    .Y(_1834_),
    .VSS(VGND),
    .A1(_1543_),
    .A2(net732));
 sg13g2_a21oi_1 _2415_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1514_),
    .A2(_1833_),
    .Y(_1835_),
    .B1(_1834_));
 sg13g2_a21oi_1 _2416_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1713_),
    .A2(_1832_),
    .Y(_1836_),
    .B1(_1835_));
 sg13g2_a22oi_1 _2417_ (.Y(_1837_),
    .B1(_1836_),
    .B2(net756),
    .A2(_1821_),
    .A1(_1675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2418_ (.A(net789),
    .B(net628),
    .Y(_1838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2419_ (.A(net763),
    .B(_1575_),
    .C(_1639_),
    .Y(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2420_ (.Y(_1840_),
    .A(\sap_3_inst.alu.flags[7] ),
    .B(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2421_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net628),
    .A2(_1840_),
    .Y(_1841_),
    .B1(_1838_));
 sg13g2_o21ai_1 _2422_ (.B1(_1530_),
    .VDD(VPWR),
    .Y(_1842_),
    .VSS(VGND),
    .A1(_1517_),
    .A2(net729));
 sg13g2_nand3_1 _2423_ (.B(_1597_),
    .C(_1646_),
    .A(net777),
    .Y(_1843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2424_ (.Y(_1844_),
    .A(net731),
    .B(_1843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2425_ (.B1(_1844_),
    .VDD(VPWR),
    .Y(_1845_),
    .VSS(VGND),
    .A1(_1724_),
    .A2(_1727_));
 sg13g2_o21ai_1 _2426_ (.B1(net731),
    .VDD(VPWR),
    .Y(_1846_),
    .VSS(VGND),
    .A1(_1441_),
    .A2(_1648_));
 sg13g2_and2_1 _2427_ (.A(net752),
    .B(_1846_),
    .X(_1847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2428_ (.B(_1602_),
    .C(_1685_),
    .A(net777),
    .Y(_1848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2429_ (.Y(_1849_),
    .A(_1565_),
    .B(net728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2430_ (.Y(_1850_),
    .A(_1569_),
    .B(_1576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2431_ (.A(_1504_),
    .B(net766),
    .C(_1524_),
    .D(_1558_),
    .Y(_1851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2432_ (.A(net737),
    .B(_1851_),
    .Y(_1852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2433_ (.B(_1849_),
    .C(_1850_),
    .A(_1848_),
    .Y(_1853_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1852_));
 sg13g2_nor2_1 _2434_ (.A(_1847_),
    .B(_1853_),
    .Y(_1854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2435_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1854_),
    .C1(net724),
    .B1(_1845_),
    .A1(net737),
    .Y(_1855_),
    .A2(_1780_));
 sg13g2_nor2_1 _2436_ (.A(_1541_),
    .B(_1678_),
    .Y(_1856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2437_ (.A(_1516_),
    .B(_1855_),
    .C(_1856_),
    .Y(_1857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2438_ (.B1(_1533_),
    .VDD(VPWR),
    .Y(_1858_),
    .VSS(VGND),
    .A1(_1842_),
    .A2(_1857_));
 sg13g2_and2_1 _2439_ (.A(net8),
    .B(_1858_),
    .X(_1859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2440_ (.Y(_1860_),
    .B1(_1809_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ),
    .A2(net637),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2441_ (.Y(_1861_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .A2(net645),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2442_ (.Y(_1862_),
    .B1(net647),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .A2(_1730_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2443_ (.Y(_1863_),
    .B1(_1807_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .A2(net650),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2444_ (.B(_1861_),
    .C(_1862_),
    .A(_1860_),
    .Y(_1864_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1863_));
 sg13g2_a221oi_1 _2445_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .C1(_1864_),
    .B1(_1811_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .Y(_1865_),
    .A2(_1806_));
 sg13g2_a21oi_1 _2446_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1805_),
    .A2(_1865_),
    .Y(_1866_),
    .B1(_1673_));
 sg13g2_or4_1 _2447_ (.A(_1820_),
    .B(_1841_),
    .C(_1859_),
    .D(_1866_),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2448_ (.A(net763),
    .B(_1570_),
    .C(_1678_),
    .Y(_1867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2449_ (.B(_1569_),
    .C(net728),
    .A(net765),
    .Y(_1868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2450_ (.A0(\sap_3_inst.alu.flags[7] ),
    .A1(net34),
    .S(_1867_),
    .X(_0032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2451_ (.Y(_1869_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .A2(net645),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2452_ (.Y(_1870_),
    .B1(net640),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .A2(net643),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2453_ (.Y(_1871_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .A2(net722),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2454_ (.Y(_1872_),
    .B1(net637),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .A2(net647),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2455_ (.Y(_1873_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .A2(net638),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2456_ (.A(_1872_),
    .B(_1873_),
    .X(_1874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2457_ (.A(net648),
    .B(_1869_),
    .C(_1870_),
    .D(_1871_),
    .X(_1875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2458_ (.Y(_1876_),
    .B1(_1874_),
    .B2(_1875_),
    .A2(net650),
    .A1(_1484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2459_ (.Y(_1877_),
    .B(_1876_),
    .A_N(_1723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2460_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1878_),
    .B(net629),
    .A(net792));
 sg13g2_nand2_1 _2461_ (.Y(_1879_),
    .A(\sap_3_inst.alu.flags[6] ),
    .B(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2462_ (.Y(_1880_),
    .A(net628),
    .B(_1879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2463_ (.Y(_1881_),
    .B1(_1878_),
    .B2(_1880_),
    .A2(_1858_),
    .A1(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2464_ (.Y(_1882_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ),
    .A2(net650),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2465_ (.Y(_1883_),
    .B1(net637),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .A2(net638),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2466_ (.Y(_1884_),
    .A(_1882_),
    .B(_1883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2467_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .C1(net643),
    .B1(net647),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ),
    .Y(_1885_),
    .A2(net722));
 sg13g2_a22oi_1 _2468_ (.Y(_1886_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .A2(net632),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2469_ (.Y(_1887_),
    .B1(net640),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .A2(net645),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2470_ (.B(_1886_),
    .C(_1887_),
    .A(_1885_),
    .Y(_1888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2471_ (.B1(net576),
    .VDD(VPWR),
    .Y(_1889_),
    .VSS(VGND),
    .A1(_1884_),
    .A2(_1888_));
 sg13g2_nand3_1 _2472_ (.B(_1881_),
    .C(_1889_),
    .A(_1877_),
    .Y(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2473_ (.A0(\sap_3_inst.alu.flags[6] ),
    .A1(net33),
    .S(_1867_),
    .X(_0031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2474_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[0][5] ),
    .B(_1801_),
    .Y(_1890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2475_ (.Y(_1891_),
    .B1(net640),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .A2(net643),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2476_ (.Y(_1892_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .A2(net645),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2477_ (.Y(_1893_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .A2(net647),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2478_ (.Y(_1894_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .A2(net722),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2479_ (.Y(_1895_),
    .A(_1893_),
    .B(_1894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2480_ (.Y(_1896_),
    .B1(net637),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .A2(net638),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2481_ (.B(_1891_),
    .C(_1892_),
    .A(net648),
    .Y(_1897_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1896_));
 sg13g2_nor2_1 _2482_ (.A(_1895_),
    .B(_1897_),
    .Y(_1898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2483_ (.A(_1890_),
    .B(_1898_),
    .Y(_1899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2484_ (.A(_1723_),
    .B(_1890_),
    .C(_1898_),
    .Y(_1900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2485_ (.A(net795),
    .B(net628),
    .Y(_1901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2486_ (.Y(_1902_),
    .A(\sap_3_inst.alu.flags[5] ),
    .B(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2487_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net629),
    .A2(_1902_),
    .Y(_1903_),
    .B1(_1901_));
 sg13g2_a22oi_1 _2488_ (.Y(_1904_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .A2(net650),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2489_ (.Y(_1905_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .A2(net645),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2490_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ),
    .C1(net643),
    .B1(net638),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .Y(_1906_),
    .A2(net722));
 sg13g2_a22oi_1 _2491_ (.Y(_1907_),
    .B1(net640),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .A2(net647),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2492_ (.Y(_1908_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .A2(net637),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2493_ (.X(_1909_),
    .A(_1906_),
    .B(_1907_),
    .C(_1908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2494_ (.B(_1905_),
    .C(_1909_),
    .A(_1904_),
    .Y(_1910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2495_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net576),
    .C1(_1903_),
    .B1(_1910_),
    .A1(net6),
    .Y(_1911_),
    .A2(_1858_));
 sg13g2_nand2b_2 _2496_ (.Y(net573),
    .B(_1911_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1900_));
 sg13g2_mux2_1 _2497_ (.A0(\sap_3_inst.alu.flags[5] ),
    .A1(net573),
    .S(_1867_),
    .X(_0030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2498_ (.Y(_1912_),
    .B1(net635),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .A2(net642),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2499_ (.Y(_1913_),
    .B1(net639),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2500_ (.Y(_1914_),
    .B1(net630),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .A2(net644),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2501_ (.A(_1912_),
    .B(_1914_),
    .X(_1915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2502_ (.Y(_1916_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .A2(net636),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2503_ (.Y(_1917_),
    .B1(net646),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ),
    .A2(net722),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2504_ (.A(net648),
    .B(_1913_),
    .C(_1916_),
    .D(_1917_),
    .X(_1918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2505_ (.Y(_1919_),
    .B1(_1915_),
    .B2(_1918_),
    .A2(net649),
    .A1(_1474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2506_ (.Y(_1920_),
    .B(_1919_),
    .A_N(_1723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2507_ (.Y(_1921_),
    .A(net5),
    .B(_1858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2508_ (.Y(_1922_),
    .A(\sap_3_inst.alu.flags[4] ),
    .B(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2509_ (.Y(_1923_),
    .A(net628),
    .B(_1922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2510_ (.B1(_1923_),
    .VDD(VPWR),
    .Y(_1924_),
    .VSS(VGND),
    .A1(net797),
    .A2(net628));
 sg13g2_a22oi_1 _2511_ (.Y(_1925_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .A2(net640),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2512_ (.Y(_1926_),
    .B1(net638),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .A2(net646),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2513_ (.Y(_1927_),
    .A(_1925_),
    .B(_1926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2514_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .C1(net642),
    .B1(net633),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ),
    .Y(_1928_),
    .A2(net722));
 sg13g2_a22oi_1 _2515_ (.Y(_1929_),
    .B1(net636),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .A2(net644),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2516_ (.Y(_1930_),
    .B1(net630),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .A2(net649),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2517_ (.B(_1929_),
    .C(_1930_),
    .A(_1928_),
    .Y(_1931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2518_ (.B1(net576),
    .VDD(VPWR),
    .Y(_1932_),
    .VSS(VGND),
    .A1(_1927_),
    .A2(_1931_));
 sg13g2_nand4_1 _2519_ (.B(_1921_),
    .C(_1924_),
    .A(_1920_),
    .Y(net21),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1932_));
 sg13g2_mux2_1 _2520_ (.A0(\sap_3_inst.alu.flags[4] ),
    .A1(net32),
    .S(_1867_),
    .X(_0029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2521_ (.B1(net724),
    .VDD(VPWR),
    .Y(_1933_),
    .VSS(VGND),
    .A1(_1543_),
    .A2(net734));
 sg13g2_a22oi_1 _2522_ (.Y(_1934_),
    .B1(net729),
    .B2(net769),
    .A2(_1675_),
    .A1(net745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2523_ (.A(net771),
    .B(_1934_),
    .Y(_1935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2524_ (.Y(_1936_),
    .A(net735),
    .B(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2525_ (.Y(_1937_),
    .B1(_1936_),
    .B2(net748),
    .A2(_1633_),
    .A1(net734),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2526_ (.A(net724),
    .B(_1935_),
    .C(_1937_),
    .Y(_1938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2527_ (.A(net741),
    .B(_1550_),
    .C(_1716_),
    .Y(_1939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2528_ (.A(net724),
    .B(_1939_),
    .Y(_1940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2529_ (.B1(_1940_),
    .VDD(VPWR),
    .Y(_1941_),
    .VSS(VGND),
    .A1(_1550_),
    .A2(net727));
 sg13g2_nand2_1 _2530_ (.Y(_1942_),
    .A(_1548_),
    .B(net735),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2531_ (.B1(_1942_),
    .VDD(VPWR),
    .Y(_1943_),
    .VSS(VGND),
    .A1(net737),
    .A2(_1938_));
 sg13g2_and2_1 _2532_ (.A(_1933_),
    .B(_1941_),
    .X(_1944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2533_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net714),
    .Y(_1945_),
    .A2(_1943_),
    .A1(_1933_));
 sg13g2_nand2_2 _2534_ (.Y(_1946_),
    .A(_1868_),
    .B(_1945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2535_ (.A(net745),
    .B(_1786_),
    .X(_1947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2536_ (.Y(_1948_),
    .B1(_1935_),
    .B2(_1551_),
    .A2(_1559_),
    .A1(_1545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2537_ (.A(_1948_),
    .B_N(net773),
    .Y(_1949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2538_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1950_),
    .B(_1949_),
    .A(_1947_));
 sg13g2_nand2b_2 _2539_ (.Y(_1951_),
    .B(_1949_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1947_));
 sg13g2_nor2_1 _2540_ (.A(_1441_),
    .B(_1948_),
    .Y(_1952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2541_ (.A(_1550_),
    .B(_1796_),
    .Y(_1953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2542_ (.A(net748),
    .B(_1633_),
    .Y(_1954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2543_ (.A(_1952_),
    .B(net721),
    .C(_1954_),
    .Y(_1955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2544_ (.A(_1952_),
    .B(net721),
    .C(_1954_),
    .X(_1956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2545_ (.A(_1442_),
    .B(_1948_),
    .Y(_1957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2546_ (.Y(_1958_),
    .A(_1956_),
    .B(_1957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2547_ (.Y(_1959_),
    .B(_1958_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1951_));
 sg13g2_nand2_2 _2548_ (.Y(_1960_),
    .A(_1950_),
    .B(_1959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2549_ (.Y(_1961_),
    .A(_1946_),
    .B(_1960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2550_ (.Y(_1962_),
    .A(\sap_3_inst.alu.flags[3] ),
    .B(_1961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2551_ (.Y(_1963_),
    .B1(net644),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .A2(net646),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2552_ (.Y(_1964_),
    .B1(net630),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .A2(net639),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2553_ (.Y(_1965_),
    .B1(net642),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .A2(net723),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2554_ (.A(_1963_),
    .B(_1965_),
    .X(_1966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2555_ (.Y(_1967_),
    .B1(net636),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2556_ (.Y(_1968_),
    .B1(net633),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ),
    .A2(net635),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2557_ (.A(net648),
    .B(_1964_),
    .C(_1967_),
    .D(_1968_),
    .X(_1969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2558_ (.Y(_1970_),
    .B1(_1966_),
    .B2(_1969_),
    .A2(net649),
    .A1(_1446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2559_ (.Y(_1971_),
    .B(_1970_),
    .A_N(_1723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2560_ (.Y(_1972_),
    .B1(_1858_),
    .B2(net4),
    .A2(_1839_),
    .A1(\sap_3_inst.alu.flags[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2561_ (.B1(_1972_),
    .VDD(VPWR),
    .Y(_1973_),
    .VSS(VGND),
    .A1(_1445_),
    .A2(net629));
 sg13g2_a22oi_1 _2562_ (.Y(_1974_),
    .B1(net646),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .A2(net649),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2563_ (.Y(_1975_),
    .B1(net633),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .A2(net723),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2564_ (.Y(_1976_),
    .B1(net639),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2565_ (.Y(_1977_),
    .B1(net630),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ),
    .A2(net636),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2566_ (.Y(_1978_),
    .B1(net635),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .A2(net644),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2567_ (.A(_1805_),
    .B(_1974_),
    .C(_1975_),
    .D(_1978_),
    .X(_1979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2568_ (.B(_1977_),
    .C(_1979_),
    .A(_1976_),
    .Y(_1980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2569_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_1980_),
    .Y(_1981_),
    .B1(_1973_));
 sg13g2_and2_1 _2570_ (.A(_1971_),
    .B(_1981_),
    .X(_1982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2571_ (.Y(net20),
    .A(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2572_ (.Y(_1983_),
    .A(_1867_),
    .B(_1982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2573_ (.B1(_1983_),
    .VDD(VPWR),
    .Y(_1984_),
    .VSS(VGND),
    .A1(net789),
    .A2(_1867_));
 sg13g2_o21ai_1 _2574_ (.B1(_1962_),
    .VDD(VPWR),
    .Y(_0028_),
    .VSS(VGND),
    .A1(_1961_),
    .A2(_1984_));
 sg13g2_nand2_1 _2575_ (.Y(_1985_),
    .A(\sap_3_inst.alu.flags[2] ),
    .B(_1961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2576_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[0][2] ),
    .B(net648),
    .Y(_1986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2577_ (.Y(_1987_),
    .B1(net633),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .A2(net635),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2578_ (.Y(_1988_),
    .B1(net630),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .A2(net639),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2579_ (.A(_1987_),
    .B(_1988_),
    .X(_1989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2580_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ),
    .C1(net649),
    .B1(net644),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ),
    .Y(_1990_),
    .A2(net723));
 sg13g2_a22oi_1 _2581_ (.Y(_1991_),
    .B1(net636),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2582_ (.Y(_1992_),
    .B1(net642),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .A2(net646),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2583_ (.X(_1993_),
    .A(_1990_),
    .B(_1991_),
    .C(_1992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _2584_ (.A2(_1993_),
    .A1(_1989_),
    .B1(_1986_),
    .X(_1994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2585_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1995_),
    .B(_1994_),
    .A(_1723_));
 sg13g2_or2_1 _2586_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1996_),
    .B(net628),
    .A(net802));
 sg13g2_nand2_1 _2587_ (.Y(_1997_),
    .A(\sap_3_inst.alu.flags[2] ),
    .B(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2588_ (.Y(_1998_),
    .A(net629),
    .B(_1997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2589_ (.Y(_1999_),
    .B1(_1996_),
    .B2(_1998_),
    .A2(_1858_),
    .A1(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2590_ (.Y(_2000_),
    .B1(net633),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2591_ (.Y(_2001_),
    .B1(net635),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ),
    .A2(net649),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2592_ (.Y(_2002_),
    .B1(net636),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .A2(net646),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2593_ (.Y(_2003_),
    .B1(net630),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .A2(net639),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2594_ (.Y(_2004_),
    .A(_2002_),
    .B(_2003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2595_ (.Y(_2005_),
    .B1(net644),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .A2(net723),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2596_ (.B(_2000_),
    .C(_2001_),
    .A(_1805_),
    .Y(_2006_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2005_));
 sg13g2_o21ai_1 _2597_ (.B1(net577),
    .VDD(VPWR),
    .Y(_2007_),
    .VSS(VGND),
    .A1(_2004_),
    .A2(_2006_));
 sg13g2_nand3_1 _2598_ (.B(_1999_),
    .C(_2007_),
    .A(_1995_),
    .Y(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2599_ (.VDD(VPWR),
    .Y(_2008_),
    .A(net19),
    .VSS(VGND));
 sg13g2_xnor2_1 _2600_ (.Y(_2009_),
    .A(net789),
    .B(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2601_ (.B(net797),
    .A(net795),
    .X(_2010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2602_ (.Y(_2011_),
    .A(_2009_),
    .B(_2010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2603_ (.B(net805),
    .A(net803),
    .X(_2012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2604_ (.B(net801),
    .A(net800),
    .X(_2013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2605_ (.Y(_2014_),
    .A(_2012_),
    .B(_2013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2606_ (.Y(_0196_),
    .A(_2011_),
    .B(_2014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2607_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1868_),
    .A2(_0196_),
    .Y(_0197_),
    .B1(_1961_));
 sg13g2_o21ai_1 _2608_ (.B1(_0197_),
    .VDD(VPWR),
    .Y(_0198_),
    .VSS(VGND),
    .A1(_1868_),
    .A2(net19));
 sg13g2_nand2_1 _2609_ (.Y(_0027_),
    .A(_1985_),
    .B(_0198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2610_ (.Y(_0199_),
    .B(_1947_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1949_));
 sg13g2_nand2_1 _2611_ (.Y(_0200_),
    .A(_1959_),
    .B(_0199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2612_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0201_),
    .B(_1950_),
    .A(net714));
 sg13g2_nand2_1 _2613_ (.Y(_0202_),
    .A(net775),
    .B(_1947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2614_ (.B(_0199_),
    .C(_0201_),
    .A(_1959_),
    .Y(_0203_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0202_));
 sg13g2_nand2_1 _2615_ (.Y(_0204_),
    .A(_1946_),
    .B(_0203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2616_ (.Y(_0205_),
    .A(net762),
    .B(_0204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2617_ (.Y(_0206_),
    .B1(net641),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .A2(net644),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2618_ (.Y(_0207_),
    .B1(net635),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .A2(net646),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2619_ (.A(_0206_),
    .B(_0207_),
    .X(_0208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2620_ (.Y(_0209_),
    .B1(net630),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .A2(net639),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2621_ (.Y(_0210_),
    .B1(net636),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .A2(net642),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2622_ (.Y(_0211_),
    .B1(net633),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .A2(net723),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2623_ (.A(net648),
    .B(_0209_),
    .C(_0210_),
    .D(_0211_),
    .X(_0212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2624_ (.Y(_0213_),
    .B1(_0208_),
    .B2(_0212_),
    .A2(net649),
    .A1(_1461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2625_ (.Y(_0214_),
    .B(_0213_),
    .A_N(_1723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2626_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0215_),
    .B(net629),
    .A(net803));
 sg13g2_nand2_1 _2627_ (.Y(_0216_),
    .A(net762),
    .B(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2628_ (.Y(_0217_),
    .A(net629),
    .B(_0216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2629_ (.Y(_0218_),
    .B1(_0215_),
    .B2(_0217_),
    .A2(_1858_),
    .A1(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2630_ (.Y(_0219_),
    .B1(net633),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .A2(net635),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2631_ (.Y(_0220_),
    .B1(net630),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .A2(net644),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2632_ (.Y(_0221_),
    .A(_0219_),
    .B(_0220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2633_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .C1(net642),
    .B1(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ),
    .Y(_0222_),
    .A2(net723));
 sg13g2_a22oi_1 _2634_ (.Y(_0223_),
    .B1(net636),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .A2(net639),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2635_ (.Y(_0224_),
    .B1(net646),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .A2(net649),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2636_ (.B(_0223_),
    .C(_0224_),
    .A(_0222_),
    .Y(_0225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2637_ (.B1(net576),
    .VDD(VPWR),
    .Y(_0226_),
    .VSS(VGND),
    .A1(_0221_),
    .A2(_0225_));
 sg13g2_nand3_1 _2638_ (.B(_0218_),
    .C(_0226_),
    .A(_0214_),
    .Y(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2639_ (.A(net18),
    .Y(_0227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2640_ (.A(\sap_3_inst.alu.carry ),
    .B(_1867_),
    .Y(_0228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2641_ (.A2(_0227_),
    .A1(_1867_),
    .B1(_0204_),
    .X(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2642_ (.B1(_0205_),
    .VDD(VPWR),
    .Y(_0026_),
    .VSS(VGND),
    .A1(_0228_),
    .A2(_0229_));
 sg13g2_nand2b_1 _2643_ (.Y(_0230_),
    .B(_1946_),
    .A_N(_1786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2644_ (.Y(_0231_),
    .A(\sap_3_inst.alu.flags[0] ),
    .B(_0230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2645_ (.Y(_0232_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .A2(net643),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2646_ (.Y(_0233_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .A2(net638),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2647_ (.Y(_0234_),
    .B1(net637),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .A2(net722),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2648_ (.A(_0233_),
    .B(_0234_),
    .X(_0235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2649_ (.Y(_0236_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .A2(net647),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2650_ (.B(_0232_),
    .C(_0236_),
    .A(net648),
    .Y(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2651_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .C1(_0237_),
    .B1(net640),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .Y(_0238_),
    .A2(net645));
 sg13g2_a221oi_1 _2652_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0238_),
    .C1(_1723_),
    .B1(_0235_),
    .A1(_1468_),
    .Y(_0239_),
    .A2(net650));
 sg13g2_or2_1 _2653_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0240_),
    .B(net628),
    .A(net806));
 sg13g2_nand2_1 _2654_ (.Y(_0241_),
    .A(\sap_3_inst.alu.flags[0] ),
    .B(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2655_ (.Y(_0242_),
    .A(net629),
    .B(_0241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2656_ (.Y(_0243_),
    .B1(_0240_),
    .B2(_0242_),
    .A2(_1858_),
    .A1(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2657_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .C1(net643),
    .B1(net631),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .Y(_0244_),
    .A2(net650));
 sg13g2_a22oi_1 _2658_ (.Y(_0245_),
    .B1(net637),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .A2(net640),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2659_ (.Y(_0246_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .A2(net722),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2660_ (.Y(_0247_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .A2(net647),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2661_ (.B(_0245_),
    .C(_0246_),
    .A(_0244_),
    .Y(_0248_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0247_));
 sg13g2_a221oi_1 _2662_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .C1(_0248_),
    .B1(net638),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .Y(_0249_),
    .A2(net645));
 sg13g2_o21ai_1 _2663_ (.B1(_0243_),
    .VDD(VPWR),
    .Y(_0250_),
    .VSS(VGND),
    .A1(_1673_),
    .A2(_0249_));
 sg13g2_or2_1 _2664_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net17),
    .B(_0250_),
    .A(_0239_));
 sg13g2_nor4_1 _2665_ (.A(net789),
    .B(net795),
    .C(net797),
    .D(net792),
    .Y(_0251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2666_ (.A(net800),
    .B(net802),
    .C(net803),
    .D(net805),
    .Y(_0252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2667_ (.B(_0251_),
    .C(_0252_),
    .A(_1960_),
    .Y(_0253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2668_ (.A(\sap_3_inst.alu.act[1] ),
    .B(\sap_3_inst.alu.act[0] ),
    .C(\sap_3_inst.alu.act[3] ),
    .D(\sap_3_inst.alu.act[2] ),
    .Y(_0254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2669_ (.A(\sap_3_inst.alu.act[5] ),
    .B(\sap_3_inst.alu.act[4] ),
    .C(\sap_3_inst.alu.act[7] ),
    .D(\sap_3_inst.alu.act[6] ),
    .Y(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2670_ (.B(_1959_),
    .C(_0254_),
    .A(_1950_),
    .Y(_0256_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0255_));
 sg13g2_nand3_1 _2671_ (.B(_0253_),
    .C(_0256_),
    .A(_1868_),
    .Y(_0257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2672_ (.B1(_0257_),
    .VDD(VPWR),
    .Y(_0258_),
    .VSS(VGND),
    .A1(_1868_),
    .A2(net31));
 sg13g2_o21ai_1 _2673_ (.B1(_0231_),
    .VDD(VPWR),
    .Y(_0025_),
    .VSS(VGND),
    .A1(_0230_),
    .A2(_0258_));
 sg13g2_nor3_1 _2674_ (.A(net741),
    .B(net766),
    .C(_1521_),
    .Y(\sap_3_inst.clock.hlt ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2675_ (.B(_1706_),
    .C(_1752_),
    .A(_1700_),
    .Y(_0259_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1826_));
 sg13g2_o21ai_1 _2676_ (.B1(_1834_),
    .VDD(VPWR),
    .Y(_0260_),
    .VSS(VGND),
    .A1(_1731_),
    .A2(_0259_));
 sg13g2_a21oi_1 _2677_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1822_),
    .A2(_0260_),
    .Y(mem_ram_we),
    .B1(_1531_));
 sg13g2_o21ai_1 _2678_ (.B1(_1618_),
    .VDD(VPWR),
    .Y(_0261_),
    .VSS(VGND),
    .A1(net744),
    .A2(_1632_));
 sg13g2_o21ai_1 _2679_ (.B1(_1613_),
    .VDD(VPWR),
    .Y(_0262_),
    .VSS(VGND),
    .A1(net744),
    .A2(_1638_));
 sg13g2_o21ai_1 _2680_ (.B1(_1608_),
    .VDD(VPWR),
    .Y(_0263_),
    .VSS(VGND),
    .A1(net744),
    .A2(_1644_));
 sg13g2_nand3_1 _2681_ (.B(_0262_),
    .C(_0263_),
    .A(_0261_),
    .Y(_0264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2682_ (.A2(net753),
    .A1(_1582_),
    .B1(net730),
    .X(_0265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2683_ (.Y(_0266_),
    .B(_1787_),
    .A_N(_1658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2684_ (.B(_1528_),
    .C(_1585_),
    .A(net743),
    .Y(_0267_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1627_));
 sg13g2_nand2b_1 _2685_ (.Y(_0268_),
    .B(net719),
    .A_N(_1704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2686_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net749),
    .A2(_0268_),
    .Y(_0269_),
    .B1(_0266_));
 sg13g2_nand2_1 _2687_ (.Y(_0270_),
    .A(_1570_),
    .B(_1587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2688_ (.B1(_1792_),
    .VDD(VPWR),
    .Y(_0271_),
    .VSS(VGND),
    .A1(net734),
    .A2(_1617_));
 sg13g2_a221oi_1 _2689_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1638_),
    .C1(_0271_),
    .B1(_0270_),
    .A1(net750),
    .Y(_0272_),
    .A2(_1644_));
 sg13g2_nand4_1 _2690_ (.B(_0265_),
    .C(_0269_),
    .A(_1825_),
    .Y(_0273_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0272_));
 sg13g2_a21oi_1 _2691_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1630_),
    .A2(_0264_),
    .Y(_0274_),
    .B1(_0273_));
 sg13g2_a221oi_1 _2692_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1685_),
    .C1(_1787_),
    .B1(_1566_),
    .A1(net735),
    .Y(_0275_),
    .A2(_1565_));
 sg13g2_nor2b_1 _2693_ (.A(_1935_),
    .B_N(_0275_),
    .Y(_0276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2694_ (.A(net736),
    .B(_0274_),
    .C(_0276_),
    .Y(_0277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2695_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net737),
    .A2(_1559_),
    .Y(_0278_),
    .B1(_0277_));
 sg13g2_nand2_1 _2696_ (.Y(_0279_),
    .A(_1940_),
    .B(_0278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2697_ (.Y(_0280_),
    .A(_1517_),
    .B(net756),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2698_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net745),
    .A2(_1712_),
    .Y(_0281_),
    .B1(_1834_));
 sg13g2_nor2_1 _2699_ (.A(_0280_),
    .B(_0281_),
    .Y(_0282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2700_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0279_),
    .C1(_1531_),
    .B1(_0282_),
    .A1(net728),
    .Y(_0283_),
    .A2(_0280_));
 sg13g2_nor2_2 _2701_ (.A(_1764_),
    .B(_0283_),
    .Y(_0284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2702_ (.A(\sap_3_inst.controller.stage[0] ),
    .B(_0284_),
    .Y(_0001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2703_ (.A(_1536_),
    .B(_0284_),
    .Y(_0002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2704_ (.Y(_0285_),
    .A(net759),
    .B(_1507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2705_ (.A(_0284_),
    .B(_0285_),
    .Y(_0003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2706_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.controller.stage[2] ),
    .A2(_1507_),
    .Y(_0286_),
    .B1(\sap_3_inst.controller.stage[3] ));
 sg13g2_nor3_1 _2707_ (.A(_1644_),
    .B(_0284_),
    .C(_0286_),
    .Y(_0004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2708_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0238_),
    .C1(_1673_),
    .B1(_0235_),
    .A1(_1468_),
    .Y(net9),
    .A2(net650));
 sg13g2_and2_1 _2709_ (.A(net576),
    .B(_0213_),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2710_ (.A(_1673_),
    .B(_1994_),
    .Y(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2711_ (.Y(_0287_),
    .A(net576),
    .B(_1970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2712_ (.VDD(VPWR),
    .Y(net12),
    .A(_0287_),
    .VSS(VGND));
 sg13g2_and2_1 _2713_ (.A(net577),
    .B(_1919_),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2714_ (.Y(_0288_),
    .A(net576),
    .B(_1899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2715_ (.VDD(VPWR),
    .Y(net14),
    .A(_0288_),
    .VSS(VGND));
 sg13g2_and2_1 _2716_ (.A(net576),
    .B(_1876_),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2717_ (.Y(_0289_),
    .A(net577),
    .B(_1819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2718_ (.VDD(VPWR),
    .Y(net16),
    .A(_0289_),
    .VSS(VGND));
 sg13g2_o21ai_1 _2719_ (.B1(_1589_),
    .VDD(VPWR),
    .Y(_0290_),
    .VSS(VGND),
    .A1(_1697_),
    .A2(_1725_));
 sg13g2_o21ai_1 _2720_ (.B1(_1573_),
    .VDD(VPWR),
    .Y(_0291_),
    .VSS(VGND),
    .A1(_1609_),
    .A2(_1648_));
 sg13g2_nor3_1 _2721_ (.A(_1661_),
    .B(_1662_),
    .C(_1696_),
    .Y(_0292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2722_ (.A(net752),
    .B(net750),
    .C(_1634_),
    .Y(_0293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2723_ (.A(net744),
    .B(_1683_),
    .C(_0293_),
    .X(_0294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2724_ (.Y(_0295_),
    .B1(_0294_),
    .B2(_1601_),
    .A2(_0291_),
    .A1(_0290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2725_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0292_),
    .A2(_0295_),
    .Y(_0296_),
    .B1(_1556_));
 sg13g2_o21ai_1 _2726_ (.B1(_1539_),
    .VDD(VPWR),
    .Y(_0297_),
    .VSS(VGND),
    .A1(_1544_),
    .A2(_0296_));
 sg13g2_nand2_1 _2727_ (.Y(_0298_),
    .A(net757),
    .B(_0297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2728_ (.Y(_0299_),
    .B1(_1538_),
    .B2(_0298_),
    .A2(_1505_),
    .A1(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2729_ (.VDD(VPWR),
    .Y(mem_mar_we),
    .A(_0299_),
    .VSS(VGND));
 sg13g2_nor2_2 _2730_ (.A(\u_ser.state[1] ),
    .B(\u_ser.state[0] ),
    .Y(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2731_ (.A0(net69),
    .A1(\sap_3_inst.out[0] ),
    .S(net813),
    .X(_0017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2732_ (.A0(net59),
    .A1(\sap_3_inst.out[1] ),
    .S(net813),
    .X(_0018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2733_ (.A0(net64),
    .A1(\sap_3_inst.out[2] ),
    .S(net813),
    .X(_0019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2734_ (.A0(net58),
    .A1(\sap_3_inst.out[3] ),
    .S(net813),
    .X(_0020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2735_ (.A0(net67),
    .A1(\sap_3_inst.out[4] ),
    .S(net813),
    .X(_0021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2736_ (.A0(net66),
    .A1(\sap_3_inst.out[5] ),
    .S(net813),
    .X(_0022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2737_ (.A0(net65),
    .A1(\sap_3_inst.out[6] ),
    .S(_0185_),
    .X(_0023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2738_ (.A0(net68),
    .A1(\sap_3_inst.out[7] ),
    .S(_0185_),
    .X(_0024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2739_ (.B(net729),
    .C(_1715_),
    .A(_1516_),
    .Y(_0300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2740_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1549_),
    .A2(_1717_),
    .Y(_0301_),
    .B1(_1551_));
 sg13g2_o21ai_1 _2741_ (.B1(net748),
    .VDD(VPWR),
    .Y(_0302_),
    .VSS(VGND),
    .A1(net763),
    .A2(_1570_));
 sg13g2_and2_1 _2742_ (.A(_1551_),
    .B(_1742_),
    .X(_0303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2743_ (.B(net728),
    .C(_1715_),
    .A(_1616_),
    .Y(_0304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2744_ (.B(_1848_),
    .C(_0303_),
    .A(_1843_),
    .Y(_0305_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0304_));
 sg13g2_a21oi_1 _2745_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1685_),
    .A2(_0302_),
    .Y(_0306_),
    .B1(_0305_));
 sg13g2_o21ai_1 _2746_ (.B1(_1713_),
    .VDD(VPWR),
    .Y(_0307_),
    .VSS(VGND),
    .A1(_0301_),
    .A2(_0306_));
 sg13g2_nor3_1 _2747_ (.A(net741),
    .B(_1515_),
    .C(_1716_),
    .Y(_0308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2748_ (.A(_1713_),
    .B(_1856_),
    .C(_0308_),
    .Y(_0309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2749_ (.Y(_0310_),
    .A(_1517_),
    .B(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2750_ (.B1(_0300_),
    .VDD(VPWR),
    .Y(_0311_),
    .VSS(VGND),
    .A1(_0309_),
    .A2(_0310_));
 sg13g2_a21oi_1 _2751_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net736),
    .A2(_1824_),
    .Y(_0312_),
    .B1(net724));
 sg13g2_o21ai_1 _2752_ (.B1(_0312_),
    .VDD(VPWR),
    .Y(_0313_),
    .VSS(VGND),
    .A1(net736),
    .A2(_1827_));
 sg13g2_o21ai_1 _2753_ (.B1(_0313_),
    .VDD(VPWR),
    .Y(_0314_),
    .VSS(VGND),
    .A1(_1543_),
    .A2(net732));
 sg13g2_nand2b_1 _2754_ (.Y(_0315_),
    .B(_1945_),
    .A_N(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2755_ (.A(_1951_),
    .B(_1958_),
    .Y(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2756_ (.A(_1947_),
    .B(_1949_),
    .X(_0317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2757_ (.A(_1955_),
    .B(_1957_),
    .Y(_0318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2758_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0319_),
    .B(_1957_),
    .A(_1955_));
 sg13g2_a21oi_1 _2759_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0317_),
    .A2(_0319_),
    .Y(_0320_),
    .B1(_0316_));
 sg13g2_o21ai_1 _2760_ (.B1(_0320_),
    .VDD(VPWR),
    .Y(_0321_),
    .VSS(VGND),
    .A1(net626),
    .A2(_0315_));
 sg13g2_nand2_1 _2761_ (.Y(_0322_),
    .A(net806),
    .B(\sap_3_inst.alu.tmp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2762_ (.B(\sap_3_inst.alu.tmp[0] ),
    .A(net806),
    .X(_0323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2763_ (.Y(_0324_),
    .A(_0317_),
    .B(_0318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2764_ (.A(net714),
    .B_N(_0324_),
    .Y(_0325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2765_ (.A(_1950_),
    .B(_1958_),
    .Y(_0326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2766_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0327_),
    .B(_1958_),
    .A(_1950_));
 sg13g2_or2_1 _2767_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0328_),
    .B(_0319_),
    .A(_0201_));
 sg13g2_inv_2 _2768_ (.Y(_0329_),
    .A(_0328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2769_ (.Y(_0330_),
    .A(_0327_),
    .B(_0328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2770_ (.Y(_0331_),
    .A(_1955_),
    .B(_1957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2771_ (.A(_0201_),
    .B(_0331_),
    .Y(_0332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2772_ (.A(_0200_),
    .B(_0330_),
    .C(net625),
    .Y(_0333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2773_ (.A(_0325_),
    .B(_0333_),
    .X(_0334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2774_ (.A(_1951_),
    .B(_0319_),
    .Y(_0335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2775_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0336_),
    .B(_0319_),
    .A(_1951_));
 sg13g2_or3_1 _2776_ (.A(net625),
    .B(net574),
    .C(_0335_),
    .X(_0337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2777_ (.A(_1956_),
    .B(_0199_),
    .Y(_0338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2778_ (.B(_1957_),
    .C(net683),
    .A(net762),
    .Y(_0339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2779_ (.A(_1955_),
    .B(_0199_),
    .Y(_0340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2780_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net803),
    .A2(net682),
    .Y(_0341_),
    .B1(net708));
 sg13g2_nor2_2 _2781_ (.A(_1951_),
    .B(_0331_),
    .Y(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2782_ (.B1(_0342_),
    .VDD(VPWR),
    .Y(_0343_),
    .VSS(VGND),
    .A1(net806),
    .A2(\sap_3_inst.alu.tmp[0] ));
 sg13g2_nor3_2 _2783_ (.A(net775),
    .B(_1951_),
    .C(_1956_),
    .Y(_0344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2784_ (.Y(_0345_),
    .B(_0344_),
    .A_N(_0322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2785_ (.A(_0339_),
    .B(_0341_),
    .C(_0343_),
    .D(_0345_),
    .X(_0346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2786_ (.Y(_0347_),
    .A(net762),
    .B(_0323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2787_ (.Y(_0348_),
    .B(net762),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0323_));
 sg13g2_xor2_1 _2788_ (.B(_0323_),
    .A(net762),
    .X(_0349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2789_ (.B1(_0346_),
    .VDD(VPWR),
    .Y(_0350_),
    .VSS(VGND),
    .A1(net805),
    .A2(_0325_));
 sg13g2_a221oi_1 _2790_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0330_),
    .C1(_0350_),
    .B1(_0349_),
    .A1(_0323_),
    .Y(_0351_),
    .A2(_0337_));
 sg13g2_nand2b_1 _2791_ (.Y(_0352_),
    .B(net708),
    .A_N(\sap_3_inst.alu.act[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2792_ (.A(net626),
    .B(_0351_),
    .Y(_0353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2793_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0353_),
    .C1(net580),
    .B1(_0352_),
    .A1(net31),
    .Y(_0354_),
    .A2(net626));
 sg13g2_a21oi_1 _2794_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1459_),
    .A2(net580),
    .Y(_0033_),
    .B1(_0354_));
 sg13g2_nand2_1 _2795_ (.Y(_0355_),
    .A(net803),
    .B(\sap_3_inst.alu.tmp[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2796_ (.B(\sap_3_inst.alu.tmp[1] ),
    .A(net804),
    .X(_0356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2797_ (.Y(_0357_),
    .A(net804),
    .B(\sap_3_inst.alu.tmp[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2798_ (.Y(_0358_),
    .B(\sap_3_inst.alu.tmp[0] ),
    .A_N(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2799_ (.Y(_0359_),
    .A(_0356_),
    .B(_0358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2800_ (.A(_0348_),
    .B(_0359_),
    .Y(_0360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2801_ (.Y(_0361_),
    .A(_0348_),
    .B(_0359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2802_ (.A(net775),
    .B(_1951_),
    .C(_1956_),
    .D(_0355_),
    .Y(_0362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2803_ (.A(_1458_),
    .B(_1550_),
    .C(_1796_),
    .Y(_0363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2804_ (.B1(_1458_),
    .VDD(VPWR),
    .Y(_0364_),
    .VSS(VGND),
    .A1(_1550_),
    .A2(_1796_));
 sg13g2_nor2b_1 _2805_ (.A(_0363_),
    .B_N(_0364_),
    .Y(_0365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2806_ (.B1(net714),
    .VDD(VPWR),
    .Y(_0366_),
    .VSS(VGND),
    .A1(net805),
    .A2(_0365_));
 sg13g2_a21oi_1 _2807_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net805),
    .A2(_0365_),
    .Y(_0367_),
    .B1(_0366_));
 sg13g2_a221oi_1 _2808_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net801),
    .C1(_0367_),
    .B1(net682),
    .A1(net806),
    .Y(_0368_),
    .A2(net683));
 sg13g2_o21ai_1 _2809_ (.B1(_0342_),
    .VDD(VPWR),
    .Y(_0369_),
    .VSS(VGND),
    .A1(net803),
    .A2(\sap_3_inst.alu.tmp[1] ));
 sg13g2_nand3_1 _2810_ (.B(_0323_),
    .C(_0356_),
    .A(net762),
    .Y(_0370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2811_ (.Y(_0371_),
    .A(_0322_),
    .B(_0357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2812_ (.Y(_0372_),
    .A(_0347_),
    .B(_0371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2813_ (.B(_0370_),
    .C(_0372_),
    .A(_0329_),
    .Y(_0373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2814_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net625),
    .C1(_0362_),
    .B1(_0359_),
    .A1(_0335_),
    .Y(_0374_),
    .A2(_0356_));
 sg13g2_o21ai_1 _2815_ (.B1(_0369_),
    .VDD(VPWR),
    .Y(_0375_),
    .VSS(VGND),
    .A1(net804),
    .A2(_0324_));
 sg13g2_a21oi_1 _2816_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0326_),
    .A2(_0361_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_nand4_1 _2817_ (.B(_0373_),
    .C(_0374_),
    .A(_0368_),
    .Y(_0377_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0376_));
 sg13g2_a21oi_1 _2818_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net574),
    .A2(_0371_),
    .Y(_0378_),
    .B1(net708));
 sg13g2_o21ai_1 _2819_ (.B1(_0378_),
    .VDD(VPWR),
    .Y(_0379_),
    .VSS(VGND),
    .A1(net574),
    .A2(_0377_));
 sg13g2_a21oi_1 _2820_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu.act[1] ),
    .A2(net708),
    .Y(_0380_),
    .B1(net626));
 sg13g2_a221oi_1 _2821_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0380_),
    .C1(net580),
    .B1(_0379_),
    .A1(_0227_),
    .Y(_0381_),
    .A2(net626));
 sg13g2_a21o_1 _2822_ (.A2(net580),
    .A1(net803),
    .B1(_0381_),
    .X(_0034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2823_ (.A(net802),
    .B(\sap_3_inst.alu.tmp[2] ),
    .X(_0382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2824_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0383_),
    .B(\sap_3_inst.alu.tmp[2] ),
    .A(net802));
 sg13g2_nor2b_2 _2825_ (.A(_0382_),
    .B_N(_0383_),
    .Y(_0384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2826_ (.A(\sap_3_inst.alu.tmp[1] ),
    .B_N(net804),
    .Y(_0385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2827_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0357_),
    .A2(_0358_),
    .Y(_0386_),
    .B1(_0385_));
 sg13g2_nor2_1 _2828_ (.A(_0384_),
    .B(_0386_),
    .Y(_0387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2829_ (.B(_0386_),
    .A(_0384_),
    .X(_0388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2830_ (.Y(_0389_),
    .B(_0360_),
    .A_N(_0388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2831_ (.B(_0388_),
    .A(_0360_),
    .X(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2832_ (.Y(_0391_),
    .A(net625),
    .B(_0388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2833_ (.Y(_0392_),
    .A(_0344_),
    .B(_0382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2834_ (.Y(_0393_),
    .A(net801),
    .B(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2835_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net805),
    .A2(_0364_),
    .Y(_0394_),
    .B1(_0363_));
 sg13g2_nor2_1 _2836_ (.A(_0393_),
    .B(_0394_),
    .Y(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2837_ (.Y(_0396_),
    .B(net714),
    .A_N(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2838_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0393_),
    .A2(_0394_),
    .Y(_0397_),
    .B1(_0396_));
 sg13g2_o21ai_1 _2839_ (.B1(_0355_),
    .VDD(VPWR),
    .Y(_0398_),
    .VSS(VGND),
    .A1(_0322_),
    .A2(_0357_));
 sg13g2_xor2_1 _2840_ (.B(_0398_),
    .A(_0384_),
    .X(_0399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2841_ (.A(_0370_),
    .B_N(_0399_),
    .Y(_0400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2842_ (.Y(_0401_),
    .A(_0370_),
    .B(_0399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2843_ (.B1(_0391_),
    .VDD(VPWR),
    .Y(_0402_),
    .VSS(VGND),
    .A1(net802),
    .A2(_0324_));
 sg13g2_a22oi_1 _2844_ (.Y(_0403_),
    .B1(_0390_),
    .B2(_0326_),
    .A2(_0384_),
    .A1(_0335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2845_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net800),
    .C1(_0397_),
    .B1(net682),
    .A1(net804),
    .Y(_0404_),
    .A2(net683));
 sg13g2_a22oi_1 _2846_ (.Y(_0405_),
    .B1(_0401_),
    .B2(_0329_),
    .A2(_0383_),
    .A1(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2847_ (.B(_0403_),
    .C(_0404_),
    .A(_0392_),
    .Y(_0406_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0405_));
 sg13g2_nor3_1 _2848_ (.A(net574),
    .B(_0402_),
    .C(_0406_),
    .Y(_0407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2849_ (.A(_0399_),
    .B_N(net574),
    .Y(_0408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2850_ (.A(net708),
    .B(_0407_),
    .C(_0408_),
    .X(_0409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2851_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu.act[2] ),
    .A2(net708),
    .Y(_0410_),
    .B1(net626));
 sg13g2_a221oi_1 _2852_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0410_),
    .C1(net580),
    .B1(_0409_),
    .A1(_2008_),
    .Y(_0411_),
    .A2(net626));
 sg13g2_a21o_1 _2853_ (.A2(net580),
    .A1(net801),
    .B1(_0411_),
    .X(_0035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2854_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net801),
    .A2(net721),
    .Y(_0412_),
    .B1(_0395_));
 sg13g2_nand2_1 _2855_ (.Y(_0413_),
    .A(net798),
    .B(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2856_ (.A(net798),
    .B(net720),
    .Y(_0414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2857_ (.Y(_0415_),
    .A(net798),
    .B(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2858_ (.B1(net714),
    .VDD(VPWR),
    .Y(_0416_),
    .VSS(VGND),
    .A1(_0412_),
    .A2(_0415_));
 sg13g2_a21oi_1 _2859_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0412_),
    .A2(_0415_),
    .Y(_0417_),
    .B1(_0416_));
 sg13g2_nand2_1 _2860_ (.Y(_0418_),
    .A(net798),
    .B(\sap_3_inst.alu.tmp[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2861_ (.B(\sap_3_inst.alu.tmp[3] ),
    .C(_0344_),
    .A(net798),
    .Y(_0419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2862_ (.B1(_0419_),
    .VDD(VPWR),
    .Y(_0420_),
    .VSS(VGND),
    .A1(net799),
    .A2(_0324_));
 sg13g2_nor2_1 _2863_ (.A(net798),
    .B(\sap_3_inst.alu.tmp[3] ),
    .Y(_0421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2864_ (.B(\sap_3_inst.alu.tmp[3] ),
    .A(net799),
    .X(_0422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2865_ (.Y(_0423_),
    .A(net799),
    .B(\sap_3_inst.alu.tmp[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2866_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0384_),
    .A2(_0398_),
    .Y(_0424_),
    .B1(_0382_));
 sg13g2_xnor2_1 _2867_ (.Y(_0425_),
    .A(_0423_),
    .B(_0424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2868_ (.VDD(VPWR),
    .Y(_0426_),
    .A(_0425_),
    .VSS(VGND));
 sg13g2_nand2_2 _2869_ (.Y(_0427_),
    .A(_0400_),
    .B(_0426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2870_ (.Y(_0428_),
    .A(_0400_),
    .B(_0425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2871_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0329_),
    .C1(_0420_),
    .B1(_0428_),
    .A1(_0335_),
    .Y(_0429_),
    .A2(_0422_));
 sg13g2_nor3_1 _2872_ (.A(_1951_),
    .B(_0331_),
    .C(_0421_),
    .Y(_0430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2873_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net796),
    .C1(_0430_),
    .B1(net682),
    .A1(net801),
    .Y(_0431_),
    .A2(net683));
 sg13g2_a21oi_1 _2874_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_1471_),
    .Y(_0432_),
    .B1(_0387_));
 sg13g2_nor2_1 _2875_ (.A(_0422_),
    .B(_0432_),
    .Y(_0433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2876_ (.Y(_0434_),
    .A(_0423_),
    .B(_0432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2877_ (.A(_0348_),
    .B(_0359_),
    .C(_0384_),
    .Y(_0435_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0422_));
 sg13g2_a21o_1 _2878_ (.A2(_0434_),
    .A1(_0389_),
    .B1(_0435_),
    .X(_0436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2879_ (.Y(_0437_),
    .B1(_0436_),
    .B2(_0326_),
    .A2(_0434_),
    .A1(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2880_ (.B(_0431_),
    .C(_0437_),
    .A(_0429_),
    .Y(_0438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2881_ (.A(net574),
    .B(_0417_),
    .C(_0438_),
    .Y(_0439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2882_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net574),
    .A2(_0425_),
    .Y(_0440_),
    .B1(net707));
 sg13g2_nand2b_1 _2883_ (.Y(_0441_),
    .B(_0440_),
    .A_N(_0439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2884_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu.act[3] ),
    .A2(net708),
    .Y(_0442_),
    .B1(net626));
 sg13g2_a221oi_1 _2885_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0442_),
    .C1(net580),
    .B1(_0441_),
    .A1(net572),
    .Y(_0443_),
    .A2(net627));
 sg13g2_a21o_1 _2886_ (.A2(net580),
    .A1(net799),
    .B1(_0443_),
    .X(_0036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2887_ (.A(net32),
    .B_N(net627),
    .Y(_0444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2888_ (.Y(_0445_),
    .A(net796),
    .B(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2889_ (.VDD(VPWR),
    .Y(_0446_),
    .A(_0445_),
    .VSS(VGND));
 sg13g2_a21oi_1 _2890_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0412_),
    .A2(_0413_),
    .Y(_0447_),
    .B1(_0414_));
 sg13g2_and2_1 _2891_ (.A(_0446_),
    .B(_0447_),
    .X(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2892_ (.B1(net714),
    .VDD(VPWR),
    .Y(_0449_),
    .VSS(VGND),
    .A1(_0446_),
    .A2(_0447_));
 sg13g2_nor2_1 _2893_ (.A(_1460_),
    .B(_1473_),
    .Y(_0450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2894_ (.Y(_0451_),
    .A(net797),
    .B(\sap_3_inst.alu.tmp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2895_ (.VDD(VPWR),
    .Y(_0452_),
    .A(_0451_),
    .VSS(VGND));
 sg13g2_nand2_1 _2896_ (.Y(_0453_),
    .A(_0344_),
    .B(_0450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2897_ (.B1(_0453_),
    .VDD(VPWR),
    .Y(_0454_),
    .VSS(VGND),
    .A1(_0336_),
    .A2(_0451_));
 sg13g2_o21ai_1 _2898_ (.B1(_0342_),
    .VDD(VPWR),
    .Y(_0455_),
    .VSS(VGND),
    .A1(net796),
    .A2(\sap_3_inst.alu.tmp[4] ));
 sg13g2_o21ai_1 _2899_ (.B1(_0455_),
    .VDD(VPWR),
    .Y(_0456_),
    .VSS(VGND),
    .A1(net796),
    .A2(_0324_));
 sg13g2_a21oi_1 _2900_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0418_),
    .A2(_0424_),
    .Y(_0457_),
    .B1(_0421_));
 sg13g2_xnor2_1 _2901_ (.Y(_0458_),
    .A(_0452_),
    .B(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2902_ (.A(_0427_),
    .B(_0458_),
    .Y(_0459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2903_ (.Y(_0460_),
    .A(_0427_),
    .B(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2904_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net798),
    .A2(_1472_),
    .Y(_0461_),
    .B1(_0433_));
 sg13g2_nor2_1 _2905_ (.A(_0452_),
    .B(_0461_),
    .Y(_0462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2906_ (.Y(_0463_),
    .A(_0451_),
    .B(_0461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2907_ (.Y(_0464_),
    .A(_0435_),
    .B(_0451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2908_ (.B(_0463_),
    .A(_0435_),
    .X(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2909_ (.Y(_0466_),
    .A(net625),
    .B(_0463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2910_ (.Y(_0467_),
    .B1(net682),
    .B2(net793),
    .A2(net683),
    .A1(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2911_ (.Y(_0468_),
    .A(_0466_),
    .B(_0467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2912_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0326_),
    .A2(_0465_),
    .Y(_0469_),
    .B1(_0468_));
 sg13g2_o21ai_1 _2913_ (.B1(_0469_),
    .VDD(VPWR),
    .Y(_0470_),
    .VSS(VGND),
    .A1(_0328_),
    .A2(_0460_));
 sg13g2_nor4_1 _2914_ (.A(net574),
    .B(_0454_),
    .C(_0456_),
    .D(_0470_),
    .Y(_0471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2915_ (.B1(_0471_),
    .VDD(VPWR),
    .Y(_0472_),
    .VSS(VGND),
    .A1(_0448_),
    .A2(_0449_));
 sg13g2_a21oi_1 _2916_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net575),
    .A2(_0458_),
    .Y(_0473_),
    .B1(net707));
 sg13g2_a221oi_1 _2917_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0473_),
    .C1(net627),
    .B1(_0472_),
    .A1(\sap_3_inst.alu.act[4] ),
    .Y(_0474_),
    .A2(net707));
 sg13g2_nor3_1 _2918_ (.A(net581),
    .B(_0444_),
    .C(_0474_),
    .Y(_0475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2919_ (.A2(net581),
    .A1(net797),
    .B1(_0475_),
    .X(_0037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2920_ (.A(net573),
    .B_N(net627),
    .Y(_0476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2921_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net796),
    .A2(net720),
    .Y(_0477_),
    .B1(_0448_));
 sg13g2_nand2_1 _2922_ (.Y(_0478_),
    .A(net793),
    .B(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2923_ (.Y(_0479_),
    .A(net793),
    .B(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2924_ (.B1(net714),
    .VDD(VPWR),
    .Y(_0480_),
    .VSS(VGND),
    .A1(_0477_),
    .A2(_0479_));
 sg13g2_a21oi_1 _2925_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0477_),
    .A2(_0479_),
    .Y(_0481_),
    .B1(_0480_));
 sg13g2_nand2_1 _2926_ (.Y(_0482_),
    .A(net793),
    .B(\sap_3_inst.alu.tmp[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2927_ (.A(net794),
    .B(\sap_3_inst.alu.tmp[5] ),
    .Y(_0483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2928_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0484_),
    .B(\sap_3_inst.alu.tmp[5] ),
    .A(net794));
 sg13g2_and2_1 _2929_ (.A(_0482_),
    .B(_0484_),
    .X(_0485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2930_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0452_),
    .A2(_0457_),
    .Y(_0486_),
    .B1(_0450_));
 sg13g2_xnor2_1 _2931_ (.Y(_0487_),
    .A(_0485_),
    .B(_0486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2932_ (.VDD(VPWR),
    .Y(_0488_),
    .A(_0487_),
    .VSS(VGND));
 sg13g2_nand2_1 _2933_ (.Y(_0489_),
    .A(_0459_),
    .B(_0487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2934_ (.Y(_0490_),
    .A(_0459_),
    .B(_0487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2935_ (.B(\sap_3_inst.alu.tmp[5] ),
    .C(_0344_),
    .A(net794),
    .Y(_0491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2936_ (.Y(_0492_),
    .B1(_0485_),
    .B2(_0335_),
    .A2(_0484_),
    .A1(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2937_ (.A(net793),
    .B(_0324_),
    .Y(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2938_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net790),
    .C1(_0493_),
    .B1(net682),
    .A1(net796),
    .Y(_0494_),
    .A2(net683));
 sg13g2_a21oi_1 _2939_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net796),
    .A2(_1473_),
    .Y(_0495_),
    .B1(_0462_));
 sg13g2_xor2_1 _2940_ (.B(_0495_),
    .A(_0485_),
    .X(_0496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2941_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0497_),
    .B(_0485_),
    .A(_0464_));
 sg13g2_or2_1 _2942_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0498_),
    .B(_0497_),
    .A(_0327_));
 sg13g2_nand4_1 _2943_ (.B(_0492_),
    .C(_0494_),
    .A(_0491_),
    .Y(_0499_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0498_));
 sg13g2_and2_1 _2944_ (.A(_0326_),
    .B(_0464_),
    .X(_0500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2945_ (.B1(_0496_),
    .VDD(VPWR),
    .Y(_0501_),
    .VSS(VGND),
    .A1(net625),
    .A2(_0500_));
 sg13g2_o21ai_1 _2946_ (.B1(_0501_),
    .VDD(VPWR),
    .Y(_0502_),
    .VSS(VGND),
    .A1(_0328_),
    .A2(_0490_));
 sg13g2_or4_1 _2947_ (.A(net575),
    .B(_0481_),
    .C(_0499_),
    .D(_0502_),
    .X(_0503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2948_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net575),
    .A2(_0488_),
    .Y(_0504_),
    .B1(net707));
 sg13g2_a221oi_1 _2949_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0504_),
    .C1(net627),
    .B1(_0503_),
    .A1(\sap_3_inst.alu.act[5] ),
    .Y(_0505_),
    .A2(net707));
 sg13g2_nor3_1 _2950_ (.A(net581),
    .B(_0476_),
    .C(_0505_),
    .Y(_0506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2951_ (.A2(net581),
    .A1(net794),
    .B1(_0506_),
    .X(_0038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2952_ (.A(net33),
    .B_N(_0311_),
    .Y(_0507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2953_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0508_),
    .B(\sap_3_inst.alu.tmp[6] ),
    .A(net791));
 sg13g2_and2_1 _2954_ (.A(net791),
    .B(\sap_3_inst.alu.tmp[6] ),
    .X(_0509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2955_ (.B(\sap_3_inst.alu.tmp[6] ),
    .A(net790),
    .X(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2956_ (.Y(_0511_),
    .A(net791),
    .B(\sap_3_inst.alu.tmp[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2957_ (.A(net794),
    .B_N(\sap_3_inst.alu.tmp[5] ),
    .Y(_0512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2958_ (.Y(_0513_),
    .B(net794),
    .A_N(\sap_3_inst.alu.tmp[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2959_ (.B1(_0513_),
    .VDD(VPWR),
    .Y(_0514_),
    .VSS(VGND),
    .A1(_0495_),
    .A2(_0512_));
 sg13g2_xnor2_1 _2960_ (.Y(_0515_),
    .A(_0510_),
    .B(_0514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2961_ (.A(_0497_),
    .B(_0515_),
    .Y(_0516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2962_ (.A(net790),
    .B(_0324_),
    .Y(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2963_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net794),
    .A2(net683),
    .Y(_0518_),
    .B1(_0517_));
 sg13g2_a22oi_1 _2964_ (.Y(_0519_),
    .B1(_0342_),
    .B2(_0508_),
    .A2(_0340_),
    .A1(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2965_ (.Y(_0520_),
    .B1(_0510_),
    .B2(_0335_),
    .A2(_0509_),
    .A1(_0344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2966_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0326_),
    .A2(_0497_),
    .Y(_0521_),
    .B1(_0332_));
 sg13g2_nand2b_1 _2967_ (.Y(_0522_),
    .B(_0515_),
    .A_N(_0521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2968_ (.A(_0518_),
    .B(_0519_),
    .C(_0520_),
    .D(_0522_),
    .X(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2969_ (.B1(_0482_),
    .VDD(VPWR),
    .Y(_0524_),
    .VSS(VGND),
    .A1(_0483_),
    .A2(_0486_));
 sg13g2_xnor2_1 _2970_ (.Y(_0525_),
    .A(_0510_),
    .B(_0524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2971_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0526_),
    .B(_0525_),
    .A(_0489_));
 sg13g2_a21oi_1 _2972_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0489_),
    .A2(_0525_),
    .Y(_0527_),
    .B1(_0328_));
 sg13g2_a221oi_1 _2973_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0527_),
    .C1(net575),
    .B1(_0526_),
    .A1(_0326_),
    .Y(_0528_),
    .A2(_0516_));
 sg13g2_nand2_1 _2974_ (.Y(_0529_),
    .A(net790),
    .B(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2975_ (.Y(_0530_),
    .A(net790),
    .B(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2976_ (.Y(_0531_),
    .A(_0477_),
    .B(_0478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2977_ (.B1(_0531_),
    .VDD(VPWR),
    .Y(_0532_),
    .VSS(VGND),
    .A1(net793),
    .A2(net721));
 sg13g2_nand2_1 _2978_ (.Y(_0533_),
    .A(_0530_),
    .B(_0532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2979_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0534_),
    .B(_0532_),
    .A(_0530_));
 sg13g2_nand3_1 _2980_ (.B(_0533_),
    .C(_0534_),
    .A(_1944_),
    .Y(_0535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2981_ (.B(_0528_),
    .C(_0535_),
    .A(_0523_),
    .Y(_0536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2982_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net575),
    .A2(_0525_),
    .Y(_0537_),
    .B1(net707));
 sg13g2_a221oi_1 _2983_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0537_),
    .C1(net627),
    .B1(_0536_),
    .A1(\sap_3_inst.alu.act[6] ),
    .Y(_0538_),
    .A2(net707));
 sg13g2_nor3_1 _2984_ (.A(net581),
    .B(_0507_),
    .C(_0538_),
    .Y(_0539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2985_ (.A2(net581),
    .A1(net791),
    .B1(_0539_),
    .X(_0039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2986_ (.Y(_0540_),
    .A(net788),
    .B(net581),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2987_ (.Y(_0541_),
    .B(_0311_),
    .A_N(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2988_ (.Y(_0542_),
    .A(_0529_),
    .B(_0534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2989_ (.Y(_0543_),
    .A(net788),
    .B(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2990_ (.Y(_0544_),
    .A(_0542_),
    .B(_0543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2991_ (.A(net787),
    .B(\sap_3_inst.alu.tmp[7] ),
    .Y(_0545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2992_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0546_),
    .B(\sap_3_inst.alu.tmp[7] ),
    .A(net787));
 sg13g2_and2_1 _2993_ (.A(net787),
    .B(\sap_3_inst.alu.tmp[7] ),
    .X(_0547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2994_ (.Y(_0548_),
    .A(net787),
    .B(\sap_3_inst.alu.tmp[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2995_ (.Y(_0549_),
    .A(_0546_),
    .B(_0548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2996_ (.A(\sap_3_inst.alu.tmp[6] ),
    .B_N(net791),
    .Y(_0550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2997_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0511_),
    .A2(_0514_),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_xnor2_1 _2998_ (.Y(_0552_),
    .A(_0549_),
    .B(_0551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2999_ (.Y(_0553_),
    .A(_0516_),
    .B(_0552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3000_ (.A(_0332_),
    .B(_0552_),
    .X(_0554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3001_ (.X(_0555_),
    .A(\sap_3_inst.alu.flags[1] ),
    .B(_1957_),
    .C(net682),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3002_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net790),
    .A2(_0338_),
    .Y(_0556_),
    .B1(_0555_));
 sg13g2_a22oi_1 _3003_ (.Y(_0557_),
    .B1(_0547_),
    .B2(_0344_),
    .A2(_0546_),
    .A1(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3004_ (.B1(_0557_),
    .VDD(VPWR),
    .Y(_0558_),
    .VSS(VGND),
    .A1(net787),
    .A2(_0324_));
 sg13g2_o21ai_1 _3005_ (.B1(_0556_),
    .VDD(VPWR),
    .Y(_0559_),
    .VSS(VGND),
    .A1(_0336_),
    .A2(_0549_));
 sg13g2_nor4_1 _3006_ (.A(net575),
    .B(_0554_),
    .C(_0558_),
    .D(_0559_),
    .Y(_0560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3007_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0510_),
    .A2(_0524_),
    .Y(_0561_),
    .B1(_0509_));
 sg13g2_xnor2_1 _3008_ (.Y(_0562_),
    .A(_0549_),
    .B(_0561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3009_ (.B(_0562_),
    .A(_0526_),
    .X(_0563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3010_ (.B1(_0560_),
    .VDD(VPWR),
    .Y(_0564_),
    .VSS(VGND),
    .A1(_0327_),
    .A2(_0553_));
 sg13g2_a221oi_1 _3011_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0329_),
    .C1(_0564_),
    .B1(_0563_),
    .A1(_1944_),
    .Y(_0565_),
    .A2(_0544_));
 sg13g2_a21o_1 _3012_ (.A2(_0562_),
    .A1(net575),
    .B1(net707),
    .X(_0566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3013_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu.act[7] ),
    .A2(_0314_),
    .Y(_0567_),
    .B1(net627));
 sg13g2_o21ai_1 _3014_ (.B1(_0567_),
    .VDD(VPWR),
    .Y(_0568_),
    .VSS(VGND),
    .A1(_0565_),
    .A2(_0566_));
 sg13g2_nand2_1 _3015_ (.Y(_0569_),
    .A(_0541_),
    .B(_0568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3016_ (.B1(_0540_),
    .VDD(VPWR),
    .Y(_0040_),
    .VSS(VGND),
    .A1(net581),
    .A2(_0569_));
 sg13g2_nand2_1 _3017_ (.Y(_0570_),
    .A(\sap_3_inst.out[0] ),
    .B(net717),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3018_ (.B1(_0570_),
    .VDD(VPWR),
    .Y(_0041_),
    .VSS(VGND),
    .A1(_1459_),
    .A2(net717));
 sg13g2_nand2_1 _3019_ (.Y(_0571_),
    .A(\sap_3_inst.out[1] ),
    .B(net717),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3020_ (.B1(_0571_),
    .VDD(VPWR),
    .Y(_0042_),
    .VSS(VGND),
    .A1(_1458_),
    .A2(net717));
 sg13g2_mux2_1 _3021_ (.A0(net801),
    .A1(\sap_3_inst.out[2] ),
    .S(net717),
    .X(_0043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3022_ (.Y(_0572_),
    .A(\sap_3_inst.out[3] ),
    .B(net717),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3023_ (.B1(_0572_),
    .VDD(VPWR),
    .Y(_0044_),
    .VSS(VGND),
    .A1(_1445_),
    .A2(net717));
 sg13g2_nand2_1 _3024_ (.Y(_0573_),
    .A(\sap_3_inst.out[4] ),
    .B(net717),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3025_ (.B1(_0573_),
    .VDD(VPWR),
    .Y(_0045_),
    .VSS(VGND),
    .A1(_1460_),
    .A2(net718));
 sg13g2_mux2_1 _3026_ (.A0(net793),
    .A1(\sap_3_inst.out[5] ),
    .S(net718),
    .X(_0046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3027_ (.A0(net790),
    .A1(\sap_3_inst.out[6] ),
    .S(net718),
    .X(_0047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3028_ (.A0(net788),
    .A1(\sap_3_inst.out[7] ),
    .S(net718),
    .X(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3029_ (.Y(_0574_),
    .A(_0202_),
    .B(_0333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3030_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0548_),
    .A2(_0561_),
    .Y(_0575_),
    .B1(_0545_));
 sg13g2_nor4_1 _3031_ (.A(_0427_),
    .B(_0451_),
    .C(_0511_),
    .D(_0549_),
    .Y(_0576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3032_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0485_),
    .A2(_0576_),
    .Y(_0577_),
    .B1(_0575_));
 sg13g2_a21oi_1 _3033_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0328_),
    .A2(_0574_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_nor4_1 _3034_ (.A(_0327_),
    .B(_0497_),
    .C(_0515_),
    .D(_0552_),
    .Y(_0579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3035_ (.A(net787),
    .B_N(\sap_3_inst.alu.tmp[7] ),
    .Y(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3036_ (.Y(_0581_),
    .B(net787),
    .A_N(\sap_3_inst.alu.tmp[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3037_ (.B1(_0581_),
    .VDD(VPWR),
    .Y(_0582_),
    .VSS(VGND),
    .A1(_0551_),
    .A2(_0580_));
 sg13g2_nor2_1 _3038_ (.A(_0326_),
    .B(net625),
    .Y(_0583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3039_ (.Y(_0584_),
    .A(net775),
    .B(_0317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3040_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu.flags[1] ),
    .A2(_1956_),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_a221oi_1 _3041_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net805),
    .C1(_0585_),
    .B1(net682),
    .A1(net789),
    .Y(_0586_),
    .A2(net683));
 sg13g2_o21ai_1 _3042_ (.B1(_0586_),
    .VDD(VPWR),
    .Y(_0587_),
    .VSS(VGND),
    .A1(_0582_),
    .A2(_0583_));
 sg13g2_nor3_1 _3043_ (.A(_0578_),
    .B(_0579_),
    .C(_0587_),
    .Y(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3044_ (.A(_1945_),
    .B_N(_0203_),
    .Y(_0589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3045_ (.B1(_0589_),
    .VDD(VPWR),
    .Y(_0590_),
    .VSS(VGND),
    .A1(_0574_),
    .A2(_0575_));
 sg13g2_nand2b_1 _3046_ (.Y(_0591_),
    .B(\sap_3_inst.alu.carry ),
    .A_N(_0589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3047_ (.B1(_0591_),
    .VDD(VPWR),
    .Y(_0049_),
    .VSS(VGND),
    .A1(_0588_),
    .A2(_0590_));
 sg13g2_nor3_1 _3048_ (.A(net736),
    .B(_1553_),
    .C(_1732_),
    .Y(_0592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3049_ (.Y(_0593_),
    .B1(_1849_),
    .B2(_0592_),
    .A2(_1780_),
    .A1(net736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3050_ (.A0(\sap_3_inst.alu.tmp[0] ),
    .A1(net31),
    .S(net715),
    .X(_0050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3051_ (.A(\sap_3_inst.alu.tmp[1] ),
    .B(net715),
    .Y(_0594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3052_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0227_),
    .A2(net715),
    .Y(_0051_),
    .B1(_0594_));
 sg13g2_nand2_1 _3053_ (.Y(_0595_),
    .A(net19),
    .B(net715),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3054_ (.B1(_0595_),
    .VDD(VPWR),
    .Y(_0052_),
    .VSS(VGND),
    .A1(_1471_),
    .A2(net715));
 sg13g2_nor2_1 _3055_ (.A(\sap_3_inst.alu.tmp[3] ),
    .B(net715),
    .Y(_0596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3056_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net572),
    .A2(net716),
    .Y(_0053_),
    .B1(_0596_));
 sg13g2_nand2_1 _3057_ (.Y(_0597_),
    .A(net32),
    .B(net716),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3058_ (.B1(_0597_),
    .VDD(VPWR),
    .Y(_0054_),
    .VSS(VGND),
    .A1(_1473_),
    .A2(net716));
 sg13g2_mux2_1 _3059_ (.A0(\sap_3_inst.alu.tmp[5] ),
    .A1(net22),
    .S(net715),
    .X(_0055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3060_ (.A0(\sap_3_inst.alu.tmp[6] ),
    .A1(net23),
    .S(net715),
    .X(_0056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3061_ (.A0(\sap_3_inst.alu.tmp[7] ),
    .A1(net24),
    .S(net716),
    .X(_0057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3062_ (.A0(net31),
    .A1(net785),
    .S(net738),
    .X(_0058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3063_ (.Y(_0598_),
    .A(net782),
    .B(net739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3064_ (.B1(_0598_),
    .VDD(VPWR),
    .Y(_0059_),
    .VSS(VGND),
    .A1(net739),
    .A2(_0227_));
 sg13g2_nor2_1 _3065_ (.A(net738),
    .B(net19),
    .Y(_0599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3066_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1444_),
    .A2(net738),
    .Y(_0060_),
    .B1(_0599_));
 sg13g2_nand2_1 _3067_ (.Y(_0600_),
    .A(net776),
    .B(net739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3068_ (.B1(_0600_),
    .VDD(VPWR),
    .Y(_0061_),
    .VSS(VGND),
    .A1(net738),
    .A2(net572));
 sg13g2_nor2_1 _3069_ (.A(net738),
    .B(net32),
    .Y(_0601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3070_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1442_),
    .A2(net738),
    .Y(_0062_),
    .B1(_0601_));
 sg13g2_mux2_1 _3071_ (.A0(net22),
    .A1(net772),
    .S(net738),
    .X(_0063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3072_ (.A0(net33),
    .A1(net770),
    .S(net738),
    .X(_0064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3073_ (.A(net739),
    .B(net34),
    .Y(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3074_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1443_),
    .A2(net739),
    .Y(_0065_),
    .B1(_0602_));
 sg13g2_a21oi_1 _3075_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1615_),
    .A2(_1749_),
    .Y(_0603_),
    .B1(net731));
 sg13g2_nand2b_1 _3076_ (.Y(_0604_),
    .B(_1851_),
    .A_N(_1746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3077_ (.B1(_0604_),
    .VDD(VPWR),
    .Y(_0605_),
    .VSS(VGND),
    .A1(_1594_),
    .A2(_1850_));
 sg13g2_a22oi_1 _3078_ (.Y(_0606_),
    .B1(_1642_),
    .B2(_1532_),
    .A2(net747),
    .A1(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3079_ (.B(net752),
    .C(net777),
    .Y(_0607_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0606_));
 sg13g2_o21ai_1 _3080_ (.B1(_0607_),
    .VDD(VPWR),
    .Y(_0608_),
    .VSS(VGND),
    .A1(_1588_),
    .A2(_1748_));
 sg13g2_o21ai_1 _3081_ (.B1(net752),
    .VDD(VPWR),
    .Y(_0609_),
    .VSS(VGND),
    .A1(_1576_),
    .A2(_1656_));
 sg13g2_a21oi_1 _3082_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net731),
    .A2(_1657_),
    .Y(_0610_),
    .B1(_1596_));
 sg13g2_a21o_1 _3083_ (.A2(_1645_),
    .A1(net733),
    .B1(_1605_),
    .X(_0611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3084_ (.B(_1549_),
    .C(net735),
    .A(net773),
    .Y(_0612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3085_ (.B(_0609_),
    .C(_0611_),
    .A(_1770_),
    .Y(_0613_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0612_));
 sg13g2_nor4_1 _3086_ (.A(_0603_),
    .B(_0605_),
    .C(_0608_),
    .D(_0613_),
    .Y(_0614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3087_ (.A(net741),
    .B(_1594_),
    .Y(_0615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3088_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net725),
    .A2(_0615_),
    .Y(_0616_),
    .B1(_1516_));
 sg13g2_o21ai_1 _3089_ (.B1(_0616_),
    .VDD(VPWR),
    .Y(_0617_),
    .VSS(VGND),
    .A1(net724),
    .A2(_0614_));
 sg13g2_a21oi_1 _3090_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1516_),
    .A2(_1746_),
    .Y(_0618_),
    .B1(_1842_));
 sg13g2_and2_1 _3091_ (.A(_0617_),
    .B(_0618_),
    .X(_0619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3092_ (.A(_1442_),
    .B(net773),
    .C(_1570_),
    .D(net731),
    .Y(_0620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3093_ (.A(_1570_),
    .B(net726),
    .Y(_0621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3094_ (.A(_1573_),
    .B(_1575_),
    .Y(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3095_ (.A(_0620_),
    .B(_0621_),
    .C(_0622_),
    .X(_0623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3096_ (.X(_0624_),
    .A(_1607_),
    .B(_1622_),
    .C(_0623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3097_ (.A(net731),
    .B(_1598_),
    .Y(_0625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3098_ (.Y(_0626_),
    .B1(_1702_),
    .B2(net731),
    .A2(_1619_),
    .A1(_1582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3099_ (.Y(_0627_),
    .A(_1577_),
    .B(_1654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3100_ (.Y(_0628_),
    .B(_1638_),
    .A_N(net753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3101_ (.Y(_0629_),
    .A(_1716_),
    .B(_1851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3102_ (.A2(_0629_),
    .A1(_0628_),
    .B1(_1442_),
    .X(_0630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3103_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1611_),
    .C1(_0610_),
    .B1(_0627_),
    .A1(net775),
    .Y(_0631_),
    .A2(_1823_));
 sg13g2_a21oi_1 _3104_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1576_),
    .A2(_1753_),
    .Y(_0632_),
    .B1(_0626_));
 sg13g2_nor4_1 _3105_ (.A(net725),
    .B(_1769_),
    .C(_1828_),
    .D(_0625_),
    .Y(_0633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3106_ (.B(_0631_),
    .C(_0632_),
    .A(_0630_),
    .Y(_0634_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0633_));
 sg13g2_and2_1 _3107_ (.A(net743),
    .B(_1711_),
    .X(_0635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3108_ (.Y(_0636_),
    .A(net743),
    .B(_1711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3109_ (.A(net741),
    .B(_1515_),
    .C(_1715_),
    .Y(_0637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3110_ (.B1(net774),
    .VDD(VPWR),
    .Y(_0638_),
    .VSS(VGND),
    .A1(_0635_),
    .A2(_0637_));
 sg13g2_a21oi_1 _3111_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net725),
    .A2(_0638_),
    .Y(_0639_),
    .B1(_1520_));
 sg13g2_o21ai_1 _3112_ (.B1(_0639_),
    .VDD(VPWR),
    .Y(_0640_),
    .VSS(VGND),
    .A1(_0624_),
    .A2(_0634_));
 sg13g2_o21ai_1 _3113_ (.B1(_1530_),
    .VDD(VPWR),
    .Y(_0641_),
    .VSS(VGND),
    .A1(\sap_3_inst.controller.stage[1] ),
    .A2(_1506_));
 sg13g2_nand3_1 _3114_ (.B(net729),
    .C(_1716_),
    .A(\sap_3_inst.controller.opcode[4] ),
    .Y(_0642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3115_ (.A2(_0642_),
    .A1(_1516_),
    .B1(_0641_),
    .X(_0643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3116_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0643_),
    .Y(_0644_),
    .A2(_0640_),
    .A1(net757));
 sg13g2_a21o_1 _3117_ (.A2(_0640_),
    .A1(net757),
    .B1(_0643_),
    .X(_0645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3118_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0646_),
    .B(_1792_),
    .A(_1441_));
 sg13g2_a22oi_1 _3119_ (.Y(_0647_),
    .B1(net727),
    .B2(_0646_),
    .A2(_1615_),
    .A1(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3120_ (.B(net745),
    .C(_1514_),
    .A(net778),
    .Y(_0648_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net764));
 sg13g2_nor4_1 _3121_ (.A(_1512_),
    .B(_1591_),
    .C(_1593_),
    .D(net727),
    .Y(_0649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3122_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net777),
    .C1(_0649_),
    .B1(_1823_),
    .A1(_1571_),
    .Y(_0650_),
    .A2(_1604_));
 sg13g2_o21ai_1 _3123_ (.B1(_1588_),
    .VDD(VPWR),
    .Y(_0651_),
    .VSS(VGND),
    .A1(net765),
    .A2(_1570_));
 sg13g2_a22oi_1 _3124_ (.Y(_0652_),
    .B1(_0651_),
    .B2(net728),
    .A2(_1685_),
    .A1(_1621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3125_ (.B(_0650_),
    .C(_0652_),
    .A(_0648_),
    .Y(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3126_ (.B1(net757),
    .VDD(VPWR),
    .Y(_0654_),
    .VSS(VGND),
    .A1(_0647_),
    .A2(_0653_));
 sg13g2_nor3_1 _3127_ (.A(net769),
    .B(net767),
    .C(_1518_),
    .Y(_0655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3128_ (.B(net729),
    .C(_0655_),
    .A(net778),
    .Y(_0656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3129_ (.A(_0654_),
    .B(_0656_),
    .X(_0657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3130_ (.Y(_0658_),
    .A(_0654_),
    .B(_0656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3131_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0656_),
    .C1(_0643_),
    .B1(_0654_),
    .A1(net757),
    .Y(_0659_),
    .A2(_0640_));
 sg13g2_and2_1 _3132_ (.A(net706),
    .B(net690),
    .X(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3133_ (.Y(_0661_),
    .A(net704),
    .B(net690),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3134_ (.A(net702),
    .B(net691),
    .Y(_0662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3135_ (.X(_0663_),
    .A(net703),
    .B(net697),
    .C(net692),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3136_ (.Y(_0664_),
    .A(net705),
    .B(_0662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3137_ (.X(_0665_),
    .A(net705),
    .B(net699),
    .C(_0658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3138_ (.VDD(VPWR),
    .Y(_0666_),
    .A(net676),
    .VSS(VGND));
 sg13g2_nand3b_1 _3139_ (.B(_1787_),
    .C(net719),
    .Y(_0667_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0621_));
 sg13g2_nor2_1 _3140_ (.A(_0622_),
    .B(_0667_),
    .Y(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3141_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1623_),
    .A2(_0668_),
    .Y(_0669_),
    .B1(_0275_));
 sg13g2_and2_1 _3142_ (.A(net742),
    .B(net726),
    .X(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3143_ (.A(_1536_),
    .B(_1642_),
    .X(_0671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3144_ (.B1(_1608_),
    .VDD(VPWR),
    .Y(_0672_),
    .VSS(VGND),
    .A1(_1632_),
    .A2(_0671_));
 sg13g2_a22oi_1 _3145_ (.Y(_0673_),
    .B1(_0670_),
    .B2(_0672_),
    .A2(_1614_),
    .A1(_1609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3146_ (.Y(_0674_),
    .B1(net730),
    .B2(net726),
    .A2(_1620_),
    .A1(net749),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3147_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1630_),
    .C1(_0674_),
    .B1(_0673_),
    .A1(net750),
    .Y(_0675_),
    .A2(_0671_));
 sg13g2_a21oi_1 _3148_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net735),
    .A2(_1616_),
    .Y(_0676_),
    .B1(_1597_));
 sg13g2_nand2_1 _3149_ (.Y(_0677_),
    .A(_1587_),
    .B(_0676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3150_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1587_),
    .A2(_0676_),
    .Y(_0678_),
    .B1(net726));
 sg13g2_nand2b_1 _3151_ (.Y(_0679_),
    .B(net752),
    .A_N(net726),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3152_ (.A(net764),
    .B(net753),
    .C(_1639_),
    .X(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3153_ (.A2(net730),
    .A1(net734),
    .B1(net753),
    .X(_0681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3154_ (.B(_0679_),
    .C(_0680_),
    .A(_1787_),
    .Y(_0682_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0681_));
 sg13g2_a221oi_1 _3155_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0677_),
    .C1(_0682_),
    .B1(_1703_),
    .A1(_1607_),
    .Y(_0683_),
    .A2(_1622_));
 sg13g2_a221oi_1 _3156_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0683_),
    .C1(_0275_),
    .B1(_0675_),
    .A1(_1623_),
    .Y(_0684_),
    .A2(_0668_));
 sg13g2_nand2_2 _3157_ (.Y(_0685_),
    .A(_1535_),
    .B(_0636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3158_ (.Y(_0686_),
    .A(net764),
    .B(_1535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3159_ (.A2(_0686_),
    .A1(_0685_),
    .B1(_0684_),
    .X(_0687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3160_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0686_),
    .C1(_0684_),
    .B1(_0685_),
    .A1(_0617_),
    .Y(_0688_),
    .A2(_0618_));
 sg13g2_and2_1 _3161_ (.A(_0659_),
    .B(net686),
    .X(_0689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3162_ (.Y(_0690_),
    .A(net690),
    .B(net686),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3163_ (.Y(_0691_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .B(net674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3164_ (.A(net704),
    .B(net702),
    .C(_0658_),
    .D(net689),
    .Y(_0692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3165_ (.Y(_0693_),
    .A(_0662_),
    .B(net686),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3166_ (.A(net700),
    .B(net691),
    .Y(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3167_ (.A(net705),
    .B(net699),
    .C(_0658_),
    .Y(_0695_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net689));
 sg13g2_nand2_1 _3168_ (.Y(_0696_),
    .A(net687),
    .B(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3169_ (.X(_0697_),
    .A(net703),
    .B(net701),
    .C(net692),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3170_ (.Y(_0698_),
    .A(net706),
    .B(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3171_ (.A(net704),
    .B(net701),
    .C(net693),
    .D(net688),
    .Y(_0699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3172_ (.B(net691),
    .C(net687),
    .A(net697),
    .Y(_0700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3173_ (.Y(_0701_),
    .B1(net664),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .A2(net665),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3174_ (.X(_0702_),
    .A(net700),
    .B(net693),
    .C(net688),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3175_ (.Y(_0703_),
    .A(_0662_),
    .B(net688),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3176_ (.X(_0704_),
    .A(net701),
    .B(net693),
    .C(net688),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3177_ (.Y(_0705_),
    .A(net688),
    .B(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3178_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .C1(net671),
    .B1(net662),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .Y(_0706_),
    .A2(net676));
 sg13g2_a22oi_1 _3179_ (.Y(_0707_),
    .B1(net657),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ),
    .A2(net681),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3180_ (.Y(_0708_),
    .B1(net667),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .A2(net678),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3181_ (.A(_0691_),
    .B(_0701_),
    .C(_0707_),
    .D(_0708_),
    .X(_0709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3182_ (.Y(_0710_),
    .B1(_0706_),
    .B2(_0709_),
    .A2(net672),
    .A1(_1468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3183_ (.Y(_0711_),
    .A(_0710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3184_ (.Y(_0712_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .B(net678),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3185_ (.Y(_0713_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .B(net675),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3186_ (.Y(_0714_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .B(net663),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3187_ (.B1(_0712_),
    .VDD(VPWR),
    .Y(_0715_),
    .VSS(VGND),
    .A1(_1497_),
    .A2(_0666_));
 sg13g2_a22oi_1 _3188_ (.Y(_0716_),
    .B1(net666),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .A2(net672),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3189_ (.B1(_0714_),
    .VDD(VPWR),
    .Y(_0717_),
    .VSS(VGND),
    .A1(_1499_),
    .A2(net620));
 sg13g2_o21ai_1 _3190_ (.B1(_0713_),
    .VDD(VPWR),
    .Y(_0718_),
    .VSS(VGND),
    .A1(_1495_),
    .A2(net613));
 sg13g2_a22oi_1 _3191_ (.Y(_0719_),
    .B1(net658),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .A2(net680),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3192_ (.Y(_0720_),
    .A(_0716_),
    .B(_0719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3193_ (.A(_0715_),
    .B(_0717_),
    .C(_0718_),
    .Y(_0721_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0720_));
 sg13g2_or4_1 _3194_ (.A(_0715_),
    .B(_0717_),
    .C(_0718_),
    .D(_0720_),
    .X(_0722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3195_ (.Y(_0723_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .B(net680),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3196_ (.B1(_0723_),
    .VDD(VPWR),
    .Y(_0724_),
    .VSS(VGND),
    .A1(_1491_),
    .A2(net619));
 sg13g2_nand2_1 _3197_ (.Y(_0725_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .B(net674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3198_ (.Y(_0726_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .B(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3199_ (.B1(_0725_),
    .VDD(VPWR),
    .Y(_0727_),
    .VSS(VGND),
    .A1(_1488_),
    .A2(net617));
 sg13g2_a22oi_1 _3200_ (.Y(_0728_),
    .B1(net655),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .A2(net664),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3201_ (.B1(_0726_),
    .VDD(VPWR),
    .Y(_0729_),
    .VSS(VGND),
    .A1(_1486_),
    .A2(net612));
 sg13g2_a22oi_1 _3202_ (.Y(_0730_),
    .B1(net677),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .A2(net679),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3203_ (.Y(_0731_),
    .A(_0728_),
    .B(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3204_ (.A(_0724_),
    .B(_0727_),
    .C(_0729_),
    .Y(_0732_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0731_));
 sg13g2_or4_1 _3205_ (.A(_0724_),
    .B(_0727_),
    .C(_0729_),
    .D(_0731_),
    .X(_0733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3206_ (.Y(_0734_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .B(net674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3207_ (.Y(_0735_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .B(net677),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3208_ (.Y(_0736_),
    .B1(net656),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .A2(net663),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3209_ (.Y(_0737_),
    .B1(net668),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .A2(net670),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3210_ (.Y(_0738_),
    .B1(net665),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ),
    .A2(net679),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3211_ (.Y(_0739_),
    .B1(net660),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .A2(net680),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3212_ (.X(_0740_),
    .A(_0736_),
    .B(_0737_),
    .C(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3213_ (.A(_0734_),
    .B(_0735_),
    .C(_0738_),
    .D(_0740_),
    .X(_0741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3214_ (.B(_0735_),
    .C(_0738_),
    .A(_0734_),
    .Y(_0742_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0740_));
 sg13g2_nand4_1 _3215_ (.B(net698),
    .C(net691),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .Y(_0743_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net686));
 sg13g2_nand4_1 _3216_ (.B(net704),
    .C(net698),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .Y(_0744_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net694));
 sg13g2_nand4_1 _3217_ (.B(net701),
    .C(net696),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .Y(_0745_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net686));
 sg13g2_nand4_1 _3218_ (.B(net704),
    .C(net701),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .Y(_0746_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net694));
 sg13g2_nand4_1 _3219_ (.B(net698),
    .C(net694),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .Y(_0747_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net686));
 sg13g2_nor2_1 _3220_ (.A(_1479_),
    .B(_0690_),
    .Y(_0748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3221_ (.B(net701),
    .C(net694),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .Y(_0749_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net689));
 sg13g2_nand4_1 _3222_ (.B(net704),
    .C(net698),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .Y(_0750_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net691));
 sg13g2_nand4_1 _3223_ (.B(net698),
    .C(net694),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .Y(_0751_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net689));
 sg13g2_nand4_1 _3224_ (.B(_0746_),
    .C(_0747_),
    .A(_0744_),
    .Y(_0752_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0750_));
 sg13g2_o21ai_1 _3225_ (.B1(_0745_),
    .VDD(VPWR),
    .Y(_0753_),
    .VSS(VGND),
    .A1(_1477_),
    .A2(_0661_));
 sg13g2_nand3_1 _3226_ (.B(_0749_),
    .C(_0751_),
    .A(_0743_),
    .Y(_0754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3227_ (.A(_0748_),
    .B(_0752_),
    .C(_0753_),
    .Y(_0755_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0754_));
 sg13g2_or4_1 _3228_ (.A(_0748_),
    .B(_0752_),
    .C(_0753_),
    .D(_0754_),
    .X(_0756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3229_ (.B(net703),
    .C(net697),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .Y(_0757_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net692));
 sg13g2_nand4_1 _3230_ (.B(net701),
    .C(net692),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .Y(_0758_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net687));
 sg13g2_and3_1 _3231_ (.X(_0759_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .B(net690),
    .C(net687),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3232_ (.B(net703),
    .C(net690),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .Y(_0760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3233_ (.Y(_0761_),
    .B1(net666),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ),
    .A2(net671),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3234_ (.Y(_0762_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .B(net676),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3235_ (.B(net697),
    .C(net691),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ),
    .Y(_0763_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net687));
 sg13g2_and4_1 _3236_ (.A(_0757_),
    .B(_0758_),
    .C(_0760_),
    .D(_0763_),
    .X(_0764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3237_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .C1(_0759_),
    .B1(net657),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .Y(_0765_),
    .A2(net661));
 sg13g2_and4_1 _3238_ (.A(_0761_),
    .B(_0762_),
    .C(_0764_),
    .D(_0765_),
    .X(_0766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3239_ (.B(net697),
    .C(net692),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ),
    .Y(_0767_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net688));
 sg13g2_nand3_1 _3240_ (.B(net703),
    .C(net690),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .Y(_0768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3241_ (.B(net701),
    .C(net692),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .Y(_0769_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net688));
 sg13g2_nand4_1 _3242_ (.B(net703),
    .C(net700),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .Y(_0770_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net693));
 sg13g2_a22oi_1 _3243_ (.Y(_0771_),
    .B1(net663),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .A2(net676),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3244_ (.Y(_0772_),
    .B1(net666),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ),
    .A2(net674),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3245_ (.Y(_0773_),
    .B1(net667),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ),
    .A2(net671),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3246_ (.A(_0767_),
    .B(_0768_),
    .C(_0769_),
    .D(_0770_),
    .X(_0774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3247_ (.A(_0771_),
    .B(_0772_),
    .C(_0773_),
    .D(_0774_),
    .X(_0775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3248_ (.B(net704),
    .C(net702),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .Y(_0776_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net694));
 sg13g2_o21ai_1 _3249_ (.B1(_0776_),
    .VDD(VPWR),
    .Y(_0777_),
    .VSS(VGND),
    .A1(_1470_),
    .A2(_0690_));
 sg13g2_nand3_1 _3250_ (.B(net705),
    .C(_0659_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .Y(_0778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3251_ (.B(net702),
    .C(net694),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .Y(_0779_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0688_));
 sg13g2_nand4_1 _3252_ (.B(net698),
    .C(net694),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .Y(_0780_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net689));
 sg13g2_nand4_1 _3253_ (.B(net702),
    .C(net695),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .Y(_0781_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net689));
 sg13g2_nand4_1 _3254_ (.B(net698),
    .C(net695),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .Y(_0782_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net686));
 sg13g2_nand4_1 _3255_ (.B(net704),
    .C(net698),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .Y(_0783_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net695));
 sg13g2_nand4_1 _3256_ (.B(net699),
    .C(net691),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .Y(_0784_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net686));
 sg13g2_and2_1 _3257_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .B(net676),
    .X(_0785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3258_ (.B(_0782_),
    .C(_0784_),
    .A(_0778_),
    .Y(_0786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3259_ (.B(_0780_),
    .C(_0781_),
    .A(_0779_),
    .Y(_0787_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0783_));
 sg13g2_nor4_1 _3260_ (.A(_0777_),
    .B(_0785_),
    .C(_0786_),
    .D(_0787_),
    .Y(_0788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _3261_ (.A(_0777_),
    .B(_0785_),
    .C(_0786_),
    .D(_0787_),
    .X(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3262_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .B(net697),
    .C(net692),
    .D(net687),
    .X(_0790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3263_ (.Y(_0791_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .B(net663),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3264_ (.B(net690),
    .C(net687),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .Y(_0792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3265_ (.B(net703),
    .C(net690),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .Y(_0793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3266_ (.B(net703),
    .C(net697),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .Y(_0794_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net691));
 sg13g2_nand4_1 _3267_ (.B(net697),
    .C(net692),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .Y(_0795_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net688));
 sg13g2_a22oi_1 _3268_ (.Y(_0796_),
    .B1(net665),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .A2(net668),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3269_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .C1(_0790_),
    .B1(net655),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .Y(_0797_),
    .A2(net679));
 sg13g2_and4_1 _3270_ (.A(_0792_),
    .B(_0793_),
    .C(_0794_),
    .D(_0795_),
    .X(_0798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3271_ (.A(_0791_),
    .B(_0796_),
    .C(_0797_),
    .D(_0798_),
    .X(_0799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3272_ (.A(_0775_),
    .B(net588),
    .X(_0800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3273_ (.Y(_0801_),
    .A(_0775_),
    .B(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3274_ (.A(_0766_),
    .B(_0775_),
    .C(net591),
    .D(net588),
    .X(_0802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3275_ (.A(_0755_),
    .B(_0802_),
    .X(_0803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3276_ (.Y(_0804_),
    .A(_0741_),
    .B(_0803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3277_ (.B(_0741_),
    .C(_0755_),
    .A(_0732_),
    .Y(_0805_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0802_));
 sg13g2_nor2_1 _3278_ (.A(_0722_),
    .B(_0805_),
    .Y(_0806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3279_ (.Y(_0807_),
    .A(_0711_),
    .B(_0806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3280_ (.Y(_0808_),
    .A(_0711_),
    .B(_0806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3281_ (.Y(_0809_),
    .A(_1608_),
    .B(_1630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3282_ (.B1(net735),
    .VDD(VPWR),
    .Y(_0810_),
    .VSS(VGND),
    .A1(_1586_),
    .A2(_1613_));
 sg13g2_a21o_1 _3283_ (.A2(_0810_),
    .A1(_0809_),
    .B1(_0670_),
    .X(_0811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3284_ (.B(_1620_),
    .C(_0676_),
    .A(net749),
    .Y(_0812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3285_ (.A(net751),
    .B(_1687_),
    .Y(_0813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3286_ (.B1(_0681_),
    .VDD(VPWR),
    .Y(_0814_),
    .VSS(VGND),
    .A1(net751),
    .A2(_1687_));
 sg13g2_or2_1 _3287_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0815_),
    .B(_0814_),
    .A(_0667_));
 sg13g2_nand2_1 _3288_ (.Y(_0816_),
    .A(_1613_),
    .B(_1697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3289_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0812_),
    .C1(_0815_),
    .B1(_1703_),
    .A1(_1613_),
    .Y(_0817_),
    .A2(_1697_));
 sg13g2_a21oi_1 _3290_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0811_),
    .A2(_0817_),
    .Y(_0818_),
    .B1(_0275_));
 sg13g2_o21ai_1 _3291_ (.B1(_1535_),
    .VDD(VPWR),
    .Y(_0819_),
    .VSS(VGND),
    .A1(net776),
    .A2(_0636_));
 sg13g2_nor2_2 _3292_ (.A(_0818_),
    .B(_0819_),
    .Y(_0820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3293_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0821_),
    .B(_0819_),
    .A(_0818_));
 sg13g2_a21o_1 _3294_ (.A2(_1654_),
    .A1(net742),
    .B1(_0809_),
    .X(_0822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3295_ (.Y(_0823_),
    .A(net750),
    .B(_1654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3296_ (.B1(_0823_),
    .VDD(VPWR),
    .Y(_0824_),
    .VSS(VGND),
    .A1(net750),
    .A2(_0622_));
 sg13g2_nand3_1 _3297_ (.B(net743),
    .C(_1711_),
    .A(net776),
    .Y(_0825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3298_ (.A(_0816_),
    .B(_0822_),
    .C(_0824_),
    .D(_0825_),
    .X(_0826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3299_ (.B(_0822_),
    .C(_0824_),
    .A(_0816_),
    .Y(_0827_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0825_));
 sg13g2_nor2_2 _3300_ (.A(net651),
    .B(net712),
    .Y(_0828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3301_ (.Y(_0829_),
    .A(net653),
    .B(net711),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3302_ (.Y(_0830_),
    .A(_0808_),
    .B(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3303_ (.Y(_0831_),
    .A(net776),
    .B(_0635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3304_ (.B(_0822_),
    .C(_0824_),
    .A(_0816_),
    .Y(_0832_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0831_));
 sg13g2_nor2_1 _3305_ (.A(net653),
    .B(net711),
    .Y(_0833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3306_ (.Y(_0834_),
    .A(net651),
    .B(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3307_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0835_),
    .B(net589),
    .A(_0775_));
 sg13g2_nor2_1 _3308_ (.A(_0766_),
    .B(_0835_),
    .Y(_0836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3309_ (.A(_0755_),
    .B(_0766_),
    .C(_0775_),
    .Y(_0837_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net589));
 sg13g2_or4_1 _3310_ (.A(_0755_),
    .B(_0766_),
    .C(_0775_),
    .D(net588),
    .X(_0838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3311_ (.Y(_0839_),
    .A(_0742_),
    .B(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3312_ (.B(_0742_),
    .C(_0837_),
    .A(_0733_),
    .Y(_0840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3313_ (.A(_0721_),
    .B(_0732_),
    .C(_0741_),
    .D(_0838_),
    .Y(_0841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3314_ (.B(_0733_),
    .C(_0742_),
    .A(_0722_),
    .Y(_0842_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0837_));
 sg13g2_nand2_1 _3315_ (.Y(_0843_),
    .A(_0710_),
    .B(_0841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3316_ (.Y(_0844_),
    .A(net590),
    .B(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3317_ (.A(net591),
    .B(_0839_),
    .Y(_0845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3318_ (.A(net591),
    .B(_0842_),
    .Y(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3319_ (.Y(_0847_),
    .A(_0710_),
    .B(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3320_ (.A(net599),
    .B(_0847_),
    .Y(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3321_ (.A(net651),
    .B(net711),
    .Y(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3322_ (.Y(_0850_),
    .A(net653),
    .B(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3323_ (.B(net729),
    .C(_1716_),
    .A(_1516_),
    .Y(_0851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3324_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1577_),
    .A2(net730),
    .Y(_0852_),
    .B1(_1620_));
 sg13g2_a21oi_1 _3325_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1643_),
    .A2(net727),
    .Y(_0853_),
    .B1(_1610_));
 sg13g2_o21ai_1 _3326_ (.B1(_0629_),
    .VDD(VPWR),
    .Y(_0854_),
    .VSS(VGND),
    .A1(net765),
    .A2(_1850_));
 sg13g2_nand2_1 _3327_ (.Y(_0855_),
    .A(_1551_),
    .B(_0611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3328_ (.B1(_1753_),
    .VDD(VPWR),
    .Y(_0856_),
    .VSS(VGND),
    .A1(_1576_),
    .A2(_1638_));
 sg13g2_nor3_1 _3329_ (.A(_1847_),
    .B(_0852_),
    .C(_0853_),
    .Y(_0857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3330_ (.A(_1769_),
    .B(_0625_),
    .C(_0854_),
    .D(_0855_),
    .Y(_0858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3331_ (.B(_0857_),
    .C(_0858_),
    .A(_0856_),
    .Y(_0859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3332_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0312_),
    .A2(_0859_),
    .Y(_0860_),
    .B1(_0637_));
 sg13g2_o21ai_1 _3333_ (.B1(_0851_),
    .VDD(VPWR),
    .Y(_0861_),
    .VSS(VGND),
    .A1(_0280_),
    .A2(_0860_));
 sg13g2_nand2b_2 _3334_ (.Y(_0862_),
    .B(_0861_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0641_));
 sg13g2_a21o_1 _3335_ (.A2(_0862_),
    .A1(net597),
    .B1(net621),
    .X(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3336_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net730),
    .A2(net726),
    .Y(_0864_),
    .B1(net753));
 sg13g2_nor4_1 _3337_ (.A(_0266_),
    .B(_0678_),
    .C(_0813_),
    .D(_0864_),
    .Y(_0865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3338_ (.B(_0675_),
    .C(_0865_),
    .A(_1624_),
    .Y(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3339_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0669_),
    .A2(_0866_),
    .Y(_0867_),
    .B1(_0685_));
 sg13g2_nand2b_1 _3340_ (.Y(_0868_),
    .B(net673),
    .A_N(net684),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3341_ (.Y(_0869_),
    .A(net597),
    .B(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3342_ (.A0(net9),
    .A1(net31),
    .S(net596),
    .X(_0870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3343_ (.A(_0848_),
    .B(net587),
    .C(_0870_),
    .Y(_0871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3344_ (.A(net653),
    .B(net712),
    .Y(_0872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3345_ (.Y(_0873_),
    .A(net652),
    .B(_0827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3346_ (.B1(net598),
    .VDD(VPWR),
    .Y(_0874_),
    .VSS(VGND),
    .A1(net592),
    .A2(net654));
 sg13g2_a22oi_1 _3347_ (.Y(_0066_),
    .B1(_0871_),
    .B2(_0830_),
    .A2(net587),
    .A1(_1468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3348_ (.Y(_0875_),
    .B1(net660),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .A2(net668),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3349_ (.Y(_0876_),
    .B1(net677),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .A2(net679),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3350_ (.B1(_0876_),
    .VDD(VPWR),
    .Y(_0877_),
    .VSS(VGND),
    .A1(_1467_),
    .A2(_0700_));
 sg13g2_a22oi_1 _3351_ (.Y(_0878_),
    .B1(net665),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .A2(net680),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3352_ (.Y(_0879_),
    .B1(net655),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ),
    .A2(net674),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3353_ (.B(_0875_),
    .C(_0878_),
    .A(net621),
    .Y(_0880_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0879_));
 sg13g2_nor2_1 _3354_ (.A(_0877_),
    .B(_0880_),
    .Y(_0881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3355_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[0][1] ),
    .B(net621),
    .Y(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3356_ (.A(_0881_),
    .B(_0882_),
    .Y(_0883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3357_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0884_),
    .B(_0882_),
    .A(_0881_));
 sg13g2_nor4_2 _3358_ (.A(_0710_),
    .B(_0722_),
    .C(_0805_),
    .Y(_0885_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0883_));
 sg13g2_xnor2_1 _3359_ (.Y(_0886_),
    .A(_0807_),
    .B(_0884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3360_ (.A(net606),
    .B(_0886_),
    .X(_0887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3361_ (.B(_0841_),
    .C(_0883_),
    .A(_0710_),
    .Y(_0888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3362_ (.A(net591),
    .B(_0888_),
    .Y(_0889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3363_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0710_),
    .A2(_0846_),
    .Y(_0890_),
    .B1(_0883_));
 sg13g2_nor2_1 _3364_ (.A(_0889_),
    .B(_0890_),
    .Y(_0891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3365_ (.A(net599),
    .B(_0891_),
    .Y(_0892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3366_ (.Y(_0893_),
    .B(net597),
    .A_N(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3367_ (.Y(_0894_),
    .B1(_0869_),
    .B2(_0893_),
    .A2(net595),
    .A1(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3368_ (.A(net586),
    .B(_0887_),
    .C(_0892_),
    .D(_0894_),
    .Y(_0895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3369_ (.Y(_0896_),
    .A(_0843_),
    .B(_0883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3370_ (.A(net591),
    .B(net589),
    .Y(_0897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3371_ (.Y(_0898_),
    .A(net590),
    .B(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3372_ (.A2(net586),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[0][1] ),
    .B1(_0895_),
    .X(_0067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3373_ (.Y(_0899_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][2] ),
    .B(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3374_ (.Y(_0900_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ),
    .B(net675),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3375_ (.Y(_0901_),
    .B1(net661),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .A2(net676),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3376_ (.Y(_0902_),
    .B1(net663),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .A2(net666),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3377_ (.Y(_0903_),
    .B1(net657),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .A2(net667),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3378_ (.Y(_0904_),
    .B1(net678),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .A2(net680),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3379_ (.A(_0900_),
    .B(_0902_),
    .C(_0903_),
    .D(_0904_),
    .X(_0905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3380_ (.B(_0901_),
    .C(_0905_),
    .A(net622),
    .Y(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3381_ (.B1(_0906_),
    .VDD(VPWR),
    .Y(_0907_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[0][2] ),
    .A2(net622));
 sg13g2_nor4_2 _3382_ (.A(_0711_),
    .B(_0842_),
    .C(_0884_),
    .Y(_0908_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0907_));
 sg13g2_xor2_1 _3383_ (.B(_0907_),
    .A(_0889_),
    .X(_0909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3384_ (.Y(_0910_),
    .A(net600),
    .B(_0909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3385_ (.Y(_0911_),
    .A(_0775_),
    .B(_0897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3386_ (.Y(_0912_),
    .B(_0910_),
    .A_N(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3387_ (.Y(_0913_),
    .A(_0885_),
    .B(_0907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3388_ (.B(_0907_),
    .A(_0885_),
    .X(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3389_ (.Y(_0915_),
    .A(net19),
    .B(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3390_ (.B1(_0869_),
    .VDD(VPWR),
    .Y(_0916_),
    .VSS(VGND),
    .A1(net11),
    .A2(_0850_));
 sg13g2_a221oi_1 _3391_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0916_),
    .C1(_0872_),
    .B1(_0915_),
    .A1(net711),
    .Y(_0917_),
    .A2(_0914_));
 sg13g2_nor2_1 _3392_ (.A(_0800_),
    .B(_0873_),
    .Y(_0918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3393_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0835_),
    .A2(_0918_),
    .Y(_0919_),
    .B1(_0917_));
 sg13g2_a21o_1 _3394_ (.A2(net589),
    .A1(net591),
    .B1(_0775_),
    .X(_0920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3395_ (.B1(_0920_),
    .VDD(VPWR),
    .Y(_0921_),
    .VSS(VGND),
    .A1(net590),
    .A2(_0801_));
 sg13g2_and4_1 _3396_ (.A(_0801_),
    .B(net651),
    .C(_0832_),
    .D(_0835_),
    .X(_0922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3397_ (.B1(_0899_),
    .VDD(VPWR),
    .Y(_0068_),
    .VSS(VGND),
    .A1(_0912_),
    .A2(_0919_));
 sg13g2_a22oi_1 _3398_ (.Y(_0923_),
    .B1(net661),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .A2(net663),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3399_ (.Y(_0924_),
    .B1(net666),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .A2(net676),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3400_ (.A(_0923_),
    .B(_0924_),
    .X(_0925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3401_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .A2(net657),
    .Y(_0926_),
    .B1(net671));
 sg13g2_a22oi_1 _3402_ (.Y(_0927_),
    .B1(net667),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ),
    .A2(net678),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3403_ (.Y(_0928_),
    .B1(net675),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .A2(net680),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3404_ (.X(_0929_),
    .A(_0926_),
    .B(_0927_),
    .C(_0928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3405_ (.Y(_0930_),
    .B1(_0925_),
    .B2(_0929_),
    .A2(net671),
    .A1(_1446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3406_ (.Y(_0931_),
    .A(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3407_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net590),
    .A2(_0908_),
    .Y(_0932_),
    .B1(_0930_));
 sg13g2_nand3_1 _3408_ (.B(_0908_),
    .C(_0930_),
    .A(net590),
    .Y(_0933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3409_ (.Y(_0934_),
    .B(_0933_),
    .A_N(_0932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3410_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0935_),
    .B(_0934_),
    .A(net598));
 sg13g2_nand3_1 _3411_ (.B(_0907_),
    .C(_0931_),
    .A(_0885_),
    .Y(_0936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3412_ (.Y(_0937_),
    .A(_0913_),
    .B(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3413_ (.A(net606),
    .B(_0937_),
    .X(_0938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3414_ (.A(_0287_),
    .B(_0869_),
    .X(_0939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3415_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net572),
    .A2(net595),
    .Y(_0940_),
    .B1(_0939_));
 sg13g2_nor3_1 _3416_ (.A(net586),
    .B(_0938_),
    .C(_0940_),
    .Y(_0941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3417_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net591),
    .A2(_0800_),
    .Y(_0942_),
    .B1(_0766_));
 sg13g2_or2_1 _3418_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0943_),
    .B(_0942_),
    .A(_0802_));
 sg13g2_nor3_1 _3419_ (.A(_0766_),
    .B(net592),
    .C(_0835_),
    .Y(_0944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3420_ (.B1(_0766_),
    .VDD(VPWR),
    .Y(_0945_),
    .VSS(VGND),
    .A1(net592),
    .A2(_0835_));
 sg13g2_nand2b_1 _3421_ (.Y(_0946_),
    .B(_0945_),
    .A_N(_0944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3422_ (.Y(_0069_),
    .B1(_0935_),
    .B2(_0941_),
    .A2(net586),
    .A1(_1446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3423_ (.Y(_0947_),
    .B1(net675),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .A2(net678),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3424_ (.A2(net676),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .B1(net671),
    .X(_0948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3425_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ),
    .C1(_0948_),
    .B1(net657),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .Y(_0949_),
    .A2(net661));
 sg13g2_a22oi_1 _3426_ (.Y(_0950_),
    .B1(net667),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .A2(net681),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3427_ (.Y(_0951_),
    .A(_0947_),
    .B(_0950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3428_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .C1(_0951_),
    .B1(net663),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .Y(_0952_),
    .A2(net666));
 sg13g2_a22oi_1 _3429_ (.Y(_0953_),
    .B1(_0949_),
    .B2(_0952_),
    .A2(net671),
    .A1(_1474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3430_ (.VDD(VPWR),
    .Y(_0954_),
    .A(_0953_),
    .VSS(VGND));
 sg13g2_nand3_1 _3431_ (.B(_0930_),
    .C(_0953_),
    .A(_0908_),
    .Y(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3432_ (.B(_0908_),
    .C(_0930_),
    .A(net590),
    .Y(_0956_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0953_));
 sg13g2_xnor2_1 _3433_ (.Y(_0957_),
    .A(_0933_),
    .B(_0953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3434_ (.B1(_0844_),
    .VDD(VPWR),
    .Y(_0958_),
    .VSS(VGND),
    .A1(_0756_),
    .A2(_0944_));
 sg13g2_a21oi_1 _3435_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net622),
    .A2(_0958_),
    .Y(_0959_),
    .B1(net598));
 sg13g2_o21ai_1 _3436_ (.B1(_0959_),
    .VDD(VPWR),
    .Y(_0960_),
    .VSS(VGND),
    .A1(net622),
    .A2(_0957_));
 sg13g2_nand4_1 _3437_ (.B(_0907_),
    .C(_0931_),
    .A(_0885_),
    .Y(_0961_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0954_));
 sg13g2_xnor2_1 _3438_ (.Y(_0962_),
    .A(_0936_),
    .B(_0953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3439_ (.Y(_0963_),
    .A(_0755_),
    .B(_0802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3440_ (.B1(net607),
    .VDD(VPWR),
    .Y(_0964_),
    .VSS(VGND),
    .A1(net671),
    .A2(_0963_));
 sg13g2_inv_1 _3441_ (.VDD(VPWR),
    .Y(_0965_),
    .A(_0964_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3442_ (.B1(_0965_),
    .VDD(VPWR),
    .Y(_0966_),
    .VSS(VGND),
    .A1(net622),
    .A2(_0962_));
 sg13g2_nand2b_1 _3443_ (.Y(_0967_),
    .B(net596),
    .A_N(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3444_ (.B1(_0967_),
    .VDD(VPWR),
    .Y(_0968_),
    .VSS(VGND),
    .A1(net13),
    .A2(net596));
 sg13g2_nand3_1 _3445_ (.B(_0966_),
    .C(_0968_),
    .A(_0960_),
    .Y(_0969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3446_ (.A0(_0969_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[0][4] ),
    .S(net586),
    .X(_0070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3447_ (.Y(_0970_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][5] ),
    .B(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3448_ (.Y(_0971_),
    .B1(net674),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .A2(net680),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3449_ (.A2(net660),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .B1(net670),
    .X(_0972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3450_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .C1(_0972_),
    .B1(net664),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .Y(_0973_),
    .A2(net668));
 sg13g2_a22oi_1 _3451_ (.Y(_0974_),
    .B1(net665),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .A2(net677),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3452_ (.Y(_0975_),
    .A(_0971_),
    .B(_0974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3453_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .C1(_0975_),
    .B1(net656),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .Y(_0976_),
    .A2(net679));
 sg13g2_a22oi_1 _3454_ (.Y(_0977_),
    .B1(_0973_),
    .B2(_0976_),
    .A2(net670),
    .A1(_1480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3455_ (.B(_0930_),
    .C(_0953_),
    .A(_0908_),
    .Y(_0978_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0977_));
 sg13g2_nand2b_1 _3456_ (.Y(_0979_),
    .B(_0977_),
    .A_N(_0956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3457_ (.Y(_0980_),
    .A(_0956_),
    .B(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3458_ (.Y(_0981_),
    .A(_0741_),
    .B(_0844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3459_ (.B1(net602),
    .VDD(VPWR),
    .Y(_0982_),
    .VSS(VGND),
    .A1(net669),
    .A2(_0981_));
 sg13g2_a21oi_1 _3460_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net669),
    .A2(_0980_),
    .Y(_0983_),
    .B1(_0982_));
 sg13g2_nand2_1 _3461_ (.Y(_0984_),
    .A(_0288_),
    .B(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3462_ (.Y(_0985_),
    .B1(_0869_),
    .B2(_0984_),
    .A2(net595),
    .A1(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3463_ (.A(net587),
    .B(_0983_),
    .C(_0985_),
    .X(_0986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3464_ (.Y(_0987_),
    .A(_0741_),
    .B(_0803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3465_ (.Y(_0988_),
    .A(_0741_),
    .B(_0838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3466_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0742_),
    .A2(_0837_),
    .Y(_0989_),
    .B1(net653));
 sg13g2_a22oi_1 _3467_ (.Y(_0990_),
    .B1(_0988_),
    .B2(_0989_),
    .A2(_0987_),
    .A1(net653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3468_ (.A(_0953_),
    .B(_0977_),
    .Y(_0991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3469_ (.A(_0885_),
    .B(_0907_),
    .C(_0931_),
    .D(_0991_),
    .X(_0992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3470_ (.Y(_0993_),
    .A(_0961_),
    .B(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3471_ (.Y(_0994_),
    .A(_0955_),
    .B(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3472_ (.A0(_0993_),
    .A1(_0994_),
    .S(net651),
    .X(_0995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3473_ (.A(net712),
    .B(_0995_),
    .Y(_0996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3474_ (.B1(net711),
    .VDD(VPWR),
    .Y(_0997_),
    .VSS(VGND),
    .A1(net669),
    .A2(_0990_));
 sg13g2_a21oi_1 _3475_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net669),
    .A2(_0995_),
    .Y(_0998_),
    .B1(_0997_));
 sg13g2_o21ai_1 _3476_ (.B1(_0970_),
    .VDD(VPWR),
    .Y(_0071_),
    .VSS(VGND),
    .A1(_0986_),
    .A2(_0998_));
 sg13g2_nand2_1 _3477_ (.Y(_0999_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .B(net674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3478_ (.Y(_1000_),
    .B1(net664),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .A2(net677),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3479_ (.Y(_1001_),
    .A(net621),
    .B(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3480_ (.Y(_1002_),
    .B1(net665),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .A2(net668),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3481_ (.Y(_1003_),
    .B1(net660),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .A2(net679),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3482_ (.Y(_1004_),
    .B1(net656),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ),
    .A2(net681),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3483_ (.B(_1002_),
    .C(_1003_),
    .A(_0999_),
    .Y(_1005_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1004_));
 sg13g2_nand2_1 _3484_ (.Y(_1006_),
    .A(_1484_),
    .B(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3485_ (.B1(_1006_),
    .VDD(VPWR),
    .Y(_1007_),
    .VSS(VGND),
    .A1(_1001_),
    .A2(_1005_));
 sg13g2_xor2_1 _3486_ (.B(_1007_),
    .A(_0992_),
    .X(_1008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3487_ (.Y(_1009_),
    .A(_0733_),
    .B(_0804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3488_ (.B1(net606),
    .VDD(VPWR),
    .Y(_1010_),
    .VSS(VGND),
    .A1(net669),
    .A2(_1009_));
 sg13g2_a21oi_1 _3489_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net669),
    .A2(_1008_),
    .Y(_1011_),
    .B1(_1010_));
 sg13g2_nor2_1 _3490_ (.A(_0978_),
    .B(_1007_),
    .Y(_1012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3491_ (.A(net591),
    .B(_0978_),
    .C(_1007_),
    .Y(_1013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3492_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1013_),
    .Y(_1014_),
    .A2(_1007_),
    .A1(_0979_));
 sg13g2_xnor2_1 _3493_ (.Y(_1015_),
    .A(_0732_),
    .B(_0845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3494_ (.B1(net602),
    .VDD(VPWR),
    .Y(_1016_),
    .VSS(VGND),
    .A1(net669),
    .A2(_1015_));
 sg13g2_inv_1 _3495_ (.VDD(VPWR),
    .Y(_1017_),
    .A(_1016_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3496_ (.B1(_1017_),
    .VDD(VPWR),
    .Y(_1018_),
    .VSS(VGND),
    .A1(net621),
    .A2(_1014_));
 sg13g2_mux2_1 _3497_ (.A0(net15),
    .A1(net33),
    .S(net595),
    .X(_1019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3498_ (.A(net587),
    .B(_1011_),
    .C(_1019_),
    .Y(_1020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3499_ (.Y(_0072_),
    .B1(_1018_),
    .B2(_1020_),
    .A2(net587),
    .A1(_1484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3500_ (.Y(_1021_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .B(net664),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3501_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .C1(net672),
    .B1(net666),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .Y(_1022_),
    .A2(net677));
 sg13g2_a22oi_1 _3502_ (.Y(_1023_),
    .B1(net662),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .A2(_0695_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3503_ (.Y(_1024_),
    .B1(net678),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .A2(net681),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3504_ (.B(_1023_),
    .C(_1024_),
    .A(_1021_),
    .Y(_1025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3505_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ),
    .C1(_1025_),
    .B1(net658),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .Y(_1026_),
    .A2(net675));
 sg13g2_a22oi_1 _3506_ (.Y(_1027_),
    .B1(_1022_),
    .B2(_1026_),
    .A2(net672),
    .A1(_1494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3507_ (.X(_1028_),
    .A(_0992_),
    .B(_1007_),
    .C(_1027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3508_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0992_),
    .A2(_1007_),
    .Y(_1029_),
    .B1(_1027_));
 sg13g2_nor2_1 _3509_ (.A(_1028_),
    .B(_1029_),
    .Y(_1030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3510_ (.A(net621),
    .B(_1028_),
    .C(_1029_),
    .Y(_1031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3511_ (.Y(_1032_),
    .A(_0721_),
    .B(_0805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3512_ (.B1(net606),
    .VDD(VPWR),
    .Y(_1033_),
    .VSS(VGND),
    .A1(net669),
    .A2(_1032_));
 sg13g2_xnor2_1 _3513_ (.Y(_1034_),
    .A(_0722_),
    .B(_0840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3514_ (.B(_0827_),
    .C(_1034_),
    .A(net621),
    .Y(_1035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3515_ (.B1(net712),
    .VDD(VPWR),
    .Y(_1036_),
    .VSS(VGND),
    .A1(_0289_),
    .A2(net595));
 sg13g2_a21oi_1 _3516_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net34),
    .A2(net595),
    .Y(_1037_),
    .B1(_1036_));
 sg13g2_a21oi_1 _3517_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net652),
    .A2(_1035_),
    .Y(_1038_),
    .B1(_1037_));
 sg13g2_o21ai_1 _3518_ (.B1(_1038_),
    .VDD(VPWR),
    .Y(_1039_),
    .VSS(VGND),
    .A1(_1031_),
    .A2(_1033_));
 sg13g2_xor2_1 _3519_ (.B(_1027_),
    .A(_1013_),
    .X(_1040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3520_ (.B1(_0721_),
    .VDD(VPWR),
    .Y(_1041_),
    .VSS(VGND),
    .A1(net592),
    .A2(_0840_));
 sg13g2_nand2b_2 _3521_ (.Y(_1042_),
    .B(_1041_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0846_));
 sg13g2_a221oi_1 _3522_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net602),
    .C1(net621),
    .B1(_1040_),
    .A1(net597),
    .Y(_1043_),
    .A2(_0862_));
 sg13g2_a22oi_1 _3523_ (.Y(_0073_),
    .B1(_1039_),
    .B2(_1043_),
    .A2(net586),
    .A1(_1494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3524_ (.A(_0700_),
    .B(net596),
    .X(_1044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3525_ (.A(net590),
    .B(net605),
    .Y(_1045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3526_ (.A(net31),
    .B(_0874_),
    .C(_1045_),
    .Y(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3527_ (.A(net592),
    .B(net598),
    .Y(_1047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3528_ (.A(net585),
    .B(_1046_),
    .C(_1047_),
    .Y(_1048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3529_ (.A2(net585),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .B1(_1048_),
    .X(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3530_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net600),
    .A2(_0898_),
    .Y(_1049_),
    .B1(net584));
 sg13g2_nor2_1 _3531_ (.A(net605),
    .B(_0898_),
    .Y(_1050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3532_ (.A(net18),
    .B(_1050_),
    .Y(_1051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3533_ (.Y(_0075_),
    .B1(_1049_),
    .B2(_1051_),
    .A2(net584),
    .A1(_1467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3534_ (.A2(_0921_),
    .A1(net607),
    .B1(net19),
    .X(_1052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3535_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net601),
    .C1(_1052_),
    .B1(_0911_),
    .A1(_0700_),
    .Y(_1053_),
    .A2(net596));
 sg13g2_a21oi_1 _3536_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1457_),
    .A2(net585),
    .Y(_0076_),
    .B1(_1053_));
 sg13g2_a21o_1 _3537_ (.A2(_0943_),
    .A1(_0828_),
    .B1(net20),
    .X(_1054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3538_ (.A(net598),
    .B(_0946_),
    .Y(_1055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3539_ (.A(net584),
    .B(_1054_),
    .C(_1055_),
    .Y(_1056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3540_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1453_),
    .A2(net584),
    .Y(_0077_),
    .B1(_1056_));
 sg13g2_nor2_1 _3541_ (.A(net32),
    .B(_0850_),
    .Y(_1057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3542_ (.B1(net601),
    .VDD(VPWR),
    .Y(_1058_),
    .VSS(VGND),
    .A1(net663),
    .A2(_0958_));
 sg13g2_o21ai_1 _3543_ (.B1(_1058_),
    .VDD(VPWR),
    .Y(_1059_),
    .VSS(VGND),
    .A1(net605),
    .A2(_0963_));
 sg13g2_nor2_2 _3544_ (.A(_1057_),
    .B(_1059_),
    .Y(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3545_ (.A0(_1060_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .S(net585),
    .X(_0078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3546_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0828_),
    .A2(_0987_),
    .Y(_1061_),
    .B1(net22));
 sg13g2_nor2_1 _3547_ (.A(net599),
    .B(_0981_),
    .Y(_1062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3548_ (.A(net584),
    .B(_1062_),
    .Y(_1063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3549_ (.Y(_0079_),
    .B1(_1061_),
    .B2(_1063_),
    .A2(net584),
    .A1(_1483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3550_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net33),
    .Y(_1064_),
    .A2(_1009_),
    .A1(net606));
 sg13g2_nand2_2 _3551_ (.Y(_1065_),
    .A(net603),
    .B(_1015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3552_ (.VDD(VPWR),
    .Y(_1066_),
    .A(_1065_),
    .VSS(VGND));
 sg13g2_nor2_1 _3553_ (.A(net584),
    .B(_1066_),
    .Y(_1067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3554_ (.Y(_0080_),
    .B1(_1064_),
    .B2(_1067_),
    .A2(net584),
    .A1(_1493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3555_ (.A(_0829_),
    .B(_1032_),
    .Y(_1068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3556_ (.A(net34),
    .B(_1068_),
    .Y(_1069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3557_ (.A(_0872_),
    .B(_1034_),
    .X(_1070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3558_ (.Y(_1071_),
    .B(_1069_),
    .A_N(_1070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3559_ (.A(net598),
    .B(_1042_),
    .Y(_1072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3560_ (.A(net585),
    .B(_1071_),
    .C(_1072_),
    .Y(_1073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3561_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1501_),
    .A2(net585),
    .Y(_0081_),
    .B1(_1073_));
 sg13g2_nand2_1 _3562_ (.Y(_1074_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .B(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3563_ (.A(net618),
    .B(net684),
    .Y(_1075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3564_ (.Y(_1076_),
    .B(net667),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net685));
 sg13g2_nor2_1 _3565_ (.A(net9),
    .B(_0828_),
    .Y(_1077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3566_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0829_),
    .A2(_1076_),
    .Y(_1078_),
    .B1(_1077_));
 sg13g2_a21o_1 _3567_ (.A2(_1076_),
    .A1(net31),
    .B1(_1078_),
    .X(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3568_ (.A(_0808_),
    .B(net713),
    .Y(_1080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3569_ (.B1(_1080_),
    .VDD(VPWR),
    .Y(_1081_),
    .VSS(VGND),
    .A1(_0695_),
    .A2(net590));
 sg13g2_a21oi_1 _3570_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1079_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(_0874_));
 sg13g2_and2_1 _3571_ (.A(net603),
    .B(_0847_),
    .X(_1083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3572_ (.Y(_1084_),
    .B(_0695_),
    .A_N(_1083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3573_ (.B1(_1074_),
    .VDD(VPWR),
    .Y(_0082_),
    .VSS(VGND),
    .A1(_1082_),
    .A2(_1084_));
 sg13g2_nand2_1 _3574_ (.Y(_1085_),
    .A(net600),
    .B(_0891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3575_ (.A(net605),
    .B(_0886_),
    .Y(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3576_ (.A(net18),
    .B_N(net684),
    .Y(_1087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3577_ (.B1(net605),
    .VDD(VPWR),
    .Y(_1088_),
    .VSS(VGND),
    .A1(net10),
    .A2(_1076_));
 sg13g2_o21ai_1 _3578_ (.B1(net668),
    .VDD(VPWR),
    .Y(_1089_),
    .VSS(VGND),
    .A1(_1087_),
    .A2(_1088_));
 sg13g2_nor2_1 _3579_ (.A(_1086_),
    .B(_1089_),
    .Y(_1090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3580_ (.Y(_0083_),
    .B1(_1085_),
    .B2(_1090_),
    .A2(net618),
    .A1(_1466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3581_ (.A0(net19),
    .A1(net11),
    .S(_1075_),
    .X(_1091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3582_ (.A(net600),
    .B(_0922_),
    .C(_1091_),
    .Y(_1092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3583_ (.A(net605),
    .B(_0914_),
    .Y(_1093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3584_ (.B1(_1093_),
    .VDD(VPWR),
    .Y(_1094_),
    .VSS(VGND),
    .A1(net668),
    .A2(_0921_));
 sg13g2_a221oi_1 _3585_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1094_),
    .C1(net618),
    .B1(_1092_),
    .A1(net600),
    .Y(_1095_),
    .A2(_0909_));
 sg13g2_a21o_1 _3586_ (.A2(net618),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .B1(_1095_),
    .X(_0084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3587_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0287_),
    .C1(_0850_),
    .B1(_1075_),
    .A1(net572),
    .Y(_1096_),
    .A2(net684));
 sg13g2_nor3_1 _3588_ (.A(net618),
    .B(_0938_),
    .C(_1096_),
    .Y(_1097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3589_ (.Y(_0085_),
    .B1(_0935_),
    .B2(_1097_),
    .A2(net618),
    .A1(_1452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3590_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .B(net667),
    .Y(_1098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3591_ (.Y(_1099_),
    .A(net601),
    .B(_0957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3592_ (.Y(_1100_),
    .A(net607),
    .B(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3593_ (.B1(net713),
    .VDD(VPWR),
    .Y(_1101_),
    .VSS(VGND),
    .A1(net13),
    .A2(_1076_));
 sg13g2_nand2b_1 _3594_ (.Y(_1102_),
    .B(net685),
    .A_N(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3595_ (.Y(_1103_),
    .B(_1102_),
    .A_N(_1101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3596_ (.B(_1099_),
    .C(_1100_),
    .A(net667),
    .Y(_1104_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1103_));
 sg13g2_nor2b_1 _3597_ (.A(_1098_),
    .B_N(_1104_),
    .Y(_0086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3598_ (.Y(_1105_),
    .B(_1076_),
    .A_N(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3599_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1106_),
    .B(net685),
    .A(net14));
 sg13g2_a221oi_1 _3600_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1106_),
    .C1(net618),
    .B1(_1105_),
    .A1(net606),
    .Y(_1107_),
    .A2(_0993_));
 sg13g2_a21oi_1 _3601_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net619),
    .A2(_0981_),
    .Y(_1108_),
    .B1(net599));
 sg13g2_nand2_1 _3602_ (.Y(_1109_),
    .A(_0980_),
    .B(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3603_ (.Y(_0087_),
    .B1(_1107_),
    .B2(_1109_),
    .A2(net619),
    .A1(_1482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3604_ (.Y(_1110_),
    .A(net602),
    .B(_1014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3605_ (.A0(net33),
    .A1(net15),
    .S(_1075_),
    .X(_1111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3606_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0732_),
    .A2(_0839_),
    .Y(_1112_),
    .B1(_0873_));
 sg13g2_nand2_1 _3607_ (.Y(_1113_),
    .A(_0840_),
    .B(_1112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3608_ (.A(net605),
    .B(_1008_),
    .Y(_1114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3609_ (.A(net619),
    .B(_1111_),
    .C(_1114_),
    .Y(_1115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3610_ (.Y(_0088_),
    .B1(_1110_),
    .B2(_1115_),
    .A2(net619),
    .A1(_1492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3611_ (.Y(_1116_),
    .A(net619),
    .B(_1042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3612_ (.B(_1040_),
    .C(_1116_),
    .A(net602),
    .Y(_1117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3613_ (.Y(_1118_),
    .B(_1076_),
    .A_N(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3614_ (.Y(_1119_),
    .A(_0289_),
    .B(_1075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3615_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1119_),
    .C1(net618),
    .B1(_1118_),
    .A1(net607),
    .Y(_1120_),
    .A2(_1030_));
 sg13g2_a22oi_1 _3616_ (.Y(_0089_),
    .B1(_1117_),
    .B2(_1120_),
    .A2(net619),
    .A1(_1500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3617_ (.A(net674),
    .B(_1075_),
    .Y(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3618_ (.Y(_1122_),
    .A(_0690_),
    .B(_1076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3619_ (.A(_1046_),
    .B(_1047_),
    .C(_1121_),
    .Y(_1123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3620_ (.A2(_1121_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .B1(_1123_),
    .X(_0090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3621_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net588),
    .A2(net651),
    .Y(_1124_),
    .B1(net600));
 sg13g2_nand2_1 _3622_ (.Y(_1125_),
    .A(_1051_),
    .B(_1124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3623_ (.Y(_1126_),
    .B(net600),
    .A_N(_0898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3624_ (.B(_1125_),
    .C(_1126_),
    .A(_1122_),
    .Y(_1127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3625_ (.B1(_1127_),
    .VDD(VPWR),
    .Y(_0091_),
    .VSS(VGND),
    .A1(_1465_),
    .A2(_1122_));
 sg13g2_nor2_1 _3626_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ),
    .B(_1122_),
    .Y(_1128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3627_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0835_),
    .C1(_1052_),
    .B1(_0918_),
    .A1(net601),
    .Y(_1129_),
    .A2(_0911_));
 sg13g2_a21oi_1 _3628_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1122_),
    .A2(_1129_),
    .Y(_0092_),
    .B1(_1128_));
 sg13g2_nor3_1 _3629_ (.A(_1054_),
    .B(_1055_),
    .C(_1121_),
    .Y(_1130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1451_),
    .A2(_1121_),
    .Y(_0093_),
    .B1(_1130_));
 sg13g2_mux2_1 _3631_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .A1(_1060_),
    .S(_1122_),
    .X(_0094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3632_ (.Y(_1131_),
    .B(_1061_),
    .A_N(_1062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3633_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .A1(_1131_),
    .S(_1122_),
    .X(_0095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3634_ (.Y(_1132_),
    .A(_1064_),
    .B(_1113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3635_ (.A(_1121_),
    .B(_1132_),
    .Y(_1133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3636_ (.Y(_0096_),
    .B1(_1133_),
    .B2(_1065_),
    .A2(_1121_),
    .A1(_1491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3637_ (.A(_1072_),
    .B(_1121_),
    .Y(_1134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3638_ (.Y(_0097_),
    .B1(_1134_),
    .B2(_1069_),
    .A2(_1121_),
    .A1(_1499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3639_ (.Y(_1135_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .B(net624),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3640_ (.Y(_1136_),
    .B(net678),
    .A_N(_1083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3641_ (.A(net623),
    .B(net684),
    .Y(_1137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3642_ (.Y(_1138_),
    .B(net678),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net685));
 sg13g2_a21oi_1 _3643_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0829_),
    .A2(_1138_),
    .Y(_1139_),
    .B1(_1077_));
 sg13g2_a21o_1 _3644_ (.A2(_1138_),
    .A1(net17),
    .B1(_1139_),
    .X(_1140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3645_ (.B1(_1080_),
    .VDD(VPWR),
    .Y(_1141_),
    .VSS(VGND),
    .A1(_0663_),
    .A2(_0789_));
 sg13g2_a21oi_1 _3646_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1140_),
    .A2(_1141_),
    .Y(_1142_),
    .B1(_0874_));
 sg13g2_o21ai_1 _3647_ (.B1(_1135_),
    .VDD(VPWR),
    .Y(_0098_),
    .VSS(VGND),
    .A1(_1136_),
    .A2(_1142_));
 sg13g2_o21ai_1 _3648_ (.B1(net597),
    .VDD(VPWR),
    .Y(_1143_),
    .VSS(VGND),
    .A1(net10),
    .A2(_1138_));
 sg13g2_nor2_1 _3649_ (.A(_1087_),
    .B(_1143_),
    .Y(_1144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3650_ (.A(net623),
    .B(_1086_),
    .C(_1144_),
    .Y(_1145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3651_ (.Y(_0099_),
    .B1(_1085_),
    .B2(_1145_),
    .A2(net623),
    .A1(_1464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3652_ (.A(net599),
    .B(_0909_),
    .Y(_1146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3653_ (.A(_1093_),
    .B(_1146_),
    .Y(_1147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3654_ (.Y(_1148_),
    .A(_2008_),
    .B(net685),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3655_ (.Y(_1149_),
    .A(_0849_),
    .B(_1138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3656_ (.B1(_1149_),
    .VDD(VPWR),
    .Y(_1150_),
    .VSS(VGND),
    .A1(_1673_),
    .A2(_1994_));
 sg13g2_a21oi_1 _3657_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1148_),
    .A2(_1150_),
    .Y(_1151_),
    .B1(net624));
 sg13g2_a22oi_1 _3658_ (.Y(_0100_),
    .B1(_1147_),
    .B2(_1151_),
    .A2(_0664_),
    .A1(_1456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3659_ (.Y(_1152_),
    .B1(_1149_),
    .B2(_0287_),
    .A2(net684),
    .A1(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3660_ (.A(net623),
    .B(_0938_),
    .C(_1152_),
    .Y(_1153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3661_ (.Y(_0101_),
    .B1(_0935_),
    .B2(_1153_),
    .A2(net623),
    .A1(_1450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3662_ (.A(_1099_),
    .B(_1100_),
    .X(_1154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3663_ (.Y(_1155_),
    .B(_1149_),
    .A_N(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3664_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1102_),
    .A2(_1155_),
    .Y(_1156_),
    .B1(net624));
 sg13g2_a22oi_1 _3665_ (.Y(_0102_),
    .B1(_1154_),
    .B2(_1156_),
    .A2(net624),
    .A1(_1479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3666_ (.Y(_1157_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .B(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3667_ (.Y(_1158_),
    .B1(_0984_),
    .B2(_1149_),
    .A2(net684),
    .A1(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3668_ (.A(net599),
    .B(_0980_),
    .Y(_1159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3669_ (.A(net623),
    .B(_1158_),
    .C(_1159_),
    .X(_1160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3670_ (.B1(_1157_),
    .VDD(VPWR),
    .Y(_0103_),
    .VSS(VGND),
    .A1(_0996_),
    .A2(_1160_));
 sg13g2_nand2_1 _3671_ (.Y(_1161_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .B(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3672_ (.A(net679),
    .B(_1009_),
    .Y(_1162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3673_ (.B1(net607),
    .VDD(VPWR),
    .Y(_1163_),
    .VSS(VGND),
    .A1(_1008_),
    .A2(_1162_));
 sg13g2_inv_1 _3674_ (.VDD(VPWR),
    .Y(_1164_),
    .A(_1163_),
    .VSS(VGND));
 sg13g2_a221oi_1 _3675_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net15),
    .C1(_0850_),
    .B1(_1137_),
    .A1(net33),
    .Y(_1165_),
    .A2(net684));
 sg13g2_nor2_1 _3676_ (.A(net624),
    .B(_1165_),
    .Y(_1166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3677_ (.B1(_1166_),
    .VDD(VPWR),
    .Y(_1167_),
    .VSS(VGND),
    .A1(net599),
    .A2(_1014_));
 sg13g2_o21ai_1 _3678_ (.B1(_1161_),
    .VDD(VPWR),
    .Y(_0104_),
    .VSS(VGND),
    .A1(_1164_),
    .A2(_1167_));
 sg13g2_o21ai_1 _3679_ (.B1(net712),
    .VDD(VPWR),
    .Y(_1168_),
    .VSS(VGND),
    .A1(_0289_),
    .A2(_1138_));
 sg13g2_a21oi_1 _3680_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net34),
    .A2(_1138_),
    .Y(_1169_),
    .B1(_1168_));
 sg13g2_nor2_1 _3681_ (.A(net652),
    .B(_1169_),
    .Y(_1170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3682_ (.B1(net607),
    .VDD(VPWR),
    .Y(_1171_),
    .VSS(VGND),
    .A1(net679),
    .A2(_1032_));
 sg13g2_o21ai_1 _3683_ (.B1(_1170_),
    .VDD(VPWR),
    .Y(_1172_),
    .VSS(VGND),
    .A1(_1030_),
    .A2(_1171_));
 sg13g2_a21oi_1 _3684_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net602),
    .A2(_1040_),
    .Y(_1173_),
    .B1(net624));
 sg13g2_a22oi_1 _3685_ (.Y(_0105_),
    .B1(_1172_),
    .B2(_1173_),
    .A2(net624),
    .A1(_1498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3686_ (.A(net677),
    .B(_1137_),
    .Y(_1174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3687_ (.A(_1046_),
    .B(_1047_),
    .C(net579),
    .Y(_1175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3688_ (.A2(net579),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .B1(_1175_),
    .X(_0106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3689_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net601),
    .C1(net18),
    .B1(_0898_),
    .A1(net588),
    .Y(_1176_),
    .A2(_0872_));
 sg13g2_nand2b_1 _3690_ (.Y(_1177_),
    .B(_1176_),
    .A_N(_1050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3691_ (.A0(_1177_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .S(net578),
    .X(_0107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3692_ (.A(net604),
    .B(_0922_),
    .C(_1052_),
    .Y(_1178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3693_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0666_),
    .A2(_0911_),
    .Y(_1179_),
    .B1(net598));
 sg13g2_nor3_1 _3694_ (.A(net578),
    .B(_1178_),
    .C(_1179_),
    .Y(_1180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3695_ (.A2(net578),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .B1(_1180_),
    .X(_0108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3696_ (.Y(_1181_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .B(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3697_ (.Y(_1182_),
    .A(_0766_),
    .B(_0835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3698_ (.Y(_1183_),
    .A(net654),
    .B(_0943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3699_ (.B1(_1183_),
    .VDD(VPWR),
    .Y(_1184_),
    .VSS(VGND),
    .A1(net654),
    .A2(_1182_));
 sg13g2_a22oi_1 _3700_ (.Y(_1185_),
    .B1(_0946_),
    .B2(net604),
    .A2(net597),
    .A1(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3701_ (.B1(_1185_),
    .VDD(VPWR),
    .Y(_1186_),
    .VSS(VGND),
    .A1(net713),
    .A2(_1184_));
 sg13g2_o21ai_1 _3702_ (.B1(_1181_),
    .VDD(VPWR),
    .Y(_0109_),
    .VSS(VGND),
    .A1(net579),
    .A2(_1186_));
 sg13g2_a21o_1 _3703_ (.A2(_0963_),
    .A1(net607),
    .B1(net32),
    .X(_1187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3704_ (.A(net598),
    .B(_0958_),
    .Y(_1188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3705_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1189_),
    .B(_1188_),
    .A(_1187_));
 sg13g2_mux2_1 _3706_ (.A0(_1189_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .S(net579),
    .X(_0110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3707_ (.Y(_1190_),
    .A(net602),
    .B(_0981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3708_ (.Y(_1191_),
    .B(net597),
    .A_N(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3709_ (.Y(_1192_),
    .A(_1190_),
    .B(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3710_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net711),
    .A2(_0990_),
    .Y(_1193_),
    .B1(_1192_));
 sg13g2_mux2_1 _3711_ (.A0(_1193_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .S(net578),
    .X(_0111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3712_ (.A(_1132_),
    .B(net578),
    .Y(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3713_ (.Y(_0112_),
    .B1(_1194_),
    .B2(_1065_),
    .A2(net578),
    .A1(_1490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3714_ (.Y(_1195_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .B(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3715_ (.A(net603),
    .B(_1071_),
    .Y(_1196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3716_ (.Y(_1197_),
    .A(net603),
    .B(_1042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3717_ (.Y(_1198_),
    .B(_1197_),
    .A_N(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3718_ (.B1(_1195_),
    .VDD(VPWR),
    .Y(_0113_),
    .VSS(VGND),
    .A1(_1196_),
    .A2(_1198_));
 sg13g2_nor3_1 _3719_ (.A(net616),
    .B(_1046_),
    .C(_1083_),
    .Y(_1199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3720_ (.A2(net616),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .B1(_1199_),
    .X(_0114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3721_ (.A(net18),
    .B(net617),
    .Y(_1200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3722_ (.Y(_0115_),
    .B1(_1085_),
    .B2(_1200_),
    .A2(net617),
    .A1(_1463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3723_ (.A(net617),
    .B(_1052_),
    .C(_1146_),
    .Y(_1201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3724_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1455_),
    .A2(net616),
    .Y(_0116_),
    .B1(_1201_));
 sg13g2_nor2_1 _3725_ (.A(net616),
    .B(_1054_),
    .Y(_1202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3726_ (.Y(_0117_),
    .B1(_0935_),
    .B2(_1202_),
    .A2(net616),
    .A1(_1449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3727_ (.A(net616),
    .B(_1187_),
    .Y(_1203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3728_ (.Y(_0118_),
    .B1(_1099_),
    .B2(_1203_),
    .A2(net616),
    .A1(_1478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3729_ (.Y(_1204_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .B(net617),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3730_ (.Y(_1205_),
    .A(net665),
    .B(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3731_ (.B1(_1204_),
    .VDD(VPWR),
    .Y(_0119_),
    .VSS(VGND),
    .A1(_1159_),
    .A2(_1205_));
 sg13g2_and2_1 _3732_ (.A(net665),
    .B(_1064_),
    .X(_1206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3733_ (.Y(_0120_),
    .B1(_1110_),
    .B2(_1206_),
    .A2(net617),
    .A1(_1489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3734_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net603),
    .A2(_1040_),
    .Y(_1207_),
    .B1(net616));
 sg13g2_a22oi_1 _3735_ (.Y(_0121_),
    .B1(_1069_),
    .B2(_1207_),
    .A2(net617),
    .A1(_1497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3736_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net680),
    .Y(_1208_),
    .A2(_1656_),
    .A1(_1595_));
 sg13g2_nor3_1 _3737_ (.A(_1046_),
    .B(_1047_),
    .C(net594),
    .Y(_1209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3738_ (.A2(net593),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .B1(_1209_),
    .X(_0122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3739_ (.A0(_1177_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .S(net593),
    .X(_0123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3740_ (.Y(_1210_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ),
    .B(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3741_ (.B1(_1210_),
    .VDD(VPWR),
    .Y(_0124_),
    .VSS(VGND),
    .A1(_1129_),
    .A2(net594));
 sg13g2_mux2_1 _3742_ (.A0(_1185_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ),
    .S(net593),
    .X(_0125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3743_ (.A0(_1189_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .S(net594),
    .X(_0126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3744_ (.Y(_1211_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ),
    .B(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3745_ (.B1(_1211_),
    .VDD(VPWR),
    .Y(_0127_),
    .VSS(VGND),
    .A1(_1192_),
    .A2(net593));
 sg13g2_nand2_1 _3746_ (.Y(_1212_),
    .A(_1064_),
    .B(_1065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3747_ (.A(net593),
    .B(_1212_),
    .Y(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3748_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1488_),
    .A2(net593),
    .Y(_0128_),
    .B1(_1213_));
 sg13g2_nor2_1 _3749_ (.A(_1072_),
    .B(net594),
    .Y(_1214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3750_ (.Y(_0129_),
    .B1(_1214_),
    .B2(_1069_),
    .A2(net594),
    .A1(_1496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3751_ (.B1(net713),
    .VDD(VPWR),
    .Y(_1215_),
    .VSS(VGND),
    .A1(net9),
    .A2(net652));
 sg13g2_a21oi_1 _3752_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0711_),
    .A2(_0842_),
    .Y(_1216_),
    .B1(_0873_));
 sg13g2_a21oi_1 _3753_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0843_),
    .A2(_1216_),
    .Y(_1217_),
    .B1(_1045_));
 sg13g2_a221oi_1 _3754_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1217_),
    .C1(net612),
    .B1(_1215_),
    .A1(net603),
    .Y(_1218_),
    .A2(_0847_));
 sg13g2_a21o_1 _3755_ (.A2(net614),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .B1(_1218_),
    .X(_0130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3756_ (.B1(net711),
    .VDD(VPWR),
    .Y(_1219_),
    .VSS(VGND),
    .A1(net651),
    .A2(_0898_));
 sg13g2_nor2_1 _3757_ (.A(net660),
    .B(net588),
    .Y(_1220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3758_ (.A(net653),
    .B(_1220_),
    .Y(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3759_ (.Y(_1222_),
    .B1(_1221_),
    .B2(_0896_),
    .A2(_1219_),
    .A1(_0893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3760_ (.A(net611),
    .B(_0892_),
    .C(_1222_),
    .Y(_1223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3761_ (.A2(net611),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .B1(_1223_),
    .X(_0131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3762_ (.Y(_1224_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .B(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3763_ (.Y(_1225_),
    .A(net660),
    .B(_0910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3764_ (.Y(_1226_),
    .A(_0888_),
    .B(_0907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3765_ (.Y(_1227_),
    .A(_0872_),
    .B(_1226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3766_ (.A(net11),
    .B(net600),
    .Y(_1228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3767_ (.B1(_1228_),
    .VDD(VPWR),
    .Y(_1229_),
    .VSS(VGND),
    .A1(_0908_),
    .A2(_1227_));
 sg13g2_a21oi_1 _3768_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net606),
    .A2(_0921_),
    .Y(_1230_),
    .B1(_1229_));
 sg13g2_o21ai_1 _3769_ (.B1(_1224_),
    .VDD(VPWR),
    .Y(_0132_),
    .VSS(VGND),
    .A1(_1225_),
    .A2(_1230_));
 sg13g2_a221oi_1 _3770_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net601),
    .C1(net611),
    .B1(_0934_),
    .A1(_0287_),
    .Y(_1231_),
    .A2(_0849_));
 sg13g2_xnor2_1 _3771_ (.Y(_1232_),
    .A(_0908_),
    .B(_0931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3772_ (.A0(_0937_),
    .A1(_1232_),
    .S(net651),
    .X(_1233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3773_ (.A2(_1184_),
    .A1(net613),
    .B1(net713),
    .X(_1234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3774_ (.B1(_1231_),
    .VDD(VPWR),
    .Y(_1235_),
    .VSS(VGND),
    .A1(_1233_),
    .A2(_1234_));
 sg13g2_o21ai_1 _3775_ (.B1(_1235_),
    .VDD(VPWR),
    .Y(_0133_),
    .VSS(VGND),
    .A1(_1448_),
    .A2(net661));
 sg13g2_a21oi_1 _3776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0908_),
    .A2(_0930_),
    .Y(_1236_),
    .B1(_0953_));
 sg13g2_nand2_1 _3777_ (.Y(_1237_),
    .A(_0872_),
    .B(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3778_ (.A(_1236_),
    .B(_1237_),
    .Y(_1238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3779_ (.A(net13),
    .B(net613),
    .C(_1238_),
    .Y(_1239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3780_ (.Y(_0134_),
    .B1(_1099_),
    .B2(_1239_),
    .A2(net613),
    .A1(_1477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3781_ (.Y(_1240_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .B(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3782_ (.B(net660),
    .C(_0984_),
    .Y(_1241_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1159_));
 sg13g2_o21ai_1 _3783_ (.B1(_1240_),
    .VDD(VPWR),
    .Y(_0135_),
    .VSS(VGND),
    .A1(_0996_),
    .A2(_1241_));
 sg13g2_o21ai_1 _3784_ (.B1(_0872_),
    .VDD(VPWR),
    .Y(_1242_),
    .VSS(VGND),
    .A1(_0978_),
    .A2(_1007_));
 sg13g2_a21oi_1 _3785_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0978_),
    .A2(_1007_),
    .Y(_1243_),
    .B1(_1242_));
 sg13g2_nor3_1 _3786_ (.A(net15),
    .B(net611),
    .C(_1243_),
    .Y(_1244_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3787_ (.Y(_0136_),
    .B1(_1110_),
    .B2(_1244_),
    .A2(net612),
    .A1(_1487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3788_ (.Y(_1245_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .B(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3789_ (.B(_1027_),
    .A(_1012_),
    .X(_1246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3790_ (.B(_0702_),
    .C(net654),
    .A(_0289_),
    .Y(_1247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3791_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net713),
    .C1(_1068_),
    .B1(_1247_),
    .A1(_0872_),
    .Y(_1248_),
    .A2(_1246_));
 sg13g2_o21ai_1 _3792_ (.B1(net662),
    .VDD(VPWR),
    .Y(_1249_),
    .VSS(VGND),
    .A1(_0834_),
    .A2(_1040_));
 sg13g2_o21ai_1 _3793_ (.B1(_1245_),
    .VDD(VPWR),
    .Y(_0137_),
    .VSS(VGND),
    .A1(_1248_),
    .A2(_1249_));
 sg13g2_nor3_1 _3794_ (.A(net613),
    .B(_1046_),
    .C(_1047_),
    .Y(_1250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3795_ (.A2(net614),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .B1(_1250_),
    .X(_0138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3796_ (.Y(_1251_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .B(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3797_ (.B1(_1251_),
    .VDD(VPWR),
    .Y(_0139_),
    .VSS(VGND),
    .A1(net611),
    .A2(_1176_));
 sg13g2_nor2_1 _3798_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ),
    .B(net661),
    .Y(_1252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3799_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net661),
    .A2(_1129_),
    .Y(_0140_),
    .B1(_1252_));
 sg13g2_nor2_1 _3800_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .B(net661),
    .Y(_1253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3801_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net662),
    .A2(_1186_),
    .Y(_0141_),
    .B1(_1253_));
 sg13g2_nor2_1 _3802_ (.A(_0756_),
    .B(_0836_),
    .Y(_1254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3803_ (.A(net654),
    .B(net713),
    .C(_0837_),
    .D(_1254_),
    .Y(_1255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3804_ (.A(net613),
    .B(_1189_),
    .C(_1255_),
    .Y(_1256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3805_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1476_),
    .A2(net613),
    .Y(_0142_),
    .B1(_1256_));
 sg13g2_mux2_1 _3806_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .A1(_1193_),
    .S(net660),
    .X(_0143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3807_ (.A(net612),
    .B(_1066_),
    .C(_1132_),
    .Y(_1257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3808_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1486_),
    .A2(net612),
    .Y(_0144_),
    .B1(_1257_));
 sg13g2_nor3_1 _3809_ (.A(net613),
    .B(_1071_),
    .C(_1072_),
    .Y(_1258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3810_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1495_),
    .A2(net614),
    .Y(_0145_),
    .B1(_1258_));
 sg13g2_nand2_1 _3811_ (.Y(_1259_),
    .A(net609),
    .B(net592),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3812_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1080_),
    .A2(_1259_),
    .Y(_1260_),
    .B1(_1077_));
 sg13g2_nor2_1 _3813_ (.A(net609),
    .B(_1083_),
    .Y(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3814_ (.B1(_1261_),
    .VDD(VPWR),
    .Y(_1262_),
    .VSS(VGND),
    .A1(_0874_),
    .A2(_1260_));
 sg13g2_o21ai_1 _3815_ (.B1(_1262_),
    .VDD(VPWR),
    .Y(_0146_),
    .VSS(VGND),
    .A1(_1469_),
    .A2(net658));
 sg13g2_nand2_1 _3816_ (.Y(_1263_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ),
    .B(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3817_ (.B(_0893_),
    .C(net655),
    .Y(_1264_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0887_));
 sg13g2_o21ai_1 _3818_ (.B1(_1263_),
    .VDD(VPWR),
    .Y(_0147_),
    .VSS(VGND),
    .A1(_0892_),
    .A2(_1264_));
 sg13g2_nor2_1 _3819_ (.A(net11),
    .B(net608),
    .Y(_1265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3820_ (.Y(_0148_),
    .B1(_1147_),
    .B2(_1265_),
    .A2(net608),
    .A1(_1454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3821_ (.A2(_1184_),
    .A1(net608),
    .B1(net713),
    .X(_1266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3822_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net601),
    .C1(net610),
    .B1(_0934_),
    .A1(_0287_),
    .Y(_1267_),
    .A2(_0849_));
 sg13g2_o21ai_1 _3823_ (.B1(_1267_),
    .VDD(VPWR),
    .Y(_1268_),
    .VSS(VGND),
    .A1(_1233_),
    .A2(_1266_));
 sg13g2_o21ai_1 _3824_ (.B1(_1268_),
    .VDD(VPWR),
    .Y(_0149_),
    .VSS(VGND),
    .A1(_1447_),
    .A2(net655));
 sg13g2_nor2_1 _3825_ (.A(net13),
    .B(net608),
    .Y(_1269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3826_ (.Y(_0150_),
    .B1(_1154_),
    .B2(_1269_),
    .A2(net608),
    .A1(_1475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3827_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net711),
    .C1(net610),
    .B1(_0995_),
    .A1(net602),
    .Y(_1270_),
    .A2(_0980_));
 sg13g2_a22oi_1 _3828_ (.Y(_0151_),
    .B1(_1270_),
    .B2(_0288_),
    .A2(net610),
    .A1(_1481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3829_ (.A(net15),
    .B(net610),
    .C(_1114_),
    .Y(_1271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3830_ (.Y(_0152_),
    .B1(_1110_),
    .B2(_1271_),
    .A2(net610),
    .A1(_1485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3831_ (.Y(_1272_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ),
    .B(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3832_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net610),
    .A2(_1032_),
    .Y(_1273_),
    .B1(net605));
 sg13g2_nand3_1 _3833_ (.B(net656),
    .C(net653),
    .A(_0289_),
    .Y(_1274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3834_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net712),
    .C1(_1070_),
    .B1(_1274_),
    .A1(_1030_),
    .Y(_1275_),
    .A2(_1273_));
 sg13g2_o21ai_1 _3835_ (.B1(net656),
    .VDD(VPWR),
    .Y(_1276_),
    .VSS(VGND),
    .A1(net599),
    .A2(_1040_));
 sg13g2_o21ai_1 _3836_ (.B1(_1272_),
    .VDD(VPWR),
    .Y(_0153_),
    .VSS(VGND),
    .A1(_1275_),
    .A2(_1276_));
 sg13g2_or2_1 _3837_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1277_),
    .B(\sap_3_inst.reg_file.array_serializer_inst.state[0] ),
    .A(\sap_3_inst.reg_file.array_serializer_inst.state[1] ));
 sg13g2_inv_2 _3838_ (.Y(_0154_),
    .A(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3839_ (.A(\sap_3_inst.reg_file.array_serializer_inst.state[0] ),
    .B_N(\sap_3_inst.reg_file.array_serializer_inst.state[1] ),
    .Y(_1278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3840_ (.A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .B(net817),
    .X(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3841_ (.Y(_1280_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .B(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3842_ (.Y(_1281_),
    .A(_1278_),
    .B(_1280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3843_ (.A(net75),
    .B_N(\sap_3_inst.reg_file.array_serializer_inst.state[0] ),
    .Y(_1282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3844_ (.A2(_1280_),
    .A1(_1278_),
    .B1(_1282_),
    .X(_0155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3845_ (.A(net817),
    .B(_1278_),
    .Y(_1283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3846_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net817),
    .A2(_0155_),
    .Y(_0156_),
    .B1(_1283_));
 sg13g2_a21oi_1 _3847_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net817),
    .A2(_0155_),
    .Y(_1284_),
    .B1(net56));
 sg13g2_nand2_1 _3848_ (.Y(_1285_),
    .A(_1278_),
    .B(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3849_ (.A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .B(_1285_),
    .Y(_1286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3850_ (.A(_1282_),
    .B(_1284_),
    .C(_1286_),
    .Y(_0157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3851_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1440_),
    .A2(_1285_),
    .Y(_0158_),
    .B1(_1282_));
 sg13g2_a21o_1 _3852_ (.A2(regFile_serial_start),
    .A1(net75),
    .B1(_0154_),
    .X(_0159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3853_ (.A(net71),
    .B(_0155_),
    .Y(_1287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3854_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net817),
    .A2(_1502_),
    .Y(_1288_),
    .B1(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ));
 sg13g2_o21ai_1 _3855_ (.B1(_1288_),
    .VDD(VPWR),
    .Y(_1289_),
    .VSS(VGND),
    .A1(net817),
    .A2(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[1] ));
 sg13g2_nor2b_1 _3856_ (.A(net817),
    .B_N(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .Y(_1290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3857_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[3] ),
    .C1(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .B1(_1290_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[4] ),
    .Y(_1291_),
    .A2(_1279_));
 sg13g2_nand2b_1 _3858_ (.Y(_1292_),
    .B(net817),
    .A_N(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3859_ (.B1(_1292_),
    .VDD(VPWR),
    .Y(_1293_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[0] ),
    .A2(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[5] ));
 sg13g2_o21ai_1 _3860_ (.B1(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .VDD(VPWR),
    .Y(_1294_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .A2(_1293_));
 sg13g2_a21oi_1 _3861_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[7] ),
    .A2(_1290_),
    .Y(_1295_),
    .B1(_1294_));
 sg13g2_a21oi_1 _3862_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1289_),
    .A2(_1291_),
    .Y(_1296_),
    .B1(_1295_));
 sg13g2_a22oi_1 _3863_ (.Y(_1297_),
    .B1(_1296_),
    .B2(_1278_),
    .A2(_1281_),
    .A1(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3864_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0155_),
    .A2(_1297_),
    .Y(_0160_),
    .B1(_1287_));
 sg13g2_nand2b_2 _3865_ (.Y(_1298_),
    .B(net815),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net816));
 sg13g2_nand2b_2 _3866_ (.Y(_1299_),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ));
 sg13g2_nor2_2 _3867_ (.A(_1298_),
    .B(_1299_),
    .Y(_1300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3868_ (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .C(_1298_),
    .Y(_1301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3869_ (.Y(_1302_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3870_ (.Y(_1303_),
    .B(net816),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net815));
 sg13g2_nor2_1 _3871_ (.A(_1302_),
    .B(_1303_),
    .Y(_1304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3872_ (.Y(_1305_),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ));
 sg13g2_nor2_2 _3873_ (.A(_1298_),
    .B(_1305_),
    .Y(_1306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3874_ (.A(net815),
    .B(net816),
    .C(_1305_),
    .Y(_1307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3875_ (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .C(_1303_),
    .Y(_1308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3876_ (.A(_1299_),
    .B(_1303_),
    .Y(_1309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3877_ (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .C(_1302_),
    .Y(_1310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3878_ (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .C(net815),
    .D(net816),
    .Y(_1311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3879_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net815),
    .A2(net816),
    .Y(_1312_),
    .B1(_1311_));
 sg13g2_a21o_1 _3880_ (.A2(net816),
    .A1(net815),
    .B1(_1311_),
    .X(_1313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3881_ (.A(_1303_),
    .B(_1305_),
    .Y(_1314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3882_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .A2(_1314_),
    .Y(_1315_),
    .B1(net808));
 sg13g2_nor2_2 _3883_ (.A(_1298_),
    .B(_1302_),
    .Y(_1316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3884_ (.A(net815),
    .B(net816),
    .C(_1299_),
    .Y(_1317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3885_ (.Y(_1318_),
    .B1(net809),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .A2(_1300_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3886_ (.Y(_1319_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .A2(_1307_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3887_ (.Y(_1320_),
    .B1(_1309_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .A2(net810),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3888_ (.Y(_1321_),
    .B1(_1306_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ),
    .A2(_1301_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3889_ (.B(_1318_),
    .C(_1320_),
    .A(_1315_),
    .Y(_1322_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1321_));
 sg13g2_a221oi_1 _3890_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .C1(_1322_),
    .B1(_1317_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .Y(_1323_),
    .A2(_1308_));
 sg13g2_a221oi_1 _3891_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1323_),
    .C1(net812),
    .B1(_1319_),
    .A1(_1468_),
    .Y(_1324_),
    .A2(net808));
 sg13g2_a21o_1 _3892_ (.A2(net811),
    .A1(net54),
    .B1(_1324_),
    .X(_0161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3893_ (.Y(_1325_),
    .B1(_1301_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .A2(_1300_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3894_ (.Y(_1326_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .A2(net810),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3895_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .A2(_1308_),
    .Y(_1327_),
    .B1(net807));
 sg13g2_a22oi_1 _3896_ (.Y(_1328_),
    .B1(_1317_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .A2(_1306_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3897_ (.Y(_1329_),
    .B1(net809),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .A2(_1309_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3898_ (.B(_1327_),
    .C(_1328_),
    .A(_1325_),
    .Y(_1330_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1329_));
 sg13g2_a221oi_1 _3899_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .C1(_1330_),
    .B1(_1314_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .Y(_1331_),
    .A2(_1307_));
 sg13g2_a221oi_1 _3900_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1331_),
    .C1(net812),
    .B1(_1326_),
    .A1(_1461_),
    .Y(_1332_),
    .A2(net807));
 sg13g2_a21o_1 _3901_ (.A2(net811),
    .A1(net55),
    .B1(_1332_),
    .X(_0162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3902_ (.Y(_1333_),
    .B1(_1317_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .A2(_1314_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3903_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .A2(_1306_),
    .Y(_1334_),
    .B1(net808));
 sg13g2_a22oi_1 _3904_ (.Y(_1335_),
    .B1(_1307_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .A2(net810),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3905_ (.Y(_1336_),
    .B1(_1309_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .A2(_1301_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3906_ (.Y(_1337_),
    .B1(net809),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ),
    .A2(_1300_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3907_ (.B(_1335_),
    .C(_1336_),
    .A(_1334_),
    .Y(_1338_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1337_));
 sg13g2_a221oi_1 _3908_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .C1(_1338_),
    .B1(_1316_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .Y(_1339_),
    .A2(_1308_));
 sg13g2_o21ai_1 _3909_ (.B1(_0154_),
    .VDD(VPWR),
    .Y(_1340_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[0][2] ),
    .A2(_1312_));
 sg13g2_a21o_1 _3910_ (.A2(_1339_),
    .A1(_1333_),
    .B1(_1340_),
    .X(_1341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3911_ (.B1(_1341_),
    .VDD(VPWR),
    .Y(_0163_),
    .VSS(VGND),
    .A1(_1502_),
    .A2(_0154_));
 sg13g2_a22oi_1 _3912_ (.Y(_1342_),
    .B1(net810),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ),
    .A2(_1300_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3913_ (.Y(_1343_),
    .B1(_1314_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .A2(_1301_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3914_ (.Y(_1344_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .A2(_1309_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3915_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .A2(_1306_),
    .Y(_1345_),
    .B1(net807));
 sg13g2_a22oi_1 _3916_ (.Y(_1346_),
    .B1(net809),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .A2(_1307_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3917_ (.B(_1343_),
    .C(_1345_),
    .A(_1342_),
    .Y(_1347_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1346_));
 sg13g2_a221oi_1 _3918_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .C1(_1347_),
    .B1(_1317_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .Y(_1348_),
    .A2(_1308_));
 sg13g2_a221oi_1 _3919_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1348_),
    .C1(net812),
    .B1(_1344_),
    .A1(_1446_),
    .Y(_1349_),
    .A2(net807));
 sg13g2_a21o_1 _3920_ (.A2(net811),
    .A1(net63),
    .B1(_1349_),
    .X(_0164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3921_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .A2(_1309_),
    .Y(_1350_),
    .B1(net808));
 sg13g2_a22oi_1 _3922_ (.Y(_1351_),
    .B1(_1317_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .A2(_1304_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3923_ (.Y(_1352_),
    .B1(_1307_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .A2(_1306_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3924_ (.Y(_1353_),
    .B1(_1314_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .A2(_1300_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3925_ (.Y(_1354_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .A2(_1310_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3926_ (.B(_1351_),
    .C(_1353_),
    .A(_1350_),
    .Y(_1355_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1354_));
 sg13g2_a221oi_1 _3927_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ),
    .C1(_1355_),
    .B1(_1308_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .Y(_1356_),
    .A2(_1301_));
 sg13g2_a221oi_1 _3928_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1356_),
    .C1(net811),
    .B1(_1352_),
    .A1(_1474_),
    .Y(_1357_),
    .A2(net808));
 sg13g2_a21o_1 _3929_ (.A2(net811),
    .A1(net50),
    .B1(_1357_),
    .X(_0165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3930_ (.Y(_1358_),
    .B1(_1317_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .A2(_1316_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3931_ (.Y(_1359_),
    .B1(net809),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .A2(_1307_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3932_ (.Y(_1360_),
    .B1(_1308_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .A2(net810),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3933_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .A2(_1314_),
    .Y(_1361_),
    .B1(net807));
 sg13g2_a22oi_1 _3934_ (.Y(_1362_),
    .B1(_1309_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .A2(_1300_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3935_ (.B(_1360_),
    .C(_1361_),
    .A(_1358_),
    .Y(_1363_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1362_));
 sg13g2_a221oi_1 _3936_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .C1(_1363_),
    .B1(_1306_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .Y(_1364_),
    .A2(_1301_));
 sg13g2_a221oi_1 _3937_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1364_),
    .C1(net812),
    .B1(_1359_),
    .A1(_1480_),
    .Y(_1365_),
    .A2(net807));
 sg13g2_a21o_1 _3938_ (.A2(net811),
    .A1(net51),
    .B1(_1365_),
    .X(_0166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3939_ (.Y(_1366_),
    .B1(_1317_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .A2(_1306_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3940_ (.Y(_1367_),
    .B1(_1309_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .A2(_1301_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3941_ (.Y(_1368_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .A2(_1307_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3942_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .A2(net810),
    .Y(_1369_),
    .B1(net807));
 sg13g2_a22oi_1 _3943_ (.Y(_1370_),
    .B1(_1314_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .A2(_1300_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3944_ (.B(_1367_),
    .C(_1369_),
    .A(_1366_),
    .Y(_1371_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1370_));
 sg13g2_a221oi_1 _3945_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .C1(_1371_),
    .B1(net809),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .Y(_1372_),
    .A2(_1308_));
 sg13g2_a221oi_1 _3946_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1372_),
    .C1(net812),
    .B1(_1368_),
    .A1(_1484_),
    .Y(_1373_),
    .A2(net807));
 sg13g2_a21o_1 _3947_ (.A2(net811),
    .A1(net53),
    .B1(_1373_),
    .X(_0167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3948_ (.Y(_1374_),
    .B1(_1314_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .A2(net809),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3949_ (.Y(_1375_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .A2(_1300_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3950_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .A2(_1309_),
    .Y(_1376_),
    .B1(net808));
 sg13g2_a22oi_1 _3951_ (.Y(_1377_),
    .B1(_1308_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .A2(_1306_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3952_ (.Y(_1378_),
    .B1(_1307_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .A2(_1301_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3953_ (.B(_1376_),
    .C(_1377_),
    .A(_1374_),
    .Y(_1379_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1378_));
 sg13g2_a221oi_1 _3954_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .C1(_1379_),
    .B1(_1317_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .Y(_1380_),
    .A2(net810));
 sg13g2_a221oi_1 _3955_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1380_),
    .C1(net812),
    .B1(_1375_),
    .A1(_1494_),
    .Y(_1381_),
    .A2(net808));
 sg13g2_a21o_1 _3956_ (.A2(net812),
    .A1(net52),
    .B1(_1381_),
    .X(_0168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3957_ (.A(net608),
    .B(_1046_),
    .C(_1047_),
    .Y(_1382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3958_ (.A2(net609),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .B1(_1382_),
    .X(_0169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3959_ (.B(_1125_),
    .C(_1126_),
    .A(net655),
    .Y(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3960_ (.B1(_1383_),
    .VDD(VPWR),
    .Y(_0170_),
    .VSS(VGND),
    .A1(_1462_),
    .A2(net655));
 sg13g2_nor2_1 _3961_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .B(net657),
    .Y(_1384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3962_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net657),
    .A2(_1129_),
    .Y(_0171_),
    .B1(_1384_));
 sg13g2_nand2_1 _3963_ (.Y(_1385_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .B(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3964_ (.B1(_1385_),
    .VDD(VPWR),
    .Y(_0172_),
    .VSS(VGND),
    .A1(net608),
    .A2(_1186_));
 sg13g2_mux2_1 _3965_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .A1(_1189_),
    .S(net657),
    .X(_0173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3966_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .A1(_1131_),
    .S(net655),
    .X(_0174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3967_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .A1(_1212_),
    .S(net656),
    .X(_0175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3968_ (.Y(_1386_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .B(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3969_ (.Y(_1387_),
    .A(net658),
    .B(_1197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3970_ (.B1(_1386_),
    .VDD(VPWR),
    .Y(_0176_),
    .VSS(VGND),
    .A1(_1196_),
    .A2(_1387_));
 sg13g2_nor3_1 _3971_ (.A(net724),
    .B(_0301_),
    .C(_0303_),
    .Y(_1388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3972_ (.A(_1856_),
    .B(_1388_),
    .Y(_1389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3973_ (.A(_0316_),
    .B_N(net709),
    .Y(_1390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3974_ (.A(_1459_),
    .B(net709),
    .Y(_1391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3975_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0323_),
    .A2(net709),
    .Y(_1392_),
    .B1(_1391_));
 sg13g2_nand2_1 _3976_ (.Y(_1393_),
    .A(\sap_3_inst.alu.act[0] ),
    .B(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3977_ (.B1(_1393_),
    .VDD(VPWR),
    .Y(_0177_),
    .VSS(VGND),
    .A1(net582),
    .A2(_1392_));
 sg13g2_nor2_1 _3978_ (.A(_1458_),
    .B(net709),
    .Y(_1394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3979_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0359_),
    .A2(net709),
    .Y(_1395_),
    .B1(_1394_));
 sg13g2_nand2_1 _3980_ (.Y(_1396_),
    .A(\sap_3_inst.alu.act[1] ),
    .B(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3981_ (.B1(_1396_),
    .VDD(VPWR),
    .Y(_0178_),
    .VSS(VGND),
    .A1(net582),
    .A2(_1395_));
 sg13g2_nor2b_1 _3982_ (.A(net709),
    .B_N(net801),
    .Y(_1397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3983_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0388_),
    .A2(net710),
    .Y(_1398_),
    .B1(_1397_));
 sg13g2_nand2_1 _3984_ (.Y(_1399_),
    .A(\sap_3_inst.alu.act[2] ),
    .B(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3985_ (.B1(_1399_),
    .VDD(VPWR),
    .Y(_0179_),
    .VSS(VGND),
    .A1(net582),
    .A2(_1398_));
 sg13g2_nor2_1 _3986_ (.A(_1445_),
    .B(net709),
    .Y(_1400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3987_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0434_),
    .A2(net709),
    .Y(_1401_),
    .B1(_1400_));
 sg13g2_nand2_1 _3988_ (.Y(_1402_),
    .A(\sap_3_inst.alu.act[3] ),
    .B(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3989_ (.B1(_1402_),
    .VDD(VPWR),
    .Y(_0180_),
    .VSS(VGND),
    .A1(net582),
    .A2(_1401_));
 sg13g2_nor2_1 _3990_ (.A(_1460_),
    .B(_1389_),
    .Y(_1403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3991_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0463_),
    .A2(net710),
    .Y(_1404_),
    .B1(_1403_));
 sg13g2_nand2_1 _3992_ (.Y(_1405_),
    .A(\sap_3_inst.alu.act[4] ),
    .B(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3993_ (.B1(_1405_),
    .VDD(VPWR),
    .Y(_0181_),
    .VSS(VGND),
    .A1(net583),
    .A2(_1404_));
 sg13g2_nand2_1 _3994_ (.Y(_1406_),
    .A(\sap_3_inst.alu.act[5] ),
    .B(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3995_ (.A(net710),
    .B_N(net793),
    .Y(_1407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3996_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0496_),
    .A2(net710),
    .Y(_1408_),
    .B1(_1407_));
 sg13g2_o21ai_1 _3997_ (.B1(_1406_),
    .VDD(VPWR),
    .Y(_0182_),
    .VSS(VGND),
    .A1(net583),
    .A2(_1408_));
 sg13g2_nand2b_1 _3998_ (.Y(_1409_),
    .B(net710),
    .A_N(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3999_ (.B1(_1409_),
    .VDD(VPWR),
    .Y(_1410_),
    .VSS(VGND),
    .A1(net790),
    .A2(net710));
 sg13g2_nand2_1 _4000_ (.Y(_1411_),
    .A(\sap_3_inst.alu.act[6] ),
    .B(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4001_ (.B1(_1411_),
    .VDD(VPWR),
    .Y(_0183_),
    .VSS(VGND),
    .A1(net583),
    .A2(_1410_));
 sg13g2_nor2b_1 _4002_ (.A(net710),
    .B_N(net788),
    .Y(_1412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4003_ (.Y(_1413_),
    .A(\sap_3_inst.alu.act[7] ),
    .B(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4004_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0552_),
    .A2(_1389_),
    .Y(_1414_),
    .B1(_1412_));
 sg13g2_o21ai_1 _4005_ (.B1(_1413_),
    .VDD(VPWR),
    .Y(_0184_),
    .VSS(VGND),
    .A1(net583),
    .A2(_1414_));
 sg13g2_nor2_2 _4006_ (.A(_1437_),
    .B(\u_ser.state[0] ),
    .Y(_1415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4007_ (.Y(_1416_),
    .A(\u_ser.bit_pos[1] ),
    .B(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4008_ (.Y(_1417_),
    .A(_1415_),
    .B(_1416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4009_ (.B1(_1415_),
    .VDD(VPWR),
    .Y(_1418_),
    .VSS(VGND),
    .A1(_1439_),
    .A2(_1416_));
 sg13g2_o21ai_1 _4010_ (.B1(_1418_),
    .VDD(VPWR),
    .Y(_0186_),
    .VSS(VGND),
    .A1(\u_ser.state[1] ),
    .A2(_1438_));
 sg13g2_nand3b_1 _4011_ (.B(\u_ser.shadow_reg[7] ),
    .C(\u_ser.bit_pos[1] ),
    .Y(_1419_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net814));
 sg13g2_nand2b_1 _4012_ (.Y(_1420_),
    .B(net814),
    .A_N(\u_ser.shadow_reg[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4013_ (.B1(_1420_),
    .VDD(VPWR),
    .Y(_1421_),
    .VSS(VGND),
    .A1(\u_ser.bit_pos[0] ),
    .A2(\u_ser.shadow_reg[5] ));
 sg13g2_o21ai_1 _4014_ (.B1(_1419_),
    .VDD(VPWR),
    .Y(_1422_),
    .VSS(VGND),
    .A1(\u_ser.bit_pos[1] ),
    .A2(_1421_));
 sg13g2_nand3_1 _4015_ (.B(_1415_),
    .C(_1422_),
    .A(\u_ser.bit_pos[2] ),
    .Y(_1423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _4016_ (.S0(net814),
    .A0(\u_ser.shadow_reg[1] ),
    .A1(\u_ser.shadow_reg[2] ),
    .A2(\u_ser.shadow_reg[3] ),
    .A3(\u_ser.shadow_reg[4] ),
    .S1(\u_ser.bit_pos[1] ),
    .X(_1424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4017_ (.B(_1415_),
    .C(_1424_),
    .A(_1439_),
    .Y(_1425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4018_ (.B1(\u_ser.shadow_reg[0] ),
    .VDD(VPWR),
    .Y(_1426_),
    .VSS(VGND),
    .A1(_1437_),
    .A2(\u_ser.state[0] ));
 sg13g2_nand4_1 _4019_ (.B(_1423_),
    .C(_1425_),
    .A(_0186_),
    .Y(_1427_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1426_));
 sg13g2_o21ai_1 _4020_ (.B1(_1427_),
    .VDD(VPWR),
    .Y(_1428_),
    .VSS(VGND),
    .A1(net78),
    .A2(_0186_));
 sg13g2_inv_1 _4021_ (.VDD(VPWR),
    .Y(_0187_),
    .A(_1428_),
    .VSS(VGND));
 sg13g2_a21o_1 _4022_ (.A2(net72),
    .A1(\u_ser.state[1] ),
    .B1(net813),
    .X(_0188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4023_ (.A(_1440_),
    .B(_1285_),
    .Y(_1429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4024_ (.B(_1429_),
    .A(net74),
    .X(_0189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4025_ (.Y(_1430_),
    .B(_1429_),
    .A_N(_1302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4026_ (.A2(_1429_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .B1(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .X(_1431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4027_ (.A(_1430_),
    .B(_1431_),
    .X(_0190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4028_ (.Y(_1432_),
    .B1(_1430_),
    .B2(net816),
    .A2(_1429_),
    .A1(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4029_ (.VDD(VPWR),
    .Y(_0191_),
    .A(_1432_),
    .VSS(VGND));
 sg13g2_a22oi_1 _4030_ (.Y(_1433_),
    .B1(_1430_),
    .B2(net815),
    .A2(_1429_),
    .A1(net810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4031_ (.VDD(VPWR),
    .Y(_0192_),
    .A(_1433_),
    .VSS(VGND));
 sg13g2_nor2_1 _4032_ (.A(net814),
    .B(_1415_),
    .Y(_1434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4033_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net814),
    .A2(_0186_),
    .Y(_0193_),
    .B1(_1434_));
 sg13g2_a21oi_1 _4034_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net814),
    .A2(_0186_),
    .Y(_1435_),
    .B1(net70));
 sg13g2_a21oi_1 _4035_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1417_),
    .A2(_0186_),
    .Y(_0194_),
    .B1(_1435_));
 sg13g2_nand3_1 _4036_ (.B(net814),
    .C(_1415_),
    .A(\u_ser.bit_pos[1] ),
    .Y(_1436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4037_ (.Y(_0195_),
    .B1(_1439_),
    .B2(_1436_),
    .A2(net61),
    .A1(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4039__4 (.VDD(VPWR),
    .Y(net40),
    .A(\clknet_leaf_0_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4040__5 (.VDD(VPWR),
    .Y(net41),
    .A(\clknet_leaf_0_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4041__6 (.VDD(VPWR),
    .Y(net42),
    .A(\clknet_leaf_2_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4042__7 (.VDD(VPWR),
    .Y(net43),
    .A(\clknet_leaf_2_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4043__8 (.VDD(VPWR),
    .Y(net44),
    .A(\clknet_leaf_2_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4044__9 (.VDD(VPWR),
    .Y(net45),
    .A(\clknet_leaf_2_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4045__10 (.VDD(VPWR),
    .Y(net46),
    .A(\clknet_leaf_1_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4046__11 (.VDD(VPWR),
    .Y(net47),
    .A(\clknet_leaf_1_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4047__12 (.VDD(VPWR),
    .Y(net48),
    .A(\clknet_leaf_0_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4048__13 (.VDD(VPWR),
    .Y(net49),
    .A(\clknet_leaf_1_sap_3_inst.alu.clk ),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_regs_0_clk_div_two (.A(\sap_3_inst.alu.clk ),
    .X(\sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _4049_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0017_),
    .Q(\u_ser.shadow_reg[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _4050_ (.RESET_B(net832),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0018_),
    .Q(\u_ser.shadow_reg[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _4051_ (.RESET_B(net836),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0019_),
    .Q(\u_ser.shadow_reg[2] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4052_ (.RESET_B(net832),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0020_),
    .Q(\u_ser.shadow_reg[3] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _4053_ (.RESET_B(net836),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0021_),
    .Q(\u_ser.shadow_reg[4] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4054_ (.RESET_B(net836),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0022_),
    .Q(\u_ser.shadow_reg[5] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4055_ (.RESET_B(net836),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0023_),
    .Q(\u_ser.shadow_reg[6] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4056_ (.RESET_B(net836),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0024_),
    .Q(\u_ser.shadow_reg[7] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4057_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0025_),
    .Q(\sap_3_inst.alu.flags[0] ),
    .CLK(net38));
 sg13g2_dfrbpq_2 _4058_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0026_),
    .Q(\sap_3_inst.alu.flags[1] ),
    .CLK(net39));
 sg13g2_dfrbpq_1 _4059_ (.RESET_B(net822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0027_),
    .Q(\sap_3_inst.alu.flags[2] ),
    .CLK(net40));
 sg13g2_dfrbpq_1 _4060_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0028_),
    .Q(\sap_3_inst.alu.flags[3] ),
    .CLK(net41));
 sg13g2_dfrbpq_1 _4061_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0001_),
    .Q(\sap_3_inst.controller.stage[0] ),
    .CLK(net42));
 sg13g2_dfrbpq_2 _4062_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0002_),
    .Q(\sap_3_inst.controller.stage[1] ),
    .CLK(net43));
 sg13g2_dfrbpq_1 _4063_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0003_),
    .Q(\sap_3_inst.controller.stage[2] ),
    .CLK(net44));
 sg13g2_dfrbpq_2 _4064_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0004_),
    .Q(\sap_3_inst.controller.stage[3] ),
    .CLK(net45));
 sg13g2_dfrbpq_1 _4065_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0029_),
    .Q(\sap_3_inst.alu.flags[4] ),
    .CLK(net46));
 sg13g2_dfrbpq_1 _4066_ (.RESET_B(net838),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0030_),
    .Q(\sap_3_inst.alu.flags[5] ),
    .CLK(net47));
 sg13g2_dfrbpq_1 _4067_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0031_),
    .Q(\sap_3_inst.alu.flags[6] ),
    .CLK(net48));
 sg13g2_dfrbpq_1 _4068_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0032_),
    .Q(\sap_3_inst.alu.flags[7] ),
    .CLK(net49));
 sg13g2_dfrbpq_1 _4069_ (.RESET_B(net832),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0033_),
    .Q(\sap_3_inst.alu.acc[0] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4070_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0034_),
    .Q(\sap_3_inst.alu.acc[1] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4071_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0035_),
    .Q(\sap_3_inst.alu.acc[2] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4072_ (.RESET_B(net838),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0036_),
    .Q(\sap_3_inst.alu.acc[3] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4073_ (.RESET_B(net838),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0037_),
    .Q(\sap_3_inst.alu.acc[4] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4074_ (.RESET_B(net838),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0038_),
    .Q(\sap_3_inst.alu.acc[5] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4075_ (.RESET_B(net839),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0039_),
    .Q(\sap_3_inst.alu.acc[6] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4076_ (.RESET_B(net839),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0040_),
    .Q(\sap_3_inst.alu.acc[7] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4077_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0041_),
    .Q(\sap_3_inst.out[0] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4078_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0042_),
    .Q(\sap_3_inst.out[1] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4079_ (.RESET_B(net836),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0043_),
    .Q(\sap_3_inst.out[2] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4080_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0044_),
    .Q(\sap_3_inst.out[3] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4081_ (.RESET_B(net837),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0045_),
    .Q(\sap_3_inst.out[4] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4082_ (.RESET_B(net837),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0046_),
    .Q(\sap_3_inst.out[5] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4083_ (.RESET_B(net837),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0047_),
    .Q(\sap_3_inst.out[6] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4084_ (.RESET_B(net840),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0048_),
    .Q(\sap_3_inst.out[7] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4085_ (.RESET_B(net838),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0049_),
    .Q(\sap_3_inst.alu.carry ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4086_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0050_),
    .Q(\sap_3_inst.alu.tmp[0] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4087_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0051_),
    .Q(\sap_3_inst.alu.tmp[1] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4088_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0052_),
    .Q(\sap_3_inst.alu.tmp[2] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4089_ (.RESET_B(net838),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0053_),
    .Q(\sap_3_inst.alu.tmp[3] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4090_ (.RESET_B(net838),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0054_),
    .Q(\sap_3_inst.alu.tmp[4] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4091_ (.RESET_B(net838),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0055_),
    .Q(\sap_3_inst.alu.tmp[5] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4092_ (.RESET_B(net839),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0056_),
    .Q(\sap_3_inst.alu.tmp[6] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4093_ (.RESET_B(net839),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0057_),
    .Q(\sap_3_inst.alu.tmp[7] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4094_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0058_),
    .Q(\sap_3_inst.controller.opcode[0] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4095_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0059_),
    .Q(\sap_3_inst.controller.opcode[1] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4096_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0060_),
    .Q(\sap_3_inst.controller.opcode[2] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4097_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0061_),
    .Q(\sap_3_inst.controller.opcode[3] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4098_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0062_),
    .Q(\sap_3_inst.controller.opcode[4] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4099_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0063_),
    .Q(\sap_3_inst.controller.opcode[5] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4100_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0064_),
    .Q(\sap_3_inst.controller.opcode[6] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4101_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0065_),
    .Q(\sap_3_inst.controller.opcode[7] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4102_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0066_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][0] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4103_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0067_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][1] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4104_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0068_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][2] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4105_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0069_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][3] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4106_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0070_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][4] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4107_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0071_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][5] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4108_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0072_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][6] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4109_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0073_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][7] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4110_ (.RESET_B(net843),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0074_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4111_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0075_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4112_ (.RESET_B(net842),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0076_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4113_ (.RESET_B(net822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0077_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4114_ (.RESET_B(net841),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0078_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4115_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0079_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4116_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0080_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4117_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0081_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4118_ (.RESET_B(net843),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4119_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0083_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4120_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0084_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4121_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0085_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4122_ (.RESET_B(net842),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0086_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4123_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0087_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4124_ (.RESET_B(net825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0088_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4125_ (.RESET_B(net826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0089_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4126_ (.RESET_B(net843),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0090_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4127_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0091_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4128_ (.RESET_B(net841),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0092_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4129_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0093_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4130_ (.RESET_B(net841),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0094_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4131_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0095_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4132_ (.RESET_B(net826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0096_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4133_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0097_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4134_ (.RESET_B(net843),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0098_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4135_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0099_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4136_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0100_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4137_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0101_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4138_ (.RESET_B(net842),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0102_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4139_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0103_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4140_ (.RESET_B(net825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0104_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4141_ (.RESET_B(net826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0105_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4142_ (.RESET_B(net844),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0106_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4143_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0107_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4144_ (.RESET_B(net842),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0108_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4145_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0109_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4146_ (.RESET_B(net841),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0110_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4147_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0111_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4148_ (.RESET_B(net826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0112_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4149_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0113_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4150_ (.RESET_B(net843),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0114_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4151_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0115_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4152_ (.RESET_B(net842),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0116_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4153_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0117_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4154_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0118_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4155_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0119_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4156_ (.RESET_B(net825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0120_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4157_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0121_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4158_ (.RESET_B(net843),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0122_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4159_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0123_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4160_ (.RESET_B(net841),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0124_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4161_ (.RESET_B(net822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0125_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4162_ (.RESET_B(net845),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0126_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4163_ (.RESET_B(net826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0127_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4164_ (.RESET_B(net826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0128_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4165_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0129_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4166_ (.RESET_B(net843),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0130_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4167_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4168_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0132_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4169_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0133_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4170_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0134_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4171_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0135_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4172_ (.RESET_B(net825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0136_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4173_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0137_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4174_ (.RESET_B(net844),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0138_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4175_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0139_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4176_ (.RESET_B(net841),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0140_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4177_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0141_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4178_ (.RESET_B(net842),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0142_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4179_ (.RESET_B(net825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0143_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4180_ (.RESET_B(net826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0144_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4181_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0145_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4182_ (.RESET_B(net843),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0146_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4183_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0147_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4184_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0148_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4185_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0149_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4186_ (.RESET_B(net842),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0150_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4187_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0151_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4188_ (.RESET_B(net825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0152_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4189_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0153_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4190_ (.RESET_B(net846),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0154_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.state[0] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _4191_ (.RESET_B(net846),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0155_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.state[1] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _4192_ (.RESET_B(net847),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0156_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[0] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _4193_ (.RESET_B(net847),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net57),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _4194_ (.RESET_B(net847),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0158_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _4195_ (.RESET_B(net846),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net76),
    .Q(regFile_serial_start),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _4196_ (.RESET_B(net846),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0160_),
    .Q(regFile_serial),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _4197_ (.RESET_B(net846),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0161_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[0] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4198_ (.RESET_B(net846),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0162_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[1] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4199_ (.RESET_B(net846),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0163_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[2] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _4200_ (.RESET_B(net841),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0164_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[3] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4201_ (.RESET_B(net846),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0165_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[4] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _4202_ (.RESET_B(net848),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0166_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[5] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _4203_ (.RESET_B(net848),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0167_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[6] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _4204_ (.RESET_B(net848),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0168_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[7] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _4205_ (.RESET_B(net844),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0169_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4206_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0170_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4207_ (.RESET_B(net841),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0171_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4208_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0172_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4209_ (.RESET_B(net845),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0173_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4210_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0174_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4211_ (.RESET_B(net826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0175_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4212_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0176_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4213_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net37),
    .Q(clk_div_out),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _4214_ (.RESET_B(net832),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0177_),
    .Q(\sap_3_inst.alu.act[0] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4215_ (.RESET_B(net832),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0178_),
    .Q(\sap_3_inst.alu.act[1] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4216_ (.RESET_B(net832),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0179_),
    .Q(\sap_3_inst.alu.act[2] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4217_ (.RESET_B(net832),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0180_),
    .Q(\sap_3_inst.alu.act[3] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4218_ (.RESET_B(net837),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0181_),
    .Q(\sap_3_inst.alu.act[4] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4219_ (.RESET_B(net837),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0182_),
    .Q(\sap_3_inst.alu.act[5] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4220_ (.RESET_B(net837),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0183_),
    .Q(\sap_3_inst.alu.act[6] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4221_ (.RESET_B(net837),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0184_),
    .Q(\sap_3_inst.alu.act[7] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4222_ (.RESET_B(net835),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net813),
    .Q(\u_ser.state[0] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _4223_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0186_),
    .Q(\u_ser.state[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _4224_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0187_),
    .Q(sap_3_outputReg_serial),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _4225_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net73),
    .Q(sap_3_outputReg_start_sync),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _4226_ (.RESET_B(net844),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0189_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _4227_ (.RESET_B(net844),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0190_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4228_ (.RESET_B(net844),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0191_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4229_ (.RESET_B(net844),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4230_ (.RESET_B(net836),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0193_),
    .Q(\u_ser.bit_pos[0] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _4231_ (.RESET_B(net836),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0194_),
    .Q(\u_ser.bit_pos[1] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4232_ (.RESET_B(net835),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net62),
    .Q(\u_ser.bit_pos[2] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_tielo heichips25_template_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net36));
 sg13g2_inv_1 _2081__1 (.VDD(VPWR),
    .Y(net37),
    .A(clknet_1_1__leaf_clk_div_out),
    .VSS(VGND));
 sg13g2_buf_1 _4235_ (.A(mem_ram_we),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _4236_ (.A(mem_mar_we),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _4237_ (.A(sap_3_outputReg_serial),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _4238_ (.A(sap_3_outputReg_start_sync),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 _4239_ (.A(regFile_serial),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 _4240_ (.A(regFile_serial_start),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_lgcp_1 \sap_3_inst.clock.clock_gate_inst  (.GATE(\sap_3_inst.clock.hlt ),
    .CLK(clknet_1_0__leaf_clk_div_out),
    .GCLK(\sap_3_inst.alu.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout572 (.A(_1982_),
    .X(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout573 (.A(net573),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout574 (.A(_0334_),
    .X(net574),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout575 (.A(_0334_),
    .X(net575),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout576 (.A(_1674_),
    .X(net576),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout577 (.A(_1674_),
    .X(net577),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout578 (.A(_1174_),
    .X(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout579 (.A(_1174_),
    .X(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout580 (.A(_0321_),
    .X(net580),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout581 (.A(_0321_),
    .X(net581),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout582 (.A(_1390_),
    .X(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout583 (.A(_1390_),
    .X(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout584 (.A(net585),
    .X(net584),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout585 (.A(_1044_),
    .X(net585),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout586 (.A(_0863_),
    .X(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout587 (.A(_0863_),
    .X(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout588 (.A(_0799_),
    .X(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout589 (.A(_0799_),
    .X(net589),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout590 (.A(_0789_),
    .X(net590),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout591 (.A(net592),
    .X(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout592 (.A(_0788_),
    .X(net592),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout593 (.A(_1208_),
    .X(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout594 (.A(_1208_),
    .X(net594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout595 (.A(net596),
    .X(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout596 (.A(_0868_),
    .X(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout597 (.A(_0849_),
    .X(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout598 (.A(_0834_),
    .X(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout599 (.A(_0834_),
    .X(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout600 (.A(net601),
    .X(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout601 (.A(net604),
    .X(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout602 (.A(net603),
    .X(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout603 (.A(net604),
    .X(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout604 (.A(_0833_),
    .X(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout605 (.A(_0829_),
    .X(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout606 (.A(net607),
    .X(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout607 (.A(_0828_),
    .X(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout608 (.A(_0705_),
    .X(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout609 (.A(_0705_),
    .X(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout610 (.A(_0705_),
    .X(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout611 (.A(net615),
    .X(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout612 (.A(net615),
    .X(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout613 (.A(net615),
    .X(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout614 (.A(net615),
    .X(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout615 (.A(_0703_),
    .X(net615),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout616 (.A(net617),
    .X(net616),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout617 (.A(_0698_),
    .X(net617),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout618 (.A(net620),
    .X(net618),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout619 (.A(net620),
    .X(net619),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout620 (.A(_0696_),
    .X(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout621 (.A(_0693_),
    .X(net621),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout622 (.A(_0693_),
    .X(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout623 (.A(net624),
    .X(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout624 (.A(_0664_),
    .X(net624),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout625 (.A(_0332_),
    .X(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout626 (.A(net627),
    .X(net626),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout627 (.A(_0311_),
    .X(net627),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout628 (.A(net629),
    .X(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout629 (.A(_1837_),
    .X(net629),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout630 (.A(_1812_),
    .X(net630),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout631 (.A(_1812_),
    .X(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout632 (.A(net633),
    .X(net632),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout633 (.A(_1811_),
    .X(net633),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout634 (.A(net635),
    .X(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout635 (.A(_1809_),
    .X(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout636 (.A(_1808_),
    .X(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout637 (.A(_1808_),
    .X(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout638 (.A(net639),
    .X(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout639 (.A(_1807_),
    .X(net639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout640 (.A(net641),
    .X(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout641 (.A(_1806_),
    .X(net641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout642 (.A(_1804_),
    .X(net642),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout643 (.A(_1804_),
    .X(net643),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout644 (.A(_1803_),
    .X(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout645 (.A(_1803_),
    .X(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout646 (.A(_1802_),
    .X(net646),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout647 (.A(_1802_),
    .X(net647),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout648 (.A(_1801_),
    .X(net648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout649 (.A(_1800_),
    .X(net649),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout650 (.A(_1800_),
    .X(net650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout651 (.A(_0821_),
    .X(net651),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout652 (.A(_0821_),
    .X(net652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout653 (.A(_0820_),
    .X(net653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout654 (.A(_0820_),
    .X(net654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout655 (.A(net659),
    .X(net655),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout656 (.A(net659),
    .X(net656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout657 (.A(net659),
    .X(net657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout658 (.A(net659),
    .X(net658),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout659 (.A(_0704_),
    .X(net659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout660 (.A(_0702_),
    .X(net660),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout661 (.A(net662),
    .X(net661),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout662 (.A(_0702_),
    .X(net662),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout663 (.A(_0699_),
    .X(net663),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout664 (.A(_0699_),
    .X(net664),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout665 (.A(_0697_),
    .X(net665),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout666 (.A(_0697_),
    .X(net666),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout667 (.A(net668),
    .X(net667),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout668 (.A(_0695_),
    .X(net668),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout669 (.A(net670),
    .X(net669),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout670 (.A(net673),
    .X(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout671 (.A(net673),
    .X(net671),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout672 (.A(net673),
    .X(net672),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout673 (.A(_0692_),
    .X(net673),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout674 (.A(_0689_),
    .X(net674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout675 (.A(_0689_),
    .X(net675),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout676 (.A(net677),
    .X(net676),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout677 (.A(_0665_),
    .X(net677),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout678 (.A(_0663_),
    .X(net678),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout679 (.A(_0663_),
    .X(net679),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout680 (.A(_0660_),
    .X(net680),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout681 (.A(_0660_),
    .X(net681),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout682 (.A(_0340_),
    .X(net682),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout683 (.A(_0338_),
    .X(net683),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout684 (.A(net685),
    .X(net684),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout685 (.A(_0867_),
    .X(net685),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout686 (.A(net687),
    .X(net686),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout687 (.A(_0688_),
    .X(net687),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout688 (.A(_0687_),
    .X(net688),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout689 (.A(_0687_),
    .X(net689),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout690 (.A(_0659_),
    .X(net690),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout691 (.A(_0658_),
    .X(net691),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout692 (.A(net696),
    .X(net692),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout693 (.A(net696),
    .X(net693),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout694 (.A(net695),
    .X(net694),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout695 (.A(net696),
    .X(net695),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout696 (.A(_0657_),
    .X(net696),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout697 (.A(net700),
    .X(net697),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout698 (.A(net699),
    .X(net698),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout699 (.A(net700),
    .X(net699),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout700 (.A(_0645_),
    .X(net700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout701 (.A(_0644_),
    .X(net701),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout702 (.A(_0644_),
    .X(net702),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout703 (.A(net706),
    .X(net703),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout704 (.A(net705),
    .X(net704),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout705 (.A(net706),
    .X(net705),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout706 (.A(_0619_),
    .X(net706),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout707 (.A(_0314_),
    .X(net707),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout708 (.A(_0314_),
    .X(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout709 (.A(net710),
    .X(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout710 (.A(_1389_),
    .X(net710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout711 (.A(_0827_),
    .X(net711),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout712 (.A(_0826_),
    .X(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout713 (.A(_0826_),
    .X(net713),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout714 (.A(_1944_),
    .X(net714),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout715 (.A(_0593_),
    .X(net715),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout716 (.A(_0593_),
    .X(net716),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout717 (.A(net719),
    .X(net717),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout718 (.A(net719),
    .X(net718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout719 (.A(_0267_),
    .X(net719),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout720 (.A(net721),
    .X(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout721 (.A(_1953_),
    .X(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout722 (.A(net723),
    .X(net722),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout723 (.A(_1730_),
    .X(net723),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout724 (.A(net725),
    .X(net724),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout725 (.A(_1714_),
    .X(net725),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout726 (.A(_1702_),
    .X(net726),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout727 (.A(_1678_),
    .X(net727),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout728 (.A(_1677_),
    .X(net728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout729 (.A(_1677_),
    .X(net729),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout730 (.A(_1633_),
    .X(net730),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout731 (.A(_1577_),
    .X(net731),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout732 (.A(_1572_),
    .X(net732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout733 (.A(_1572_),
    .X(net733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout734 (.A(_1560_),
    .X(net734),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout735 (.A(_1559_),
    .X(net735),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout736 (.A(_1552_),
    .X(net736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout737 (.A(_1552_),
    .X(net737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout738 (.A(net739),
    .X(net738),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout739 (.A(_1533_),
    .X(net739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout740 (.A(net741),
    .X(net740),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout741 (.A(net742),
    .X(net741),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout742 (.A(_1510_),
    .X(net742),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout743 (.A(net744),
    .X(net743),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout744 (.A(net745),
    .X(net744),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout745 (.A(_1509_),
    .X(net745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout746 (.A(_1631_),
    .X(net746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout747 (.A(_1631_),
    .X(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout748 (.A(_1605_),
    .X(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout749 (.A(_1600_),
    .X(net749),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout750 (.A(_1599_),
    .X(net750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout751 (.A(_1596_),
    .X(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout752 (.A(_1595_),
    .X(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout753 (.A(_1588_),
    .X(net753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout754 (.A(_1557_),
    .X(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout755 (.A(_1532_),
    .X(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout756 (.A(_1521_),
    .X(net756),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout757 (.A(_1517_),
    .X(net757),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout758 (.A(_1503_),
    .X(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout759 (.A(\sap_3_inst.controller.stage[2] ),
    .X(net759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout760 (.A(\sap_3_inst.controller.stage[1] ),
    .X(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout761 (.A(\sap_3_inst.controller.stage[0] ),
    .X(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout762 (.A(\sap_3_inst.alu.flags[1] ),
    .X(net762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout763 (.A(net764),
    .X(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout764 (.A(_1519_),
    .X(net764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout765 (.A(_1518_),
    .X(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout766 (.A(net767),
    .X(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout767 (.A(_1513_),
    .X(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout768 (.A(\sap_3_inst.controller.opcode[7] ),
    .X(net768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout769 (.A(\sap_3_inst.controller.opcode[7] ),
    .X(net769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout770 (.A(\sap_3_inst.controller.opcode[6] ),
    .X(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout771 (.A(\sap_3_inst.controller.opcode[6] ),
    .X(net771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout772 (.A(net773),
    .X(net772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout773 (.A(\sap_3_inst.controller.opcode[5] ),
    .X(net773),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout774 (.A(net775),
    .X(net774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout775 (.A(\sap_3_inst.controller.opcode[4] ),
    .X(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout776 (.A(net779),
    .X(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout777 (.A(net779),
    .X(net777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout778 (.A(net779),
    .X(net778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout779 (.A(\sap_3_inst.controller.opcode[3] ),
    .X(net779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout780 (.A(net781),
    .X(net780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout781 (.A(\sap_3_inst.controller.opcode[2] ),
    .X(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout782 (.A(net784),
    .X(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout783 (.A(net784),
    .X(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout784 (.A(\sap_3_inst.controller.opcode[1] ),
    .X(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout785 (.A(net786),
    .X(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout786 (.A(\sap_3_inst.controller.opcode[0] ),
    .X(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout787 (.A(net788),
    .X(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout788 (.A(net789),
    .X(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout789 (.A(\sap_3_inst.alu.acc[7] ),
    .X(net789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout790 (.A(net792),
    .X(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout791 (.A(net792),
    .X(net791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout792 (.A(\sap_3_inst.alu.acc[6] ),
    .X(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout793 (.A(net795),
    .X(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout794 (.A(net795),
    .X(net794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout795 (.A(\sap_3_inst.alu.acc[5] ),
    .X(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout796 (.A(net797),
    .X(net796),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout797 (.A(\sap_3_inst.alu.acc[4] ),
    .X(net797),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout798 (.A(net800),
    .X(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout799 (.A(net800),
    .X(net799),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout800 (.A(\sap_3_inst.alu.acc[3] ),
    .X(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout801 (.A(\sap_3_inst.alu.acc[2] ),
    .X(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout802 (.A(\sap_3_inst.alu.acc[2] ),
    .X(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout803 (.A(\sap_3_inst.alu.acc[1] ),
    .X(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout804 (.A(\sap_3_inst.alu.acc[1] ),
    .X(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout805 (.A(net806),
    .X(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout806 (.A(\sap_3_inst.alu.acc[0] ),
    .X(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout807 (.A(net808),
    .X(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout808 (.A(_1313_),
    .X(net808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout809 (.A(_1310_),
    .X(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout810 (.A(_1304_),
    .X(net810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout811 (.A(net812),
    .X(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout812 (.A(_1277_),
    .X(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout813 (.A(_0185_),
    .X(net813),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout814 (.A(net79),
    .X(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout815 (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .X(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout816 (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .X(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout817 (.A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[0] ),
    .X(net817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout818 (.A(net820),
    .X(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout819 (.A(net820),
    .X(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout820 (.A(net822),
    .X(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout821 (.A(net822),
    .X(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout822 (.A(rst_n),
    .X(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout823 (.A(net830),
    .X(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout824 (.A(net827),
    .X(net824),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout825 (.A(net827),
    .X(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout826 (.A(net827),
    .X(net826),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout827 (.A(net830),
    .X(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout828 (.A(net829),
    .X(net828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout829 (.A(net830),
    .X(net829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout830 (.A(rst_n),
    .X(net830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout831 (.A(net832),
    .X(net831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout832 (.A(net835),
    .X(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout833 (.A(net835),
    .X(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout834 (.A(net835),
    .X(net834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout835 (.A(net849),
    .X(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout836 (.A(net837),
    .X(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout837 (.A(net840),
    .X(net837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout838 (.A(net840),
    .X(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout839 (.A(net840),
    .X(net839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout840 (.A(net849),
    .X(net840),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout841 (.A(net842),
    .X(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout842 (.A(net845),
    .X(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout843 (.A(net844),
    .X(net843),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout844 (.A(net845),
    .X(net844),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout845 (.A(net849),
    .X(net845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout846 (.A(net847),
    .X(net846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout847 (.A(net848),
    .X(net847),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout848 (.A(net849),
    .X(net848),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout849 (.A(rst_n),
    .X(net849),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net31),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net32),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net33),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net34),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout31 (.A(net17),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout32 (.A(net21),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout33 (.A(net23),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout34 (.A(net24),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_template_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net35));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload1 (.VDD(VPWR),
    .A(clknet_3_1__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_1 clkload2 (.A(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload3 (.VDD(VPWR),
    .A(clknet_3_3__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload4 (.VDD(VPWR),
    .A(clknet_3_5__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload5 (.VDD(VPWR),
    .A(clknet_3_6__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload6 (.VDD(VPWR),
    .A(clknet_3_7__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk_div_out (.A(clk_div_out),
    .X(clknet_0_clk_div_out),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_clk_div_out (.A(clknet_0_clk_div_out),
    .X(clknet_1_0__leaf_clk_div_out),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_1__f_clk_div_out (.A(clknet_0_clk_div_out),
    .X(clknet_1_1__leaf_clk_div_out),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload7 (.A(clknet_1_1__leaf_clk_div_out),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_leaf_0_sap_3_inst.alu.clk  (.A(\clknet_1_0__leaf_sap_3_inst.alu.clk ),
    .X(\clknet_leaf_0_sap_3_inst.alu.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_leaf_1_sap_3_inst.alu.clk  (.A(\clknet_1_1__leaf_sap_3_inst.alu.clk ),
    .X(\clknet_leaf_1_sap_3_inst.alu.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_leaf_2_sap_3_inst.alu.clk  (.A(\clknet_1_0__leaf_sap_3_inst.alu.clk ),
    .X(\clknet_leaf_2_sap_3_inst.alu.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_0_sap_3_inst.alu.clk  (.A(\sap_3_inst.alu.clk ),
    .X(\clknet_0_sap_3_inst.alu.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_1_0__f_sap_3_inst.alu.clk  (.A(\clknet_0_sap_3_inst.alu.clk ),
    .X(\clknet_1_0__leaf_sap_3_inst.alu.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_1_1__f_sap_3_inst.alu.clk  (.A(\clknet_0_sap_3_inst.alu.clk ),
    .X(\clknet_1_1__leaf_sap_3_inst.alu.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload8 (.A(\clknet_1_1__leaf_sap_3_inst.alu.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_0_sap_3_inst.alu.clk_regs  (.A(\sap_3_inst.alu.clk_regs ),
    .X(\clknet_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_0_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_0_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_1_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_1_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_2_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_2_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_3_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_3_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_4_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_4_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_5_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_5_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_6_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_6_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_7_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_7_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_8_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_8_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_9_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_9_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_10_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_10_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_11_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_11_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_12_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_12_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_13_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_13_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_14_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_14_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_15_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_15_0_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_0__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_0_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_1__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_0_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_2__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_1_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_3__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_1_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_4__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_2_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_5__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_2_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_6__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_3_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_7__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_3_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_8__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_4_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_9__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_4_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_10__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_5_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_11__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_5_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_12__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_6_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_13__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_6_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_14__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_7_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_15__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_7_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_16__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_8_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_17__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_8_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_18__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_9_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_19__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_9_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_20__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_10_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_21__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_10_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_22__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_11_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_23__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_11_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_24__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_12_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_25__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_12_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_26__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_13_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_27__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_13_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_28__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_14_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_29__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_14_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_30__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_15_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_31__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_15_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload9 (.VDD(VPWR),
    .A(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload10 (.VDD(VPWR),
    .A(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload11 (.VDD(VPWR),
    .A(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload12 (.VDD(VPWR),
    .A(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload13 (.VDD(VPWR),
    .A(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload14 (.VDD(VPWR),
    .A(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ),
    .VSS(VGND));
 sg13g2_buf_1 clkload15 (.A(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload16 (.VDD(VPWR),
    .A(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ),
    .VSS(VGND));
 sg13g2_buf_1 clkload17 (.A(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload18 (.VDD(VPWR),
    .A(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload19 (.VDD(VPWR),
    .A(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold2 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold3 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold4 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold5 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold6 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold7 (.A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0157_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_ser.shadow_reg[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_ser.shadow_reg[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold11 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_ser.state[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0195_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold14 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u_ser.shadow_reg[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_ser.shadow_reg[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold17 (.A(\u_ser.shadow_reg[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_ser.shadow_reg[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_ser.shadow_reg[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold20 (.A(\u_ser.shadow_reg[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_ser.bit_pos[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold22 (.A(regFile_serial),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold23 (.A(sap_3_outputReg_start_sync),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0188_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold25 (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold26 (.A(\sap_3_inst.reg_file.array_serializer_inst.state[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0159_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold28 (.A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold29 (.A(sap_3_outputReg_serial),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold30 (.A(\u_ser.bit_pos[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net79));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_1027 (.VDD(VPWR),
    .VSS(VGND));
 assign uo_out[6] = net35;
 assign uo_out[7] = net36;
endmodule
