* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_lgcp_1 abstract view
.subckt sg13g2_lgcp_1 GATE CLK GCLK VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
X_3155_ _0690_ _1569_ _0275_ _0691_ VPWR VGND sg13g2_a21o_2
XFILLER_28_918 VPWR VGND sg13g2_decap_8
X_3086_ VGND VPWR _0611_ _0621_ _0622_ _0275_ sg13g2_a21oi_1
X_2106_ net719 net718 _1527_ VPWR VGND sg13g2_and2_1
XFILLER_36_962 VPWR VGND sg13g2_decap_8
X_2037_ _1460_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[0\] VPWR VGND
+ sg13g2_inv_2
XFILLER_23_612 VPWR VGND sg13g2_decap_8
XFILLER_22_122 VPWR VGND sg13g2_fill_2
X_3988_ _1406_ VPWR _0184_ VGND net548 _1405_ sg13g2_o21ai_1
XFILLER_23_689 VPWR VGND sg13g2_decap_8
X_2939_ VGND VPWR _0472_ _0501_ _0502_ _0500_ sg13g2_a21oi_1
XFILLER_19_929 VPWR VGND sg13g2_decap_8
XFILLER_46_759 VPWR VGND sg13g2_decap_8
XFILLER_45_214 VPWR VGND sg13g2_fill_1
XFILLER_26_450 VPWR VGND sg13g2_decap_8
XFILLER_27_984 VPWR VGND sg13g2_decap_8
XFILLER_42_965 VPWR VGND sg13g2_decap_8
XFILLER_14_656 VPWR VGND sg13g2_decap_8
XFILLER_13_155 VPWR VGND sg13g2_fill_2
XFILLER_41_486 VPWR VGND sg13g2_decap_8
XFILLER_6_855 VPWR VGND sg13g2_decap_8
XFILLER_10_895 VPWR VGND sg13g2_decap_8
XFILLER_3_23 VPWR VGND sg13g2_decap_8
XFILLER_49_542 VPWR VGND sg13g2_decap_8
XFILLER_3_1018 VPWR VGND sg13g2_decap_8
XFILLER_37_737 VPWR VGND sg13g2_decap_8
XFILLER_33_921 VPWR VGND sg13g2_decap_8
X_3911_ _1346_ _1347_ _1345_ _1349_ VPWR VGND _1348_ sg13g2_nand4_1
X_3842_ _1287_ net63 _1281_ VPWR VGND sg13g2_nand2_1
XFILLER_20_604 VPWR VGND sg13g2_decap_8
XFILLER_33_998 VPWR VGND sg13g2_decap_8
XFILLER_32_497 VPWR VGND sg13g2_decap_8
X_3773_ net14 net598 _1239_ _1240_ VPWR VGND sg13g2_nor3_1
X_2724_ net57 sap_3_inst.out\[3\] net766 _0021_ VPWR VGND sg13g2_mux2_1
X_2655_ net754 net744 net756 net746 _0249_ VPWR VGND sg13g2_nor4_1
X_2586_ _1988_ VPWR _1997_ VGND net567 _1996_ sg13g2_o21ai_1
XFILLER_28_715 VPWR VGND sg13g2_decap_8
X_4187_ net794 VGND VPWR _0165_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[3\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
X_3207_ _0743_ _1460_ net615 VPWR VGND sg13g2_nand2_1
X_3138_ _0614_ _0628_ net680 _0674_ VPWR VGND sg13g2_nand3_1
X_3069_ _0604_ VPWR _0605_ VGND _1607_ _0600_ sg13g2_o21ai_1
XFILLER_23_431 VPWR VGND sg13g2_decap_8
XFILLER_24_932 VPWR VGND sg13g2_decap_8
XFILLER_11_648 VPWR VGND sg13g2_decap_8
XFILLER_23_486 VPWR VGND sg13g2_decap_8
XFILLER_7_608 VPWR VGND sg13g2_decap_8
XFILLER_3_836 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
Xfanout650 _0729_ net650 VPWR VGND sg13g2_buf_8
Xfanout672 _1947_ net672 VPWR VGND sg13g2_buf_8
Xfanout683 _1714_ net683 VPWR VGND sg13g2_buf_1
Xfanout694 _1530_ net694 VPWR VGND sg13g2_buf_8
Xfanout661 _0625_ net661 VPWR VGND sg13g2_buf_2
XFILLER_19_726 VPWR VGND sg13g2_decap_8
XFILLER_46_556 VPWR VGND sg13g2_decap_8
XFILLER_27_781 VPWR VGND sg13g2_decap_8
XFILLER_34_718 VPWR VGND sg13g2_decap_8
XFILLER_42_762 VPWR VGND sg13g2_decap_8
XFILLER_15_976 VPWR VGND sg13g2_decap_8
XFILLER_30_913 VPWR VGND sg13g2_decap_8
XFILLER_6_652 VPWR VGND sg13g2_decap_8
XFILLER_5_140 VPWR VGND sg13g2_fill_2
XFILLER_10_692 VPWR VGND sg13g2_decap_8
X_2440_ _1859_ net620 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] net634
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2371_ _1772_ _1790_ _1792_ VPWR VGND sg13g2_nor2_1
X_4110_ net776 VGND VPWR _0088_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\]
+ clknet_5_9__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4041_ net788 VGND VPWR _0023_ u_ser.shadow_reg\[5\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_37_534 VPWR VGND sg13g2_decap_8
XFILLER_33_795 VPWR VGND sg13g2_decap_8
XFILLER_21_968 VPWR VGND sg13g2_decap_8
X_3825_ net15 net605 _1117_ _1275_ VPWR VGND sg13g2_nor3_1
X_3756_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] _1226_ net655 _0132_
+ VPWR VGND sg13g2_mux2_1
X_2707_ _0286_ _1653_ _0285_ VPWR VGND sg13g2_nand2_1
X_3687_ _1040_ _1041_ _1181_ _1183_ VPWR VGND sg13g2_nor3_1
X_2638_ _0233_ net625 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] _1799_
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_0_806 VPWR VGND sg13g2_decap_8
X_2569_ _1980_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] net634
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_28_512 VPWR VGND sg13g2_decap_8
XFILLER_16_718 VPWR VGND sg13g2_decap_8
XFILLER_28_589 VPWR VGND sg13g2_decap_8
XFILLER_43_537 VPWR VGND sg13g2_decap_8
XFILLER_12_924 VPWR VGND sg13g2_decap_8
XFILLER_3_633 VPWR VGND sg13g2_decap_8
XFILLER_2_143 VPWR VGND sg13g2_fill_1
XFILLER_19_523 VPWR VGND sg13g2_decap_8
XFILLER_47_843 VPWR VGND sg13g2_decap_8
XFILLER_0_57 VPWR VGND sg13g2_decap_8
XFILLER_34_515 VPWR VGND sg13g2_decap_8
XFILLER_15_773 VPWR VGND sg13g2_decap_8
XFILLER_14_283 VPWR VGND sg13g2_fill_1
XFILLER_30_710 VPWR VGND sg13g2_decap_8
XFILLER_30_787 VPWR VGND sg13g2_decap_8
XFILLER_31_1023 VPWR VGND sg13g2_decap_4
X_3610_ VPWR VGND _1122_ net661 _1121_ net666 _1123_ _1027_ sg13g2_a221oi_1
X_3541_ net22 _1063_ _1064_ VPWR VGND sg13g2_nor2_1
XFILLER_7_972 VPWR VGND sg13g2_decap_8
X_3472_ net575 _1001_ _1002_ VPWR VGND sg13g2_nor2_2
XFILLER_9_1013 VPWR VGND sg13g2_decap_8
X_2423_ VPWR VGND _1842_ _1715_ _1841_ net689 _1844_ _1743_ sg13g2_a221oi_1
X_2354_ _1774_ net697 net682 _1775_ VPWR VGND sg13g2_a21o_1
XFILLER_29_0 VPWR VGND sg13g2_fill_1
X_2285_ VPWR VGND net724 _1571_ _1705_ _1586_ _1706_ _1604_ sg13g2_a221oi_1
X_4024_ _0196_ _1434_ _1431_ _1433_ net58 VPWR VGND sg13g2_a22oi_1
XFILLER_38_865 VPWR VGND sg13g2_decap_8
XFILLER_25_548 VPWR VGND sg13g2_decap_8
XFILLER_40_529 VPWR VGND sg13g2_decap_8
XFILLER_21_765 VPWR VGND sg13g2_decap_8
XFILLER_33_592 VPWR VGND sg13g2_decap_8
X_3808_ net604 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] _1262_ _0148_
+ VPWR VGND sg13g2_a21o_1
X_3739_ _1215_ VPWR _0126_ VGND _1442_ _1211_ sg13g2_o21ai_1
XFILLER_0_603 VPWR VGND sg13g2_decap_8
XFILLER_29_832 VPWR VGND sg13g2_decap_8
XFILLER_16_515 VPWR VGND sg13g2_decap_8
XFILLER_18_64 VPWR VGND sg13g2_fill_1
XFILLER_28_375 VPWR VGND sg13g2_fill_1
XFILLER_44_857 VPWR VGND sg13g2_decap_8
XFILLER_12_721 VPWR VGND sg13g2_decap_8
XFILLER_15_1018 VPWR VGND sg13g2_decap_8
XFILLER_7_213 VPWR VGND sg13g2_fill_2
XFILLER_11_275 VPWR VGND sg13g2_fill_2
XFILLER_12_798 VPWR VGND sg13g2_decap_8
XFILLER_8_769 VPWR VGND sg13g2_decap_8
XFILLER_4_964 VPWR VGND sg13g2_decap_8
XFILLER_39_607 VPWR VGND sg13g2_decap_8
XFILLER_47_640 VPWR VGND sg13g2_decap_8
X_2070_ VPWR _1493_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_35_835 VPWR VGND sg13g2_decap_8
XFILLER_34_345 VPWR VGND sg13g2_fill_2
XFILLER_15_570 VPWR VGND sg13g2_decap_8
X_2972_ VGND VPWR net745 net672 _0534_ _0502_ sg13g2_a21oi_1
XFILLER_30_584 VPWR VGND sg13g2_decap_8
X_3524_ net575 _0906_ _1050_ VPWR VGND sg13g2_nor2_2
X_3455_ _0766_ VPWR _0986_ VGND net559 _0853_ sg13g2_o21ai_1
X_2406_ _1826_ _1827_ VPWR VGND sg13g2_inv_4
X_3386_ net560 _0918_ _0919_ VPWR VGND sg13g2_nor2_1
X_2337_ _1758_ _1682_ _1757_ VPWR VGND sg13g2_nand2_1
X_2268_ net707 VPWR _1689_ VGND _1687_ _1688_ sg13g2_o21ai_1
XFILLER_29_128 VPWR VGND sg13g2_fill_2
X_4007_ _1422_ VPWR _1423_ VGND net77 _0187_ sg13g2_o21ai_1
XFILLER_38_662 VPWR VGND sg13g2_decap_8
X_2199_ _1437_ net730 _1620_ VPWR VGND sg13g2_nor2_2
XFILLER_26_835 VPWR VGND sg13g2_decap_8
XFILLER_25_389 VPWR VGND sg13g2_fill_1
XFILLER_21_562 VPWR VGND sg13g2_decap_8
XFILLER_1_912 VPWR VGND sg13g2_decap_8
XFILLER_49_927 VPWR VGND sg13g2_decap_8
Xhold30 sap_3_outputReg_serial VPWR VGND net77 sg13g2_dlygate4sd3_1
XFILLER_0_477 VPWR VGND sg13g2_decap_8
XFILLER_1_989 VPWR VGND sg13g2_decap_8
XFILLER_48_437 VPWR VGND sg13g2_decap_8
XFILLER_35_109 VPWR VGND sg13g2_fill_2
XFILLER_17_857 VPWR VGND sg13g2_decap_8
XFILLER_44_654 VPWR VGND sg13g2_decap_8
XFILLER_32_805 VPWR VGND sg13g2_decap_8
XFILLER_40_893 VPWR VGND sg13g2_decap_8
XFILLER_12_595 VPWR VGND sg13g2_decap_8
XFILLER_8_566 VPWR VGND sg13g2_decap_8
XFILLER_4_761 VPWR VGND sg13g2_decap_8
X_3240_ _0772_ _0773_ _0770_ _0776_ VPWR VGND _0774_ sg13g2_nand4_1
XFILLER_6_1027 VPWR VGND sg13g2_fill_2
XFILLER_6_1016 VPWR VGND sg13g2_decap_8
X_3171_ VGND VPWR net697 _1614_ _0707_ net682 sg13g2_a21oi_1
X_2122_ _1543_ net725 net727 VPWR VGND sg13g2_nand2b_1
X_2053_ VPWR _1476_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] VGND
+ sg13g2_inv_1
XFILLER_35_632 VPWR VGND sg13g2_decap_8
X_2955_ _0492_ _0516_ _0518_ VPWR VGND sg13g2_nor2_1
X_2886_ _0451_ _0426_ _0450_ VPWR VGND sg13g2_nand2_1
X_3507_ net562 sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[7\] _1035_ _0074_
+ VPWR VGND sg13g2_a21o_1
XFILLER_44_1011 VPWR VGND sg13g2_decap_8
X_3438_ _0967_ _0968_ _0969_ VPWR VGND sg13g2_and2_1
X_3369_ net11 net571 _0903_ VPWR VGND sg13g2_nor2_1
XFILLER_39_971 VPWR VGND sg13g2_decap_8
XFILLER_45_429 VPWR VGND sg13g2_decap_8
XFILLER_26_632 VPWR VGND sg13g2_decap_8
XFILLER_38_470 VPWR VGND sg13g2_fill_1
XFILLER_25_120 VPWR VGND sg13g2_fill_2
XFILLER_14_838 VPWR VGND sg13g2_decap_8
XFILLER_25_153 VPWR VGND sg13g2_fill_1
XFILLER_41_668 VPWR VGND sg13g2_decap_8
X_4025__3 VPWR net37 clknet_leaf_2_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_5_558 VPWR VGND sg13g2_decap_8
Xoutput20 net20 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_49_724 VPWR VGND sg13g2_decap_8
XFILLER_1_786 VPWR VGND sg13g2_decap_8
XFILLER_37_919 VPWR VGND sg13g2_decap_8
XFILLER_17_654 VPWR VGND sg13g2_decap_8
XFILLER_45_996 VPWR VGND sg13g2_decap_8
XFILLER_44_451 VPWR VGND sg13g2_decap_8
XFILLER_16_164 VPWR VGND sg13g2_fill_1
XFILLER_32_602 VPWR VGND sg13g2_decap_8
XFILLER_32_679 VPWR VGND sg13g2_decap_8
XFILLER_40_690 VPWR VGND sg13g2_decap_8
XFILLER_9_831 VPWR VGND sg13g2_decap_8
X_2740_ net713 _0306_ _0308_ _0309_ VPWR VGND sg13g2_or3_1
XFILLER_31_189 VPWR VGND sg13g2_fill_2
X_2671_ _0263_ _1569_ _1786_ VPWR VGND sg13g2_nand2b_1
X_3223_ _0759_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] net655 VPWR
+ VGND sg13g2_nand2_1
XFILLER_39_212 VPWR VGND sg13g2_fill_2
X_3154_ _0674_ VPWR _0690_ VGND _0683_ _0689_ sg13g2_o21ai_1
X_3085_ _0263_ _0617_ _0619_ _0620_ _0621_ VPWR VGND sg13g2_nor4_1
X_2105_ _1525_ VPWR _1526_ VGND _1509_ _1515_ sg13g2_o21ai_1
X_2036_ VPWR _1459_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] VGND
+ sg13g2_inv_1
XFILLER_36_941 VPWR VGND sg13g2_decap_8
X_3987_ _1406_ sap_3_inst.alu.act\[6\] net548 VPWR VGND sg13g2_nand2_1
XFILLER_23_668 VPWR VGND sg13g2_decap_8
X_2938_ _0471_ VPWR _0501_ VGND net747 net671 sg13g2_o21ai_1
X_2869_ _0323_ _0431_ _0435_ VPWR VGND sg13g2_nor2_1
XFILLER_2_539 VPWR VGND sg13g2_decap_8
XFILLER_19_908 VPWR VGND sg13g2_decap_8
XFILLER_46_738 VPWR VGND sg13g2_decap_8
XFILLER_27_963 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_42_944 VPWR VGND sg13g2_decap_8
XFILLER_14_635 VPWR VGND sg13g2_decap_8
XFILLER_41_465 VPWR VGND sg13g2_decap_8
XFILLER_13_167 VPWR VGND sg13g2_fill_1
XFILLER_6_834 VPWR VGND sg13g2_decap_8
XFILLER_5_311 VPWR VGND sg13g2_fill_2
XFILLER_10_874 VPWR VGND sg13g2_decap_8
XFILLER_47_9 VPWR VGND sg13g2_fill_1
XFILLER_3_13 VPWR VGND sg13g2_fill_1
XFILLER_49_521 VPWR VGND sg13g2_decap_8
XFILLER_1_583 VPWR VGND sg13g2_decap_8
XFILLER_37_716 VPWR VGND sg13g2_decap_8
XFILLER_49_598 VPWR VGND sg13g2_decap_8
XFILLER_17_462 VPWR VGND sg13g2_fill_1
XFILLER_18_985 VPWR VGND sg13g2_decap_8
XFILLER_33_900 VPWR VGND sg13g2_decap_8
XFILLER_45_793 VPWR VGND sg13g2_decap_8
X_3910_ _1348_ _1306_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] _1302_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_977 VPWR VGND sg13g2_decap_8
X_3841_ VGND VPWR net769 _0156_ _1286_ net72 sg13g2_a21oi_1
X_3772_ net574 _1238_ _1239_ VPWR VGND sg13g2_nor2_1
X_2723_ net62 sap_3_inst.out\[2\] net766 _0020_ VPWR VGND sg13g2_mux2_1
X_2654_ _1566_ _1940_ _0248_ VPWR VGND sg13g2_nor2_1
X_2585_ _1991_ _1995_ _1996_ VPWR VGND sg13g2_nor2_1
XFILLER_41_1025 VPWR VGND sg13g2_decap_4
X_4186_ net793 VGND VPWR _0164_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[2\]
+ clknet_3_3__leaf_clk sg13g2_dfrbpq_1
X_3206_ _0741_ VPWR _0742_ VGND _1461_ net590 sg13g2_o21ai_1
X_3137_ _0673_ _0658_ _0670_ VPWR VGND sg13g2_nand2_1
XFILLER_27_226 VPWR VGND sg13g2_fill_2
XFILLER_43_719 VPWR VGND sg13g2_decap_8
X_3068_ _1601_ VPWR _0604_ VGND _1581_ _1626_ sg13g2_o21ai_1
XFILLER_24_911 VPWR VGND sg13g2_decap_8
X_2019_ VPWR _1442_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_35_281 VPWR VGND sg13g2_fill_1
XFILLER_23_465 VPWR VGND sg13g2_decap_8
XFILLER_24_988 VPWR VGND sg13g2_decap_8
XFILLER_11_627 VPWR VGND sg13g2_decap_8
XFILLER_12_33 VPWR VGND sg13g2_fill_2
XFILLER_3_815 VPWR VGND sg13g2_decap_8
Xfanout651 net652 net651 VPWR VGND sg13g2_buf_8
Xfanout640 net642 net640 VPWR VGND sg13g2_buf_8
Xfanout673 _0260_ net673 VPWR VGND sg13g2_buf_8
Xfanout684 _1674_ net684 VPWR VGND sg13g2_buf_8
XFILLER_19_705 VPWR VGND sg13g2_decap_8
Xfanout662 _1746_ net662 VPWR VGND sg13g2_buf_8
Xfanout695 _1530_ net695 VPWR VGND sg13g2_buf_8
XFILLER_46_535 VPWR VGND sg13g2_decap_8
XFILLER_18_226 VPWR VGND sg13g2_fill_2
XFILLER_27_760 VPWR VGND sg13g2_decap_8
XFILLER_42_741 VPWR VGND sg13g2_decap_8
XFILLER_14_421 VPWR VGND sg13g2_fill_2
XFILLER_15_955 VPWR VGND sg13g2_decap_8
XFILLER_18_1027 VPWR VGND sg13g2_fill_2
XFILLER_30_969 VPWR VGND sg13g2_decap_8
XFILLER_10_671 VPWR VGND sg13g2_decap_8
XFILLER_6_631 VPWR VGND sg13g2_decap_8
X_2370_ VPWR _1791_ _1790_ VGND sg13g2_inv_1
X_4040_ net788 VGND VPWR _0022_ u_ser.shadow_reg\[4\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_37_513 VPWR VGND sg13g2_decap_8
XFILLER_49_395 VPWR VGND sg13g2_decap_8
XFILLER_24_218 VPWR VGND sg13g2_fill_2
XFILLER_45_590 VPWR VGND sg13g2_decap_8
XFILLER_18_782 VPWR VGND sg13g2_decap_8
XFILLER_32_240 VPWR VGND sg13g2_fill_1
XFILLER_33_774 VPWR VGND sg13g2_decap_8
XFILLER_21_947 VPWR VGND sg13g2_decap_8
X_3824_ _1270_ VPWR _0152_ VGND _1271_ _1274_ sg13g2_o21ai_1
XFILLER_20_457 VPWR VGND sg13g2_fill_1
X_3755_ _1224_ _1225_ _1226_ VPWR VGND _1144_ sg13g2_nand3b_1
X_2706_ VGND VPWR _1616_ _0284_ _0285_ net696 sg13g2_a21oi_1
X_3686_ _1182_ net569 VPWR VGND net647 sg13g2_nand2b_2
X_2637_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] net639
+ net622 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] _0232_ net678 sg13g2_a221oi_1
X_2568_ _1979_ net620 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] net626
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2499_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] net621
+ net638 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] _1914_ net677 sg13g2_a221oi_1
X_4169_ net795 VGND VPWR _0147_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\]
+ clknet_5_29__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_43_516 VPWR VGND sg13g2_decap_8
XFILLER_28_568 VPWR VGND sg13g2_decap_8
XFILLER_12_903 VPWR VGND sg13g2_decap_8
XFILLER_24_785 VPWR VGND sg13g2_decap_8
Xclkbuf_4_12_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_12_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_7_439 VPWR VGND sg13g2_fill_1
XFILLER_23_98 VPWR VGND sg13g2_fill_1
XFILLER_3_612 VPWR VGND sg13g2_decap_8
XFILLER_2_122 VPWR VGND sg13g2_decap_4
XFILLER_3_689 VPWR VGND sg13g2_decap_8
XFILLER_47_822 VPWR VGND sg13g2_decap_8
XFILLER_19_502 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_47_899 VPWR VGND sg13g2_decap_8
XFILLER_0_36 VPWR VGND sg13g2_decap_8
XFILLER_19_579 VPWR VGND sg13g2_decap_8
XFILLER_15_752 VPWR VGND sg13g2_decap_8
XFILLER_30_766 VPWR VGND sg13g2_decap_8
XFILLER_31_1002 VPWR VGND sg13g2_decap_8
X_3540_ net583 _0975_ _1063_ VPWR VGND sg13g2_nor2_2
XFILLER_7_951 VPWR VGND sg13g2_decap_8
XFILLER_11_991 VPWR VGND sg13g2_decap_8
X_3471_ _1000_ VPWR _1001_ VGND net560 _0855_ sg13g2_o21ai_1
X_2422_ _1843_ net689 _1743_ VPWR VGND sg13g2_nand2_1
X_2353_ _1436_ _1563_ _1774_ VPWR VGND sg13g2_nor2_2
X_2284_ _1584_ net708 _1703_ _1705_ VPWR VGND sg13g2_nor3_1
X_4023_ net767 _1410_ u_ser.bit_pos\[1\] _1431_ VPWR VGND sg13g2_nand3_1
XFILLER_38_844 VPWR VGND sg13g2_decap_8
XFILLER_25_527 VPWR VGND sg13g2_decap_8
XFILLER_40_508 VPWR VGND sg13g2_decap_8
XFILLER_33_571 VPWR VGND sg13g2_decap_8
XFILLER_21_744 VPWR VGND sg13g2_decap_8
X_3807_ VPWR VGND _1261_ net603 _0884_ net577 _1262_ _0874_ sg13g2_a221oi_1
X_3738_ _1055_ _1211_ _1054_ _1215_ VPWR VGND sg13g2_nand3_1
X_3669_ VGND VPWR net581 _0999_ _1167_ net597 sg13g2_a21oi_1
Xclkbuf_4_4_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_4_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_0_659 VPWR VGND sg13g2_decap_8
XFILLER_48_619 VPWR VGND sg13g2_decap_8
XFILLER_29_811 VPWR VGND sg13g2_decap_8
XFILLER_29_888 VPWR VGND sg13g2_decap_8
XFILLER_44_836 VPWR VGND sg13g2_decap_8
XFILLER_12_700 VPWR VGND sg13g2_decap_8
XFILLER_24_582 VPWR VGND sg13g2_decap_8
XFILLER_31_519 VPWR VGND sg13g2_decap_8
XFILLER_34_75 VPWR VGND sg13g2_fill_2
XFILLER_12_777 VPWR VGND sg13g2_decap_8
XFILLER_8_748 VPWR VGND sg13g2_decap_8
XFILLER_4_943 VPWR VGND sg13g2_decap_8
XFILLER_3_486 VPWR VGND sg13g2_decap_8
XFILLER_19_365 VPWR VGND sg13g2_fill_1
XFILLER_35_814 VPWR VGND sg13g2_decap_8
XFILLER_47_696 VPWR VGND sg13g2_decap_8
XFILLER_46_173 VPWR VGND sg13g2_fill_2
XFILLER_43_880 VPWR VGND sg13g2_decap_8
X_2971_ net542 net617 _0533_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_519 VPWR VGND sg13g2_decap_8
XFILLER_30_563 VPWR VGND sg13g2_decap_8
X_3523_ net19 _1048_ _1049_ VPWR VGND sg13g2_nor2_2
X_3454_ VGND VPWR net578 _0983_ _0985_ net562 sg13g2_a21oi_1
XFILLER_41_0 VPWR VGND sg13g2_fill_1
X_2405_ VGND VPWR _1515_ _1825_ _1826_ _1813_ sg13g2_a21oi_1
X_3385_ _0872_ _0895_ _0857_ _0918_ VPWR VGND _0917_ sg13g2_nand4_1
X_2336_ _1757_ net696 net706 VPWR VGND sg13g2_nand2_1
X_2267_ VGND VPWR _1688_ _1638_ _1577_ sg13g2_or2_1
XFILLER_38_641 VPWR VGND sg13g2_decap_8
X_4006_ _1418_ _1420_ _0187_ _1422_ VPWR VGND _1421_ sg13g2_nand4_1
XFILLER_26_814 VPWR VGND sg13g2_decap_8
X_2198_ _1619_ net680 _1586_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_1019 VPWR VGND sg13g2_decap_8
XFILLER_21_541 VPWR VGND sg13g2_decap_8
XFILLER_49_906 VPWR VGND sg13g2_decap_8
XFILLER_1_968 VPWR VGND sg13g2_decap_8
XFILLER_48_416 VPWR VGND sg13g2_decap_8
Xhold31 sap_3_inst.reg_file.array_serializer_inst.word_index\[3\] VPWR VGND net78
+ sg13g2_dlygate4sd3_1
XFILLER_0_456 VPWR VGND sg13g2_decap_8
XFILLER_29_53 VPWR VGND sg13g2_fill_2
Xhold20 _0161_ VPWR VGND net67 sg13g2_dlygate4sd3_1
XFILLER_44_633 VPWR VGND sg13g2_decap_8
XFILLER_17_836 VPWR VGND sg13g2_decap_8
XFILLER_29_685 VPWR VGND sg13g2_decap_8
XFILLER_45_41 VPWR VGND sg13g2_fill_2
XFILLER_16_368 VPWR VGND sg13g2_fill_1
XFILLER_25_891 VPWR VGND sg13g2_decap_8
XFILLER_40_872 VPWR VGND sg13g2_decap_8
XFILLER_8_545 VPWR VGND sg13g2_decap_8
XFILLER_12_574 VPWR VGND sg13g2_decap_8
XFILLER_6_57 VPWR VGND sg13g2_fill_2
XFILLER_4_740 VPWR VGND sg13g2_decap_8
X_3170_ _0696_ _0701_ _0703_ _0705_ _0706_ VPWR VGND sg13g2_nor4_1
X_2121_ _1439_ net727 _1542_ VPWR VGND sg13g2_nor2_1
X_2052_ _1475_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[5\] VPWR VGND
+ sg13g2_inv_2
XFILLER_48_983 VPWR VGND sg13g2_decap_8
XFILLER_35_611 VPWR VGND sg13g2_decap_8
XFILLER_47_493 VPWR VGND sg13g2_decap_8
XFILLER_35_688 VPWR VGND sg13g2_decap_8
X_2954_ _0492_ _0516_ _0517_ VPWR VGND sg13g2_and2_1
X_2885_ _0450_ _0447_ _0448_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_883 VPWR VGND sg13g2_decap_8
X_3506_ VPWR VGND _1034_ net562 _1030_ _1022_ _1035_ _1026_ sg13g2_a221oi_1
X_3437_ _0968_ _1475_ net612 VPWR VGND sg13g2_nand2_1
X_3368_ net19 _0838_ _0902_ VPWR VGND sg13g2_nor2_1
X_2319_ VPWR _1740_ _1739_ VGND sg13g2_inv_1
XFILLER_45_408 VPWR VGND sg13g2_decap_8
Xheichips25_template_33 VPWR VGND uo_out[6] sg13g2_tielo
X_3299_ VGND VPWR _1569_ _0834_ _0835_ _0275_ sg13g2_a21oi_1
XFILLER_39_950 VPWR VGND sg13g2_decap_8
XFILLER_26_611 VPWR VGND sg13g2_decap_8
XFILLER_14_817 VPWR VGND sg13g2_decap_8
XFILLER_26_688 VPWR VGND sg13g2_decap_8
XFILLER_41_647 VPWR VGND sg13g2_decap_8
XFILLER_40_146 VPWR VGND sg13g2_fill_2
XFILLER_21_360 VPWR VGND sg13g2_fill_1
XFILLER_22_883 VPWR VGND sg13g2_decap_8
XFILLER_5_537 VPWR VGND sg13g2_decap_8
XFILLER_31_76 VPWR VGND sg13g2_fill_2
Xoutput21 net21 uio_out[4] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_oe[1] VPWR VGND sg13g2_buf_1
XFILLER_49_703 VPWR VGND sg13g2_decap_8
XFILLER_1_765 VPWR VGND sg13g2_decap_8
Xclkbuf_5_6__f_sap_3_inst.alu.clk_regs clknet_4_3_0_sap_3_inst.alu.clk_regs clknet_5_6__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_29_482 VPWR VGND sg13g2_decap_8
XFILLER_44_430 VPWR VGND sg13g2_decap_8
XFILLER_17_633 VPWR VGND sg13g2_decap_8
XFILLER_45_975 VPWR VGND sg13g2_decap_8
XFILLER_31_113 VPWR VGND sg13g2_fill_2
XFILLER_32_658 VPWR VGND sg13g2_decap_8
XFILLER_9_810 VPWR VGND sg13g2_decap_8
XFILLER_13_894 VPWR VGND sg13g2_decap_8
X_2670_ VGND VPWR net673 _0261_ _0262_ net708 sg13g2_a21oi_1
XFILLER_9_887 VPWR VGND sg13g2_decap_8
X_3222_ _0758_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] net606 VPWR
+ VGND sg13g2_nand2_1
X_3153_ _0685_ _0688_ _0689_ VPWR VGND net680 sg13g2_nand3b_1
X_2104_ _1518_ _1520_ _1516_ _1525_ VPWR VGND _1522_ sg13g2_nand4_1
XFILLER_48_780 VPWR VGND sg13g2_decap_8
X_3084_ VGND VPWR _0616_ _0618_ _0620_ _1703_ sg13g2_a21oi_1
XFILLER_27_419 VPWR VGND sg13g2_fill_2
XFILLER_36_920 VPWR VGND sg13g2_decap_8
X_2035_ VPWR _1458_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] VGND
+ sg13g2_inv_1
XFILLER_36_997 VPWR VGND sg13g2_decap_8
XFILLER_23_647 VPWR VGND sg13g2_decap_8
XFILLER_11_809 VPWR VGND sg13g2_decap_8
X_3986_ VGND VPWR net746 net663 _1405_ _1404_ sg13g2_a21oi_1
X_2937_ _0500_ net745 net671 VPWR VGND sg13g2_xnor2_1
XFILLER_31_680 VPWR VGND sg13g2_decap_8
X_2868_ _0428_ VPWR _0434_ VGND net564 _0433_ sg13g2_o21ai_1
X_2799_ _0367_ _0355_ _0320_ VPWR VGND sg13g2_nand2b_1
XFILLER_2_518 VPWR VGND sg13g2_decap_8
Xfanout800 net801 net800 VPWR VGND sg13g2_buf_8
Xclkbuf_5_13__f_sap_3_inst.alu.clk_regs clknet_4_6_0_sap_3_inst.alu.clk_regs clknet_5_13__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_46_717 VPWR VGND sg13g2_decap_8
XFILLER_27_942 VPWR VGND sg13g2_decap_8
XFILLER_42_923 VPWR VGND sg13g2_decap_8
XFILLER_14_614 VPWR VGND sg13g2_decap_8
XFILLER_41_422 VPWR VGND sg13g2_fill_2
XFILLER_26_485 VPWR VGND sg13g2_decap_8
XFILLER_22_680 VPWR VGND sg13g2_decap_8
XFILLER_10_853 VPWR VGND sg13g2_decap_8
XFILLER_6_813 VPWR VGND sg13g2_decap_8
XFILLER_49_500 VPWR VGND sg13g2_decap_8
XFILLER_1_562 VPWR VGND sg13g2_decap_8
XFILLER_3_58 VPWR VGND sg13g2_fill_2
XFILLER_49_577 VPWR VGND sg13g2_decap_8
XFILLER_18_964 VPWR VGND sg13g2_decap_8
XFILLER_45_772 VPWR VGND sg13g2_decap_8
XFILLER_33_956 VPWR VGND sg13g2_decap_8
X_3840_ VGND VPWR net769 _0156_ _0157_ _1285_ sg13g2_a21oi_1
X_3771_ _1238_ _0955_ _0969_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_639 VPWR VGND sg13g2_decap_8
X_2722_ net61 sap_3_inst.out\[1\] net766 _0019_ VPWR VGND sg13g2_mux2_1
XFILLER_13_691 VPWR VGND sg13g2_decap_8
XFILLER_9_684 VPWR VGND sg13g2_decap_8
X_2653_ _0237_ _0240_ _0247_ net17 VPWR VGND sg13g2_or3_1
X_2584_ _1993_ _1994_ _1992_ _1995_ VPWR VGND sg13g2_nand3_1
XFILLER_41_1004 VPWR VGND sg13g2_decap_8
X_4185_ net793 VGND VPWR _0163_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[1\]
+ clknet_3_3__leaf_clk sg13g2_dfrbpq_1
X_3205_ _0741_ net588 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] net641
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] VPWR VGND sg13g2_a22oi_1
X_3136_ _0657_ net665 _0672_ VPWR VGND sg13g2_nor2_2
X_3067_ _1582_ _1662_ _0603_ VPWR VGND sg13g2_nor2_1
X_2018_ VPWR _1441_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_23_400 VPWR VGND sg13g2_decap_8
XFILLER_23_411 VPWR VGND sg13g2_fill_2
XFILLER_36_794 VPWR VGND sg13g2_decap_8
XFILLER_11_606 VPWR VGND sg13g2_decap_8
XFILLER_24_967 VPWR VGND sg13g2_decap_8
X_3969_ _1392_ _1393_ _0311_ _1394_ VPWR VGND sg13g2_nand3_1
Xfanout630 _1798_ net630 VPWR VGND sg13g2_buf_8
Xfanout641 net642 net641 VPWR VGND sg13g2_buf_8
Xfanout663 net664 net663 VPWR VGND sg13g2_buf_8
Xfanout674 _0260_ net674 VPWR VGND sg13g2_buf_8
Xfanout685 _1674_ net685 VPWR VGND sg13g2_buf_8
Xfanout652 net654 net652 VPWR VGND sg13g2_buf_8
XFILLER_46_514 VPWR VGND sg13g2_decap_8
Xfanout696 net701 net696 VPWR VGND sg13g2_buf_8
XFILLER_42_720 VPWR VGND sg13g2_decap_8
XFILLER_14_400 VPWR VGND sg13g2_fill_2
XFILLER_15_934 VPWR VGND sg13g2_decap_8
XFILLER_18_1006 VPWR VGND sg13g2_decap_8
XFILLER_42_797 VPWR VGND sg13g2_decap_8
XFILLER_14_488 VPWR VGND sg13g2_decap_8
XFILLER_30_948 VPWR VGND sg13g2_decap_8
XFILLER_6_610 VPWR VGND sg13g2_decap_8
XFILLER_10_650 VPWR VGND sg13g2_decap_8
XFILLER_6_687 VPWR VGND sg13g2_decap_8
XFILLER_5_142 VPWR VGND sg13g2_fill_1
XFILLER_2_882 VPWR VGND sg13g2_decap_8
XFILLER_49_374 VPWR VGND sg13g2_decap_8
XFILLER_18_761 VPWR VGND sg13g2_decap_8
XFILLER_25_709 VPWR VGND sg13g2_decap_8
XFILLER_37_569 VPWR VGND sg13g2_decap_8
XFILLER_33_753 VPWR VGND sg13g2_decap_8
X_3823_ VPWR VGND _0633_ _1109_ _1273_ _0973_ _1274_ _1272_ sg13g2_a221oi_1
XFILLER_21_926 VPWR VGND sg13g2_decap_8
X_3754_ _1045_ VPWR _1225_ VGND net10 net666 sg13g2_o21ai_1
X_2705_ net707 _1628_ _0284_ VPWR VGND sg13g2_nor2_1
X_3685_ net647 net569 _1181_ VPWR VGND sg13g2_nor2b_2
X_2636_ _0229_ _0230_ _0231_ VPWR VGND sg13g2_and2_1
X_2567_ _1978_ sap_3_inst.alu.flags\[2\] _1955_ VPWR VGND sg13g2_nand2b_1
X_2498_ _1911_ _1912_ _1913_ VPWR VGND sg13g2_and2_1
X_4168_ net776 VGND VPWR _0146_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_547 VPWR VGND sg13g2_decap_8
X_3119_ _1502_ _1831_ _0654_ _0655_ VPWR VGND sg13g2_or3_1
X_4099_ net786 VGND VPWR _0077_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_24_764 VPWR VGND sg13g2_decap_8
XFILLER_36_591 VPWR VGND sg13g2_decap_8
XFILLER_12_959 VPWR VGND sg13g2_decap_8
XFILLER_23_33 VPWR VGND sg13g2_fill_1
XFILLER_3_668 VPWR VGND sg13g2_decap_8
XFILLER_47_801 VPWR VGND sg13g2_decap_8
XFILLER_47_878 VPWR VGND sg13g2_decap_8
XFILLER_46_344 VPWR VGND sg13g2_decap_8
XFILLER_19_558 VPWR VGND sg13g2_decap_8
XFILLER_46_388 VPWR VGND sg13g2_decap_8
XFILLER_15_731 VPWR VGND sg13g2_decap_8
XFILLER_42_594 VPWR VGND sg13g2_decap_8
XFILLER_30_745 VPWR VGND sg13g2_decap_8
XFILLER_11_970 VPWR VGND sg13g2_decap_8
XFILLER_7_930 VPWR VGND sg13g2_decap_8
XFILLER_6_484 VPWR VGND sg13g2_decap_8
X_3470_ _0757_ VPWR _1000_ VGND net559 _0854_ sg13g2_o21ai_1
X_2421_ _1835_ _1836_ _1837_ _1839_ _1842_ VPWR VGND sg13g2_nor4_1
X_2352_ VPWR _1773_ _1772_ VGND sg13g2_inv_1
X_2283_ _1704_ _1559_ _1647_ VPWR VGND sg13g2_nand2_1
X_4022_ VGND VPWR _1412_ _0187_ _0195_ _1430_ sg13g2_a21oi_1
XFILLER_38_823 VPWR VGND sg13g2_decap_8
XFILLER_25_506 VPWR VGND sg13g2_decap_8
XFILLER_21_723 VPWR VGND sg13g2_decap_8
XFILLER_33_550 VPWR VGND sg13g2_decap_8
X_3806_ net10 _1086_ _1261_ VPWR VGND sg13g2_nor2_1
X_3737_ _0125_ _1214_ _1049_ net556 _1449_ VPWR VGND sg13g2_a22oi_1
X_3668_ _1161_ VPWR _0104_ VGND _1165_ _1166_ sg13g2_o21ai_1
X_3599_ _1104_ VPWR _0088_ VGND _1111_ _1113_ sg13g2_o21ai_1
X_2619_ _0216_ net620 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] net637
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_0_638 VPWR VGND sg13g2_decap_8
XFILLER_44_815 VPWR VGND sg13g2_decap_8
XFILLER_29_867 VPWR VGND sg13g2_decap_8
XFILLER_24_561 VPWR VGND sg13g2_decap_8
XFILLER_12_756 VPWR VGND sg13g2_decap_8
XFILLER_8_727 VPWR VGND sg13g2_decap_8
XFILLER_4_922 VPWR VGND sg13g2_decap_8
XFILLER_4_999 VPWR VGND sg13g2_decap_8
XFILLER_3_465 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_47_675 VPWR VGND sg13g2_decap_8
XFILLER_34_347 VPWR VGND sg13g2_fill_1
X_2970_ net554 net745 _0532_ _0040_ VPWR VGND sg13g2_a21o_1
XFILLER_30_542 VPWR VGND sg13g2_decap_8
X_3522_ VGND VPWR _0822_ _0907_ _1048_ net583 sg13g2_a21oi_1
X_3453_ _0984_ net578 _0983_ VPWR VGND sg13g2_nand2_1
X_2404_ VGND VPWR net683 _1820_ _1825_ _1824_ sg13g2_a21oi_1
X_3384_ VPWR _0917_ _0916_ VGND sg13g2_inv_1
X_2335_ _1583_ net681 net723 _1756_ VPWR VGND _1646_ sg13g2_nand4_1
X_2266_ net714 _1634_ _1687_ VPWR VGND sg13g2_nor2_1
XFILLER_38_620 VPWR VGND sg13g2_decap_8
X_2197_ _1586_ net680 _1618_ VPWR VGND sg13g2_nor2b_1
X_4005_ u_ser.shadow_reg\[0\] VPWR _1421_ VGND u_ser.state\[0\] _1433_ sg13g2_o21ai_1
XFILLER_37_174 VPWR VGND sg13g2_fill_1
XFILLER_38_697 VPWR VGND sg13g2_decap_8
XFILLER_41_829 VPWR VGND sg13g2_decap_8
XFILLER_13_509 VPWR VGND sg13g2_decap_8
XFILLER_21_520 VPWR VGND sg13g2_decap_8
XFILLER_14_1020 VPWR VGND sg13g2_decap_8
XFILLER_21_597 VPWR VGND sg13g2_decap_8
XFILLER_5_719 VPWR VGND sg13g2_decap_8
XFILLER_0_435 VPWR VGND sg13g2_decap_8
XFILLER_1_947 VPWR VGND sg13g2_decap_8
Xhold32 sap_3_inst.reg_file.array_serializer_inst.word_index\[2\] VPWR VGND net79
+ sg13g2_dlygate4sd3_1
Xhold10 u_ser.shadow_reg\[3\] VPWR VGND net57 sg13g2_dlygate4sd3_1
Xhold21 sap_3_outputReg_start_sync VPWR VGND net68 sg13g2_dlygate4sd3_1
XFILLER_21_1024 VPWR VGND sg13g2_decap_4
XFILLER_29_664 VPWR VGND sg13g2_decap_8
XFILLER_44_612 VPWR VGND sg13g2_decap_8
XFILLER_17_815 VPWR VGND sg13g2_decap_8
XFILLER_16_336 VPWR VGND sg13g2_fill_1
XFILLER_16_358 VPWR VGND sg13g2_fill_2
XFILLER_44_689 VPWR VGND sg13g2_decap_8
XFILLER_25_870 VPWR VGND sg13g2_decap_8
XFILLER_40_851 VPWR VGND sg13g2_decap_8
XFILLER_12_553 VPWR VGND sg13g2_decap_8
XFILLER_8_524 VPWR VGND sg13g2_decap_8
XFILLER_6_36 VPWR VGND sg13g2_decap_4
XFILLER_4_796 VPWR VGND sg13g2_decap_8
X_2120_ _1540_ net698 net712 _1541_ VPWR VGND sg13g2_a21o_1
XFILLER_48_962 VPWR VGND sg13g2_decap_8
X_2051_ VPWR _1474_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_47_472 VPWR VGND sg13g2_decap_8
XFILLER_19_174 VPWR VGND sg13g2_fill_2
XFILLER_23_829 VPWR VGND sg13g2_decap_8
XFILLER_35_667 VPWR VGND sg13g2_decap_8
X_2953_ _0515_ _0507_ _0516_ VPWR VGND sg13g2_xor2_1
XFILLER_22_328 VPWR VGND sg13g2_fill_1
XFILLER_31_862 VPWR VGND sg13g2_decap_8
X_2884_ _0447_ _0448_ _0449_ VPWR VGND sg13g2_and2_1
XFILLER_30_372 VPWR VGND sg13g2_fill_2
X_3505_ net578 _1031_ _1033_ _1034_ VPWR VGND sg13g2_nor3_1
X_3436_ _0965_ _0966_ _0967_ VPWR VGND _0964_ sg13g2_nand3b_1
X_3367_ _0901_ _0900_ net584 _0898_ net577 VPWR VGND sg13g2_a22oi_1
X_2318_ net683 VPWR _1739_ VGND _1509_ _1545_ sg13g2_o21ai_1
Xheichips25_template_34 VPWR VGND uo_out[7] sg13g2_tielo
X_3298_ _0674_ VPWR _0834_ VGND _0683_ _0833_ sg13g2_o21ai_1
X_2249_ VGND VPWR _1569_ _1669_ _1670_ _1572_ sg13g2_a21oi_1
XFILLER_38_494 VPWR VGND sg13g2_decap_8
XFILLER_26_667 VPWR VGND sg13g2_decap_8
XFILLER_41_626 VPWR VGND sg13g2_decap_8
XFILLER_25_177 VPWR VGND sg13g2_fill_2
XFILLER_22_862 VPWR VGND sg13g2_decap_8
XFILLER_5_516 VPWR VGND sg13g2_decap_8
Xoutput22 net22 uio_out[5] VPWR VGND sg13g2_buf_1
Xoutput9 net9 uio_oe[0] VPWR VGND sg13g2_buf_1
Xoutput11 net11 uio_oe[2] VPWR VGND sg13g2_buf_1
XFILLER_1_744 VPWR VGND sg13g2_decap_8
XFILLER_49_759 VPWR VGND sg13g2_decap_8
XFILLER_17_612 VPWR VGND sg13g2_decap_8
XFILLER_29_461 VPWR VGND sg13g2_decap_8
XFILLER_45_954 VPWR VGND sg13g2_decap_8
XFILLER_17_689 VPWR VGND sg13g2_decap_8
XFILLER_44_486 VPWR VGND sg13g2_decap_8
XFILLER_31_125 VPWR VGND sg13g2_fill_1
XFILLER_32_637 VPWR VGND sg13g2_decap_8
XFILLER_13_873 VPWR VGND sg13g2_decap_8
XFILLER_31_169 VPWR VGND sg13g2_fill_1
XFILLER_9_866 VPWR VGND sg13g2_decap_8
XFILLER_4_593 VPWR VGND sg13g2_decap_8
X_3221_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] _0756_
+ net609 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] _0757_ net615 sg13g2_a221oi_1
X_3152_ VPWR VGND _1589_ _0687_ _1932_ _1615_ _0688_ _1704_ sg13g2_a221oi_1
X_2103_ net738 net725 net727 _1524_ VPWR VGND sg13g2_or3_1
X_3083_ _0614_ _0615_ _0612_ _0619_ VPWR VGND sg13g2_nand3_1
X_2034_ _1457_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[1\] VPWR VGND
+ sg13g2_inv_2
XFILLER_36_976 VPWR VGND sg13g2_decap_8
XFILLER_23_626 VPWR VGND sg13g2_decap_8
X_3985_ _0510_ net663 _1404_ VPWR VGND sg13g2_nor2_1
XFILLER_22_158 VPWR VGND sg13g2_fill_1
X_2936_ _0499_ net747 net555 _0039_ VPWR VGND sg13g2_mux2_1
X_2867_ _0433_ _0392_ _0431_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_1012 VPWR VGND sg13g2_decap_8
X_2798_ _0321_ _0355_ net720 _0366_ VPWR VGND sg13g2_nand3_1
Xclkbuf_1_0__f_clk_div_out clknet_0_clk_div_out clknet_1_0__leaf_clk_div_out VPWR
+ VGND sg13g2_buf_8
Xfanout801 rst_n net801 VPWR VGND sg13g2_buf_8
X_3419_ VGND VPWR _0788_ _0849_ _0951_ _0776_ sg13g2_a21oi_1
XFILLER_27_921 VPWR VGND sg13g2_decap_8
XFILLER_42_902 VPWR VGND sg13g2_decap_8
XFILLER_26_464 VPWR VGND sg13g2_decap_8
XFILLER_27_998 VPWR VGND sg13g2_decap_8
XFILLER_42_979 VPWR VGND sg13g2_decap_8
XFILLER_42_87 VPWR VGND sg13g2_fill_1
XFILLER_10_832 VPWR VGND sg13g2_decap_8
XFILLER_42_98 VPWR VGND sg13g2_fill_1
XFILLER_6_869 VPWR VGND sg13g2_decap_8
XFILLER_1_541 VPWR VGND sg13g2_decap_8
XFILLER_49_556 VPWR VGND sg13g2_decap_8
XFILLER_18_943 VPWR VGND sg13g2_decap_8
XFILLER_45_751 VPWR VGND sg13g2_decap_8
XFILLER_33_935 VPWR VGND sg13g2_decap_8
X_3770_ _0135_ _1102_ _1237_ net598 _1471_ VPWR VGND sg13g2_a22oi_1
XFILLER_13_670 VPWR VGND sg13g2_decap_8
XFILLER_20_618 VPWR VGND sg13g2_decap_8
XFILLER_34_1012 VPWR VGND sg13g2_decap_8
XFILLER_41_990 VPWR VGND sg13g2_decap_8
X_2721_ net70 sap_3_inst.out\[0\] net766 _0018_ VPWR VGND sg13g2_mux2_1
XFILLER_9_663 VPWR VGND sg13g2_decap_8
X_2652_ VGND VPWR _0243_ _0246_ _0247_ net566 sg13g2_a21oi_1
X_2583_ _1994_ net620 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] net632
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_880 VPWR VGND sg13g2_decap_8
X_3204_ _0713_ _0731_ _0740_ VPWR VGND sg13g2_nor2_2
X_4184_ net794 VGND VPWR _0162_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[0\]
+ clknet_3_6__leaf_clk sg13g2_dfrbpq_1
X_3135_ _0671_ _0660_ _0669_ VPWR VGND sg13g2_nand2_1
XFILLER_28_729 VPWR VGND sg13g2_decap_8
X_3066_ VPWR VGND _1716_ net689 _1839_ net723 _0602_ _1838_ sg13g2_a221oi_1
X_2017_ _1440_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[3\] VPWR VGND
+ sg13g2_inv_2
XFILLER_36_773 VPWR VGND sg13g2_decap_8
XFILLER_24_946 VPWR VGND sg13g2_decap_8
XFILLER_23_445 VPWR VGND sg13g2_decap_8
X_3968_ _1393_ _1938_ _0315_ VPWR VGND sg13g2_nand2_1
X_2919_ _0483_ _0482_ _2008_ _0478_ net563 VPWR VGND sg13g2_a22oi_1
X_3899_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] _1308_
+ _1338_ net762 sg13g2_a21oi_1
Xfanout642 _0737_ net642 VPWR VGND sg13g2_buf_8
Xfanout620 _1803_ net620 VPWR VGND sg13g2_buf_8
Xfanout631 net632 net631 VPWR VGND sg13g2_buf_8
Xfanout664 _1391_ net664 VPWR VGND sg13g2_buf_8
Xfanout675 _1857_ net675 VPWR VGND sg13g2_buf_8
Xfanout653 net654 net653 VPWR VGND sg13g2_buf_8
Xfanout686 _1582_ net686 VPWR VGND sg13g2_buf_8
Xfanout697 net701 net697 VPWR VGND sg13g2_buf_1
XFILLER_18_228 VPWR VGND sg13g2_fill_1
XFILLER_15_913 VPWR VGND sg13g2_decap_8
XFILLER_33_209 VPWR VGND sg13g2_fill_2
XFILLER_14_423 VPWR VGND sg13g2_fill_1
XFILLER_26_272 VPWR VGND sg13g2_fill_2
XFILLER_27_795 VPWR VGND sg13g2_decap_8
XFILLER_42_776 VPWR VGND sg13g2_decap_8
XFILLER_41_253 VPWR VGND sg13g2_fill_1
XFILLER_30_927 VPWR VGND sg13g2_decap_8
XFILLER_23_990 VPWR VGND sg13g2_decap_8
XFILLER_6_666 VPWR VGND sg13g2_decap_8
XFILLER_2_861 VPWR VGND sg13g2_decap_8
XFILLER_49_353 VPWR VGND sg13g2_decap_8
XFILLER_37_548 VPWR VGND sg13g2_decap_8
XFILLER_18_740 VPWR VGND sg13g2_decap_8
XFILLER_21_905 VPWR VGND sg13g2_decap_8
XFILLER_33_732 VPWR VGND sg13g2_decap_8
X_3822_ net14 net661 net602 _1273_ VPWR VGND sg13g2_or3_1
X_3753_ _0873_ _1223_ _0844_ _1224_ VPWR VGND sg13g2_nand3_1
X_3684_ _0106_ _1179_ _1180_ net597 _1495_ VPWR VGND sg13g2_a22oi_1
X_2704_ _1514_ net699 _1508_ _0001_ VPWR VGND sg13g2_nand3_1
X_2635_ _0230_ net624 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] net635
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2566_ sap_3_inst.alu.flags\[3\] _1977_ _1955_ _0029_ VPWR VGND sg13g2_mux2_1
X_2497_ _1912_ net625 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] net633
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4167_ net780 VGND VPWR _0145_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\]
+ clknet_5_13__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3118_ VGND VPWR net731 _1716_ _0654_ net702 sg13g2_a21oi_1
XFILLER_28_526 VPWR VGND sg13g2_decap_8
X_4098_ net786 VGND VPWR _0076_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\]
+ clknet_5_25__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3049_ _0591_ VPWR _0060_ VGND net693 _0225_ sg13g2_o21ai_1
XFILLER_15_209 VPWR VGND sg13g2_fill_1
XFILLER_36_570 VPWR VGND sg13g2_decap_8
XFILLER_24_743 VPWR VGND sg13g2_decap_8
XFILLER_12_938 VPWR VGND sg13g2_decap_8
XFILLER_8_909 VPWR VGND sg13g2_decap_8
XFILLER_20_982 VPWR VGND sg13g2_decap_8
XFILLER_3_647 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_135 VPWR VGND sg13g2_fill_1
XFILLER_47_857 VPWR VGND sg13g2_decap_8
XFILLER_46_301 VPWR VGND sg13g2_fill_2
XFILLER_19_537 VPWR VGND sg13g2_decap_8
XFILLER_46_367 VPWR VGND sg13g2_decap_8
XFILLER_15_710 VPWR VGND sg13g2_decap_8
XFILLER_34_529 VPWR VGND sg13g2_decap_8
XFILLER_14_220 VPWR VGND sg13g2_fill_2
XFILLER_27_592 VPWR VGND sg13g2_decap_8
XFILLER_42_573 VPWR VGND sg13g2_decap_8
XFILLER_15_787 VPWR VGND sg13g2_decap_8
XFILLER_30_724 VPWR VGND sg13g2_decap_8
XFILLER_7_986 VPWR VGND sg13g2_decap_8
X_2420_ _1833_ VPWR _1841_ VGND _1602_ _1840_ sg13g2_o21ai_1
XFILLER_9_1027 VPWR VGND sg13g2_fill_2
X_2351_ _1570_ _1771_ _1503_ _1772_ VPWR VGND sg13g2_nand3_1
X_2282_ _1703_ net704 net714 net710 net711 VPWR VGND sg13g2_a22oi_1
X_4021_ VGND VPWR net767 _0187_ _1430_ net71 sg13g2_a21oi_1
XFILLER_38_802 VPWR VGND sg13g2_decap_8
XFILLER_38_879 VPWR VGND sg13g2_decap_8
XFILLER_21_702 VPWR VGND sg13g2_decap_8
XFILLER_21_779 VPWR VGND sg13g2_decap_8
X_3805_ net604 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] _1260_ _0147_
+ VPWR VGND sg13g2_a21o_1
XFILLER_20_267 VPWR VGND sg13g2_fill_1
X_3736_ _1050_ net556 _1214_ VPWR VGND sg13g2_nor2_1
X_3667_ _1166_ net651 _1112_ VPWR VGND sg13g2_nand2_1
XFILLER_47_1011 VPWR VGND sg13g2_decap_8
X_3598_ _1113_ net592 _1112_ VPWR VGND sg13g2_nand2_1
X_2618_ _0215_ net2 _1847_ VPWR VGND sg13g2_nand2_1
XFILLER_0_617 VPWR VGND sg13g2_decap_8
X_2549_ _1962_ _1959_ _1960_ _1961_ VPWR VGND sg13g2_and3_1
X_4219_ net784 VGND VPWR net59 u_ser.bit_pos\[2\] clknet_3_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_29_846 VPWR VGND sg13g2_decap_8
XFILLER_16_529 VPWR VGND sg13g2_decap_8
XFILLER_24_540 VPWR VGND sg13g2_decap_8
XFILLER_12_735 VPWR VGND sg13g2_decap_8
XFILLER_8_706 VPWR VGND sg13g2_decap_8
XFILLER_7_227 VPWR VGND sg13g2_fill_2
XFILLER_4_901 VPWR VGND sg13g2_decap_8
XFILLER_3_400 VPWR VGND sg13g2_fill_2
XFILLER_4_978 VPWR VGND sg13g2_decap_8
XFILLER_3_444 VPWR VGND sg13g2_decap_8
XFILLER_47_654 VPWR VGND sg13g2_decap_8
XFILLER_46_120 VPWR VGND sg13g2_fill_2
XFILLER_35_849 VPWR VGND sg13g2_decap_8
XFILLER_28_890 VPWR VGND sg13g2_decap_8
XFILLER_15_584 VPWR VGND sg13g2_decap_8
XFILLER_30_521 VPWR VGND sg13g2_decap_8
XFILLER_30_598 VPWR VGND sg13g2_decap_8
X_3521_ _1047_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] net557 _0076_
+ VPWR VGND sg13g2_mux2_1
XFILLER_7_783 VPWR VGND sg13g2_decap_8
X_3452_ _0983_ _0956_ _0970_ VPWR VGND sg13g2_xnor2_1
X_2403_ VGND VPWR _1510_ _1821_ _1824_ _1823_ sg13g2_a21oi_1
X_3383_ _0915_ VPWR _0916_ VGND _0910_ _0914_ sg13g2_o21ai_1
X_2334_ net699 _1565_ net742 _1755_ VPWR VGND _1754_ sg13g2_nand4_1
X_2265_ net733 _1616_ _1642_ _1686_ VPWR VGND sg13g2_or3_1
X_4004_ _1410_ _1419_ _1434_ _1420_ VPWR VGND sg13g2_nand3_1
X_2196_ _1594_ _1601_ _1608_ _1613_ _1617_ VPWR VGND sg13g2_nor4_1
XFILLER_37_142 VPWR VGND sg13g2_fill_2
XFILLER_38_676 VPWR VGND sg13g2_decap_8
XFILLER_26_849 VPWR VGND sg13g2_decap_8
XFILLER_37_186 VPWR VGND sg13g2_fill_2
XFILLER_41_808 VPWR VGND sg13g2_decap_8
XFILLER_34_893 VPWR VGND sg13g2_decap_8
XFILLER_21_576 VPWR VGND sg13g2_decap_8
X_3719_ _1204_ _0921_ _1203_ net595 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_0_403 VPWR VGND sg13g2_fill_1
XFILLER_1_926 VPWR VGND sg13g2_decap_8
Xhold22 _0189_ VPWR VGND net69 sg13g2_dlygate4sd3_1
Xhold11 u_ser.state\[0\] VPWR VGND net58 sg13g2_dlygate4sd3_1
Xhold33 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[0\] VPWR VGND net80 sg13g2_dlygate4sd3_1
XFILLER_21_1003 VPWR VGND sg13g2_decap_8
XFILLER_29_643 VPWR VGND sg13g2_decap_8
XFILLER_28_164 VPWR VGND sg13g2_fill_1
XFILLER_44_668 VPWR VGND sg13g2_decap_8
XFILLER_32_819 VPWR VGND sg13g2_decap_8
XFILLER_40_830 VPWR VGND sg13g2_decap_8
XFILLER_8_503 VPWR VGND sg13g2_decap_8
XFILLER_12_532 VPWR VGND sg13g2_decap_8
XFILLER_4_775 VPWR VGND sg13g2_decap_8
XFILLER_0_981 VPWR VGND sg13g2_decap_8
XFILLER_48_941 VPWR VGND sg13g2_decap_8
X_2050_ VPWR _1473_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_47_451 VPWR VGND sg13g2_decap_8
XFILLER_35_646 VPWR VGND sg13g2_decap_8
Xclkbuf_5_21__f_sap_3_inst.alu.clk_regs clknet_4_10_0_sap_3_inst.alu.clk_regs clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_23_808 VPWR VGND sg13g2_decap_8
XFILLER_37_1010 VPWR VGND sg13g2_decap_8
X_2952_ _0478_ VPWR _0515_ VGND _0449_ _0514_ sg13g2_o21ai_1
XFILLER_16_893 VPWR VGND sg13g2_decap_8
XFILLER_31_841 VPWR VGND sg13g2_decap_8
X_2883_ VGND VPWR _0416_ _0424_ _0448_ _0417_ sg13g2_a21oi_1
X_3504_ net574 _1032_ _1033_ VPWR VGND sg13g2_nor2_1
XFILLER_7_580 VPWR VGND sg13g2_decap_8
X_3435_ _0966_ net592 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] net640
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_44_1025 VPWR VGND sg13g2_decap_4
X_3366_ _0900_ _0882_ _0894_ VPWR VGND sg13g2_xnor2_1
X_3297_ _0686_ _0832_ _0612_ _0833_ VPWR VGND sg13g2_nand3_1
X_2317_ _1736_ _1737_ _1699_ _1738_ VPWR VGND sg13g2_nand3_1
X_2248_ _1619_ VPWR _1669_ VGND _1632_ _1668_ sg13g2_o21ai_1
XFILLER_39_985 VPWR VGND sg13g2_decap_8
X_2179_ VPWR _1600_ _1599_ VGND sg13g2_inv_1
XFILLER_26_646 VPWR VGND sg13g2_decap_8
XFILLER_41_605 VPWR VGND sg13g2_decap_8
XFILLER_25_145 VPWR VGND sg13g2_fill_1
XFILLER_15_57 VPWR VGND sg13g2_fill_2
XFILLER_22_841 VPWR VGND sg13g2_decap_8
XFILLER_34_690 VPWR VGND sg13g2_decap_8
XFILLER_40_148 VPWR VGND sg13g2_fill_1
Xoutput23 net23 uio_out[6] VPWR VGND sg13g2_buf_1
Xoutput12 net12 uio_oe[3] VPWR VGND sg13g2_buf_1
XFILLER_1_723 VPWR VGND sg13g2_decap_8
XFILLER_49_738 VPWR VGND sg13g2_decap_8
XFILLER_45_933 VPWR VGND sg13g2_decap_8
XFILLER_44_465 VPWR VGND sg13g2_decap_8
XFILLER_17_668 VPWR VGND sg13g2_decap_8
XFILLER_31_115 VPWR VGND sg13g2_fill_1
XFILLER_32_616 VPWR VGND sg13g2_decap_8
XFILLER_13_852 VPWR VGND sg13g2_decap_8
XFILLER_9_845 VPWR VGND sg13g2_decap_8
XFILLER_4_572 VPWR VGND sg13g2_decap_8
XFILLER_28_1009 VPWR VGND sg13g2_decap_8
X_3220_ _0753_ _0754_ _0752_ _0756_ VPWR VGND _0755_ sg13g2_nand4_1
X_3151_ _1438_ _1590_ _0638_ _0687_ VPWR VGND sg13g2_nor3_2
X_2102_ net738 net725 net727 _1523_ VPWR VGND sg13g2_nor3_1
XFILLER_39_226 VPWR VGND sg13g2_fill_1
X_3082_ _1596_ _1599_ net707 _1661_ _0618_ VPWR VGND sg13g2_nor4_1
X_2033_ VPWR _1456_ net760 VGND sg13g2_inv_1
XFILLER_36_955 VPWR VGND sg13g2_decap_8
XFILLER_23_605 VPWR VGND sg13g2_decap_8
X_3984_ _1403_ sap_3_inst.alu.act\[5\] net548 _0183_ VPWR VGND sg13g2_mux2_1
XFILLER_16_690 VPWR VGND sg13g2_decap_8
X_2935_ VGND VPWR _1899_ net616 _0499_ _0498_ sg13g2_a21oi_1
X_2866_ _0432_ _0431_ VPWR VGND _0392_ sg13g2_nand2b_2
X_2797_ VPWR VGND _0333_ _0364_ _0355_ net759 _0365_ net573 sg13g2_a221oi_1
XFILLER_7_91 VPWR VGND sg13g2_fill_2
X_3418_ _0950_ _0838_ net13 VPWR VGND sg13g2_nand2b_1
X_3349_ _0884_ net584 _0883_ VPWR VGND sg13g2_nand2_2
XFILLER_27_900 VPWR VGND sg13g2_decap_8
XFILLER_39_782 VPWR VGND sg13g2_decap_8
XFILLER_26_443 VPWR VGND sg13g2_decap_8
XFILLER_27_977 VPWR VGND sg13g2_decap_8
XFILLER_42_958 VPWR VGND sg13g2_decap_8
XFILLER_14_649 VPWR VGND sg13g2_decap_8
XFILLER_41_479 VPWR VGND sg13g2_decap_8
XFILLER_10_811 VPWR VGND sg13g2_decap_8
XFILLER_10_888 VPWR VGND sg13g2_decap_8
XFILLER_6_848 VPWR VGND sg13g2_decap_8
XFILLER_1_520 VPWR VGND sg13g2_decap_8
XFILLER_49_535 VPWR VGND sg13g2_decap_8
XFILLER_1_597 VPWR VGND sg13g2_decap_8
XFILLER_45_730 VPWR VGND sg13g2_decap_8
XFILLER_18_922 VPWR VGND sg13g2_decap_8
XFILLER_33_914 VPWR VGND sg13g2_decap_8
XFILLER_18_999 VPWR VGND sg13g2_decap_8
X_2720_ u_ser.state\[0\] u_ser.state\[1\] _0186_ VPWR VGND sg13g2_nor2_2
XFILLER_9_642 VPWR VGND sg13g2_decap_8
X_2651_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] _0245_
+ net619 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] _0246_ net623 sg13g2_a221oi_1
X_2582_ _1993_ net628 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] net636
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] VPWR VGND sg13g2_a22oi_1
X_3203_ _0739_ net659 _0719_ VPWR VGND sg13g2_nand2_1
X_4183_ net799 VGND VPWR net67 regFile_serial clknet_3_6__leaf_clk sg13g2_dfrbpq_1
X_3134_ _0660_ _0669_ _0670_ VPWR VGND sg13g2_and2_1
XFILLER_28_708 VPWR VGND sg13g2_decap_8
X_3065_ _1594_ VPWR _0601_ VGND _1581_ _1646_ sg13g2_o21ai_1
X_2016_ VPWR _1439_ net725 VGND sg13g2_inv_1
XFILLER_36_752 VPWR VGND sg13g2_decap_8
XFILLER_24_925 VPWR VGND sg13g2_decap_8
Xclkbuf_5_18__f_sap_3_inst.alu.clk_regs clknet_4_9_0_sap_3_inst.alu.clk_regs clknet_5_18__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_23_424 VPWR VGND sg13g2_decap_8
X_3967_ _1392_ net617 net664 VPWR VGND sg13g2_nand2b_1
XFILLER_23_479 VPWR VGND sg13g2_decap_8
X_2918_ _0432_ _0447_ _0479_ _0482_ VPWR VGND sg13g2_nor3_1
XFILLER_32_980 VPWR VGND sg13g2_decap_8
X_3898_ _1337_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] _1311_
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2849_ net753 sap_3_inst.alu.tmp\[3\] _0415_ VPWR VGND sg13g2_and2_1
XFILLER_3_829 VPWR VGND sg13g2_decap_8
Xfanout610 _0715_ net610 VPWR VGND sg13g2_buf_8
Xfanout632 _1797_ net632 VPWR VGND sg13g2_buf_8
Xfanout621 net622 net621 VPWR VGND sg13g2_buf_8
Xfanout643 net645 net643 VPWR VGND sg13g2_buf_8
Xfanout676 _1857_ net676 VPWR VGND sg13g2_buf_1
Xfanout665 _0671_ net665 VPWR VGND sg13g2_buf_8
Xfanout654 _0726_ net654 VPWR VGND sg13g2_buf_8
Xfanout687 net688 net687 VPWR VGND sg13g2_buf_8
Xfanout698 net701 net698 VPWR VGND sg13g2_buf_8
XFILLER_19_719 VPWR VGND sg13g2_decap_8
XFILLER_46_549 VPWR VGND sg13g2_decap_8
XFILLER_2_1022 VPWR VGND sg13g2_decap_8
XFILLER_27_774 VPWR VGND sg13g2_decap_8
XFILLER_42_755 VPWR VGND sg13g2_decap_8
XFILLER_15_969 VPWR VGND sg13g2_decap_8
XFILLER_30_906 VPWR VGND sg13g2_decap_8
XFILLER_6_645 VPWR VGND sg13g2_decap_8
XFILLER_10_685 VPWR VGND sg13g2_decap_8
XFILLER_2_840 VPWR VGND sg13g2_decap_8
XFILLER_49_332 VPWR VGND sg13g2_decap_8
XFILLER_37_527 VPWR VGND sg13g2_decap_8
XFILLER_18_796 VPWR VGND sg13g2_decap_8
XFILLER_33_711 VPWR VGND sg13g2_decap_8
X_3821_ VGND VPWR net602 _0975_ _1272_ net583 sg13g2_a21oi_1
XFILLER_33_788 VPWR VGND sg13g2_decap_8
X_3752_ _1223_ _0871_ _0857_ VPWR VGND sg13g2_nand2b_1
X_3683_ net651 _1125_ _1180_ VPWR VGND sg13g2_and2_1
X_2703_ net565 _1810_ net16 VPWR VGND sg13g2_nor2b_2
X_2634_ _0229_ net629 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] net633
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2565_ VGND VPWR net675 _1975_ _1977_ _1976_ sg13g2_a21oi_1
X_2496_ _1911_ net623 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] net635
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_4_81 VPWR VGND sg13g2_fill_1
X_4166_ net776 VGND VPWR _0144_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_505 VPWR VGND sg13g2_decap_8
X_3117_ _0653_ net702 _0652_ VPWR VGND sg13g2_nand2_1
X_4097_ net797 VGND VPWR _0075_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\]
+ clknet_5_29__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3048_ _0591_ sap_3_inst.controller.opcode\[1\] net693 VPWR VGND sg13g2_nand2_1
XFILLER_24_722 VPWR VGND sg13g2_decap_8
XFILLER_12_917 VPWR VGND sg13g2_decap_8
XFILLER_24_799 VPWR VGND sg13g2_decap_8
XFILLER_20_961 VPWR VGND sg13g2_decap_8
XFILLER_3_626 VPWR VGND sg13g2_decap_8
XFILLER_2_147 VPWR VGND sg13g2_decap_4
XFILLER_24_1023 VPWR VGND sg13g2_decap_4
XFILLER_47_836 VPWR VGND sg13g2_decap_8
XFILLER_19_516 VPWR VGND sg13g2_decap_8
XFILLER_34_508 VPWR VGND sg13g2_decap_8
XFILLER_27_571 VPWR VGND sg13g2_decap_8
XFILLER_42_552 VPWR VGND sg13g2_decap_8
XFILLER_15_766 VPWR VGND sg13g2_decap_8
XFILLER_30_703 VPWR VGND sg13g2_decap_8
XFILLER_31_1016 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_7_965 VPWR VGND sg13g2_decap_8
Xsap_3_inst.clock.clock_gate_inst _0001_ clknet_1_1__leaf_clk_div_out sap_3_inst.alu.clk
+ VPWR VGND sg13g2_lgcp_1
X_2350_ _1619_ VPWR _1771_ VGND _1763_ _1770_ sg13g2_o21ai_1
XFILLER_9_1006 VPWR VGND sg13g2_decap_8
X_2281_ net689 _1664_ _1700_ _1701_ _1702_ VPWR VGND sg13g2_nor4_1
X_4020_ VGND VPWR net767 _0187_ _0194_ _1429_ sg13g2_a21oi_1
XFILLER_38_858 VPWR VGND sg13g2_decap_8
XFILLER_18_593 VPWR VGND sg13g2_decap_8
XFILLER_33_585 VPWR VGND sg13g2_decap_8
XFILLER_21_758 VPWR VGND sg13g2_decap_8
X_3804_ net605 _0861_ _1259_ _1260_ VPWR VGND sg13g2_nor3_1
X_3735_ net556 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] _1213_ _0124_
+ VPWR VGND sg13g2_a21o_1
X_3666_ _1110_ _1162_ _1164_ _1165_ VPWR VGND sg13g2_nor3_1
X_3597_ _1112_ net579 VPWR VGND _0983_ sg13g2_nand2b_2
X_2617_ _0214_ _1828_ net720 _1827_ net757 VPWR VGND sg13g2_a22oi_1
X_2548_ _1961_ net626 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] net628
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2479_ _1896_ _1893_ _1894_ _1895_ VPWR VGND sg13g2_and3_1
X_4218_ net784 VGND VPWR _0195_ u_ser.bit_pos\[1\] clknet_3_2__leaf_clk sg13g2_dfrbpq_2
XFILLER_29_825 VPWR VGND sg13g2_decap_8
X_4149_ net779 VGND VPWR _0127_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\]
+ clknet_5_15__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4028__6 VPWR net40 clknet_leaf_0_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_16_508 VPWR VGND sg13g2_decap_8
XFILLER_37_891 VPWR VGND sg13g2_decap_8
XFILLER_12_714 VPWR VGND sg13g2_decap_8
XFILLER_24_596 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_3_0__leaf_clk clkload0/X VPWR VGND sg13g2_buf_1
XFILLER_4_957 VPWR VGND sg13g2_decap_8
XFILLER_47_633 VPWR VGND sg13g2_decap_8
XFILLER_46_154 VPWR VGND sg13g2_fill_2
XFILLER_34_305 VPWR VGND sg13g2_fill_1
XFILLER_35_828 VPWR VGND sg13g2_decap_8
XFILLER_15_563 VPWR VGND sg13g2_decap_8
XFILLER_43_894 VPWR VGND sg13g2_decap_8
XFILLER_30_500 VPWR VGND sg13g2_decap_8
XFILLER_30_577 VPWR VGND sg13g2_decap_8
X_3520_ _0876_ net580 _1046_ _1047_ VPWR VGND sg13g2_a21o_2
XFILLER_10_290 VPWR VGND sg13g2_fill_1
XFILLER_7_762 VPWR VGND sg13g2_decap_8
X_3451_ net559 _0918_ net552 _0970_ _0982_ VPWR VGND sg13g2_or4_1
X_2402_ _1823_ _1715_ _1822_ VPWR VGND sg13g2_nand2_1
X_3382_ _0915_ _1440_ net615 VPWR VGND sg13g2_nand2_1
XFILLER_3_990 VPWR VGND sg13g2_decap_8
X_2333_ _1754_ _1511_ _1569_ VPWR VGND sg13g2_nand2_1
X_2264_ VGND VPWR _1685_ _1651_ _1616_ sg13g2_or2_1
X_2195_ _1523_ _1614_ _1506_ _1616_ VPWR VGND sg13g2_nand3_1
X_4003_ net767 u_ser.shadow_reg\[1\] u_ser.shadow_reg\[2\] u_ser.shadow_reg\[3\] u_ser.shadow_reg\[4\]
+ u_ser.bit_pos\[1\] _1419_ VPWR VGND sg13g2_mux4_1
XFILLER_38_655 VPWR VGND sg13g2_decap_8
XFILLER_25_316 VPWR VGND sg13g2_fill_2
XFILLER_26_828 VPWR VGND sg13g2_decap_8
XFILLER_1_93 VPWR VGND sg13g2_decap_4
XFILLER_19_880 VPWR VGND sg13g2_decap_8
XFILLER_34_872 VPWR VGND sg13g2_decap_8
XFILLER_21_555 VPWR VGND sg13g2_decap_8
X_3718_ VGND VPWR _1975_ _1053_ _1203_ net595 sg13g2_a21oi_1
X_3649_ _1150_ net546 net568 VPWR VGND sg13g2_nand2_1
XFILLER_1_905 VPWR VGND sg13g2_decap_8
Xhold23 u_ser.shadow_reg\[0\] VPWR VGND net70 sg13g2_dlygate4sd3_1
Xhold12 _0196_ VPWR VGND net59 sg13g2_dlygate4sd3_1
XFILLER_29_622 VPWR VGND sg13g2_decap_8
Xhold34 _0157_ VPWR VGND net81 sg13g2_dlygate4sd3_1
XFILLER_44_647 VPWR VGND sg13g2_decap_8
XFILLER_29_699 VPWR VGND sg13g2_decap_8
XFILLER_45_66 VPWR VGND sg13g2_fill_2
XFILLER_12_511 VPWR VGND sg13g2_decap_8
XFILLER_24_393 VPWR VGND sg13g2_decap_8
XFILLER_40_886 VPWR VGND sg13g2_decap_8
XFILLER_12_588 VPWR VGND sg13g2_decap_8
XFILLER_8_559 VPWR VGND sg13g2_decap_8
XFILLER_6_27 VPWR VGND sg13g2_fill_2
XFILLER_4_754 VPWR VGND sg13g2_decap_8
XFILLER_6_1009 VPWR VGND sg13g2_decap_8
XFILLER_48_920 VPWR VGND sg13g2_decap_8
XFILLER_0_960 VPWR VGND sg13g2_decap_8
XFILLER_47_430 VPWR VGND sg13g2_decap_8
XFILLER_48_997 VPWR VGND sg13g2_decap_8
XFILLER_19_176 VPWR VGND sg13g2_fill_1
XFILLER_19_198 VPWR VGND sg13g2_decap_4
XFILLER_35_625 VPWR VGND sg13g2_decap_8
XFILLER_16_872 VPWR VGND sg13g2_decap_8
X_2951_ sap_3_inst.alu.tmp\[4\] net750 _0477_ _0514_ VPWR VGND sg13g2_a21o_1
XFILLER_31_820 VPWR VGND sg13g2_decap_8
XFILLER_43_691 VPWR VGND sg13g2_decap_8
XFILLER_15_393 VPWR VGND sg13g2_fill_2
X_2882_ sap_3_inst.alu.tmp\[4\] net750 _0447_ VPWR VGND sg13g2_xor2_1
XFILLER_31_897 VPWR VGND sg13g2_decap_8
X_3503_ _1032_ _0751_ _0855_ VPWR VGND sg13g2_xnor2_1
X_3434_ _0965_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] net587 VPWR
+ VGND sg13g2_nand2_1
XFILLER_44_1004 VPWR VGND sg13g2_decap_8
X_3365_ _0899_ net577 _0898_ VPWR VGND sg13g2_nand2_1
X_2316_ _1737_ net739 _1701_ VPWR VGND sg13g2_nand2_1
X_3296_ VGND VPWR _1589_ _0676_ _0832_ _1657_ sg13g2_a21oi_1
X_2247_ _1650_ _1653_ _1645_ _1668_ VPWR VGND _1667_ sg13g2_nand4_1
XFILLER_39_964 VPWR VGND sg13g2_decap_8
X_2178_ net738 _1517_ _1562_ _1599_ VPWR VGND sg13g2_nor3_2
XFILLER_26_625 VPWR VGND sg13g2_decap_8
XFILLER_22_820 VPWR VGND sg13g2_decap_8
XFILLER_25_179 VPWR VGND sg13g2_fill_1
XFILLER_22_897 VPWR VGND sg13g2_decap_8
XFILLER_21_374 VPWR VGND sg13g2_fill_2
XFILLER_1_702 VPWR VGND sg13g2_decap_8
Xoutput24 net24 uio_out[7] VPWR VGND sg13g2_buf_1
Xoutput13 net13 uio_oe[4] VPWR VGND sg13g2_buf_1
XFILLER_49_717 VPWR VGND sg13g2_decap_8
XFILLER_1_779 VPWR VGND sg13g2_decap_8
XFILLER_5_1020 VPWR VGND sg13g2_decap_8
XFILLER_45_912 VPWR VGND sg13g2_decap_8
XFILLER_17_647 VPWR VGND sg13g2_decap_8
XFILLER_29_496 VPWR VGND sg13g2_decap_8
XFILLER_45_989 VPWR VGND sg13g2_decap_8
XFILLER_44_444 VPWR VGND sg13g2_decap_8
XFILLER_16_146 VPWR VGND sg13g2_fill_1
XFILLER_13_831 VPWR VGND sg13g2_decap_8
XFILLER_9_824 VPWR VGND sg13g2_decap_8
XFILLER_40_683 VPWR VGND sg13g2_decap_8
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_4_551 VPWR VGND sg13g2_decap_8
X_3150_ net680 _0685_ _0686_ VPWR VGND sg13g2_nor2b_1
X_2101_ net735 net737 _1522_ VPWR VGND sg13g2_nor2_2
X_3081_ net695 _1588_ _1622_ _0617_ VPWR VGND sg13g2_nor3_1
X_2032_ _1455_ net757 VPWR VGND sg13g2_inv_2
XFILLER_48_794 VPWR VGND sg13g2_decap_8
XFILLER_36_934 VPWR VGND sg13g2_decap_8
XFILLER_35_499 VPWR VGND sg13g2_decap_8
X_3983_ _0488_ net748 net663 _1403_ VPWR VGND sg13g2_mux2_1
X_2934_ VPWR VGND _0497_ _0310_ _0496_ sap_3_inst.alu.act\[5\] _0498_ net669 sg13g2_a221oi_1
X_2865_ _0431_ _0423_ _0429_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_694 VPWR VGND sg13g2_decap_8
X_2796_ net618 _0197_ _0353_ _0364_ VPWR VGND sg13g2_nor3_1
X_3417_ _0949_ _1920_ net571 VPWR VGND sg13g2_nand2_1
X_3348_ _0883_ _0827_ _0872_ VPWR VGND sg13g2_xnor2_1
X_3279_ _0658_ _0671_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] _0815_
+ VPWR VGND net659 sg13g2_nand4_1
XFILLER_39_761 VPWR VGND sg13g2_decap_8
XFILLER_26_422 VPWR VGND sg13g2_decap_8
XFILLER_27_956 VPWR VGND sg13g2_decap_8
XFILLER_42_937 VPWR VGND sg13g2_decap_8
XFILLER_14_628 VPWR VGND sg13g2_decap_8
XFILLER_26_68 VPWR VGND sg13g2_fill_2
XFILLER_26_499 VPWR VGND sg13g2_decap_8
XFILLER_41_458 VPWR VGND sg13g2_decap_8
XFILLER_13_127 VPWR VGND sg13g2_fill_2
XFILLER_22_694 VPWR VGND sg13g2_decap_8
XFILLER_6_827 VPWR VGND sg13g2_decap_8
XFILLER_10_867 VPWR VGND sg13g2_decap_8
XFILLER_49_514 VPWR VGND sg13g2_decap_8
XFILLER_1_576 VPWR VGND sg13g2_decap_8
XFILLER_18_901 VPWR VGND sg13g2_decap_8
XFILLER_37_709 VPWR VGND sg13g2_decap_8
XFILLER_18_978 VPWR VGND sg13g2_decap_8
XFILLER_45_786 VPWR VGND sg13g2_decap_8
XFILLER_40_480 VPWR VGND sg13g2_decap_8
XFILLER_9_621 VPWR VGND sg13g2_decap_8
X_2650_ _0242_ _0244_ _0241_ _0245_ VPWR VGND sg13g2_nand3_1
XFILLER_8_186 VPWR VGND sg13g2_fill_1
XFILLER_9_698 VPWR VGND sg13g2_decap_8
X_2581_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] net622
+ net624 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] _1992_ net679 sg13g2_a221oi_1
X_3202_ _0713_ _0720_ _0738_ VPWR VGND sg13g2_nor2_1
XFILLER_41_1018 VPWR VGND sg13g2_decap_8
X_4182_ net799 VGND VPWR net76 regFile_serial_start clknet_3_6__leaf_clk sg13g2_dfrbpq_1
X_3133_ net702 VPWR _0669_ VGND _0665_ _0668_ sg13g2_o21ai_1
X_3064_ _1635_ net684 _0600_ VPWR VGND sg13g2_nor2_1
XFILLER_48_591 VPWR VGND sg13g2_decap_8
X_2015_ _1438_ net729 VPWR VGND sg13g2_inv_2
XFILLER_24_904 VPWR VGND sg13g2_decap_8
XFILLER_36_731 VPWR VGND sg13g2_decap_8
X_3966_ _1391_ _1390_ _1845_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_458 VPWR VGND sg13g2_decap_8
X_2917_ _0481_ _0476_ _0480_ VPWR VGND sg13g2_nand2_1
X_3897_ _1336_ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] _1302_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_31_491 VPWR VGND sg13g2_decap_8
X_2848_ _0414_ _0410_ _0412_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_808 VPWR VGND sg13g2_decap_8
X_2779_ _0348_ _0336_ _0341_ VPWR VGND sg13g2_nand2_1
Xfanout622 _1802_ net622 VPWR VGND sg13g2_buf_8
Xfanout611 _0715_ net611 VPWR VGND sg13g2_buf_8
Xfanout600 _0724_ net600 VPWR VGND sg13g2_buf_8
Xfanout633 net634 net633 VPWR VGND sg13g2_buf_8
Xfanout666 _0632_ net666 VPWR VGND sg13g2_buf_8
Xfanout655 net658 net655 VPWR VGND sg13g2_buf_8
Xfanout644 net645 net644 VPWR VGND sg13g2_buf_1
Xfanout688 _1558_ net688 VPWR VGND sg13g2_buf_8
Xfanout699 net700 net699 VPWR VGND sg13g2_buf_1
Xfanout677 net679 net677 VPWR VGND sg13g2_buf_8
XFILLER_46_528 VPWR VGND sg13g2_decap_8
XFILLER_2_1001 VPWR VGND sg13g2_decap_8
XFILLER_27_753 VPWR VGND sg13g2_decap_8
XFILLER_42_734 VPWR VGND sg13g2_decap_8
XFILLER_15_948 VPWR VGND sg13g2_decap_8
XFILLER_22_491 VPWR VGND sg13g2_decap_8
XFILLER_6_624 VPWR VGND sg13g2_decap_8
XFILLER_10_664 VPWR VGND sg13g2_decap_8
XFILLER_49_311 VPWR VGND sg13g2_decap_8
XFILLER_2_896 VPWR VGND sg13g2_decap_8
XFILLER_37_506 VPWR VGND sg13g2_decap_8
XFILLER_49_388 VPWR VGND sg13g2_decap_8
XFILLER_18_775 VPWR VGND sg13g2_decap_8
XFILLER_45_583 VPWR VGND sg13g2_decap_8
XFILLER_32_222 VPWR VGND sg13g2_fill_1
X_3820_ _1271_ net606 _1112_ VPWR VGND sg13g2_nand2_1
XFILLER_33_767 VPWR VGND sg13g2_decap_8
XFILLER_14_992 VPWR VGND sg13g2_decap_8
X_3751_ net601 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] _1222_ _0131_
+ VPWR VGND sg13g2_a21o_1
X_2702_ net565 _1866_ net15 VPWR VGND sg13g2_nor2b_2
X_3682_ _1174_ VPWR _1179_ VGND _1176_ _1178_ sg13g2_o21ai_1
XFILLER_9_495 VPWR VGND sg13g2_decap_8
X_2633_ _0027_ _0205_ _0228_ VPWR VGND sg13g2_nand2_1
X_2564_ net743 net675 _1976_ VPWR VGND sg13g2_nor2_1
X_2495_ _1910_ net5 _1847_ VPWR VGND sg13g2_nand2_1
X_4165_ net779 VGND VPWR _0143_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\]
+ clknet_5_14__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3116_ _0649_ _0641_ _0651_ _0652_ VPWR VGND sg13g2_a21o_2
X_4096_ net775 VGND VPWR _0074_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[7\]
+ clknet_5_10__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
XFILLER_43_509 VPWR VGND sg13g2_decap_8
X_3047_ net31 sap_3_inst.controller.opcode\[0\] net692 _0059_ VPWR VGND sg13g2_mux2_1
XFILLER_24_701 VPWR VGND sg13g2_decap_8
XFILLER_24_778 VPWR VGND sg13g2_decap_8
X_3949_ VPWR VGND _1382_ net765 _1379_ _1490_ _1383_ net763 sg13g2_a221oi_1
XFILLER_20_940 VPWR VGND sg13g2_decap_8
XFILLER_3_605 VPWR VGND sg13g2_decap_8
XFILLER_24_1002 VPWR VGND sg13g2_decap_8
XFILLER_47_815 VPWR VGND sg13g2_decap_8
XFILLER_46_358 VPWR VGND sg13g2_decap_4
XFILLER_0_29 VPWR VGND sg13g2_decap_8
XFILLER_27_550 VPWR VGND sg13g2_decap_8
XFILLER_42_531 VPWR VGND sg13g2_decap_8
XFILLER_14_222 VPWR VGND sg13g2_fill_1
XFILLER_15_745 VPWR VGND sg13g2_decap_8
XFILLER_30_759 VPWR VGND sg13g2_decap_8
XFILLER_7_944 VPWR VGND sg13g2_decap_8
XFILLER_10_450 VPWR VGND sg13g2_fill_1
XFILLER_11_984 VPWR VGND sg13g2_decap_8
XFILLER_6_498 VPWR VGND sg13g2_decap_8
XFILLER_2_693 VPWR VGND sg13g2_decap_8
X_2280_ _1544_ net709 _1701_ VPWR VGND sg13g2_and2_1
XFILLER_38_837 VPWR VGND sg13g2_decap_8
XFILLER_46_892 VPWR VGND sg13g2_decap_8
XFILLER_45_380 VPWR VGND sg13g2_decap_8
XFILLER_18_572 VPWR VGND sg13g2_decap_8
XFILLER_33_564 VPWR VGND sg13g2_decap_8
XFILLER_21_737 VPWR VGND sg13g2_decap_8
X_3803_ net9 _1138_ _1258_ _1259_ VPWR VGND sg13g2_nor3_1
X_3734_ _1184_ _1185_ net556 _1213_ VPWR VGND sg13g2_nor3_1
X_3665_ VGND VPWR _1899_ net568 _1164_ _1163_ sg13g2_a21oi_1
Xclkbuf_4_15_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_15_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2616_ _0213_ _0209_ _0212_ net637 _1457_ VPWR VGND sg13g2_a22oi_1
X_3596_ _1105_ _1107_ _1110_ _1111_ VPWR VGND sg13g2_nor3_1
X_2547_ _1960_ net620 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] net630
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2478_ _1895_ net619 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] net627
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4217_ net788 VGND VPWR _0194_ u_ser.bit_pos\[0\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_29_804 VPWR VGND sg13g2_decap_8
X_4148_ net795 VGND VPWR _0126_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\]
+ clknet_5_28__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_44_829 VPWR VGND sg13g2_decap_8
X_4079_ net791 VGND VPWR _0057_ sap_3_inst.alu.tmp\[6\] clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_37_870 VPWR VGND sg13g2_decap_8
XFILLER_24_575 VPWR VGND sg13g2_decap_8
XFILLER_7_229 VPWR VGND sg13g2_fill_1
Xclkload1 VPWR clkload1/Y clknet_3_1__leaf_clk VGND sg13g2_inv_1
XFILLER_3_402 VPWR VGND sg13g2_fill_1
XFILLER_4_936 VPWR VGND sg13g2_decap_8
XFILLER_3_479 VPWR VGND sg13g2_decap_8
XFILLER_47_612 VPWR VGND sg13g2_decap_8
XFILLER_47_689 VPWR VGND sg13g2_decap_8
XFILLER_35_807 VPWR VGND sg13g2_decap_8
XFILLER_15_542 VPWR VGND sg13g2_decap_8
XFILLER_43_873 VPWR VGND sg13g2_decap_8
XFILLER_30_556 VPWR VGND sg13g2_decap_8
XFILLER_7_741 VPWR VGND sg13g2_decap_8
XFILLER_11_781 VPWR VGND sg13g2_decap_8
X_3450_ _0981_ _0980_ _0977_ VPWR VGND sg13g2_nand2b_1
X_2401_ _1822_ _1540_ _1577_ VPWR VGND sg13g2_nand2_1
X_3381_ _0911_ _0912_ net611 _0914_ VPWR VGND _0913_ sg13g2_nand4_1
X_2332_ _1607_ _1658_ _1753_ VPWR VGND sg13g2_nor2_1
XFILLER_2_490 VPWR VGND sg13g2_decap_8
Xclkbuf_4_7_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_7_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_4002_ _1410_ _1417_ u_ser.bit_pos\[2\] _1418_ VPWR VGND sg13g2_nand3_1
X_2263_ VGND VPWR _1684_ _1630_ net700 sg13g2_or2_1
X_2194_ _1609_ _1614_ _1615_ VPWR VGND sg13g2_and2_1
XFILLER_38_634 VPWR VGND sg13g2_decap_8
XFILLER_26_807 VPWR VGND sg13g2_decap_8
XFILLER_37_188 VPWR VGND sg13g2_fill_1
XFILLER_34_851 VPWR VGND sg13g2_decap_8
X_4034__12 VPWR net46 clknet_leaf_1_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_21_534 VPWR VGND sg13g2_decap_8
XFILLER_33_394 VPWR VGND sg13g2_fill_1
X_3717_ _1198_ VPWR _0117_ VGND _1201_ _1202_ sg13g2_o21ai_1
X_3648_ _1149_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] net597 VPWR
+ VGND sg13g2_nand2_1
X_4030__8 VPWR net42 clknet_leaf_3_sap_3_inst.alu.clk VGND sg13g2_inv_1
X_3579_ _1096_ _1078_ net12 VPWR VGND sg13g2_nand2b_1
XFILLER_48_409 VPWR VGND sg13g2_decap_8
XFILLER_0_449 VPWR VGND sg13g2_decap_8
Xhold13 u_ser.shadow_reg\[7\] VPWR VGND net60 sg13g2_dlygate4sd3_1
Xhold35 sap_3_inst.reg_file.array_serializer_inst.word_index\[0\] VPWR VGND net82
+ sg13g2_dlygate4sd3_1
Xhold24 u_ser.bit_pos\[1\] VPWR VGND net71 sg13g2_dlygate4sd3_1
XFILLER_29_601 VPWR VGND sg13g2_decap_8
XFILLER_17_829 VPWR VGND sg13g2_decap_8
XFILLER_29_678 VPWR VGND sg13g2_decap_8
XFILLER_44_626 VPWR VGND sg13g2_decap_8
XFILLER_28_199 VPWR VGND sg13g2_fill_2
XFILLER_24_350 VPWR VGND sg13g2_fill_2
XFILLER_25_884 VPWR VGND sg13g2_decap_8
XFILLER_40_865 VPWR VGND sg13g2_decap_8
XFILLER_12_567 VPWR VGND sg13g2_decap_8
XFILLER_8_538 VPWR VGND sg13g2_decap_8
XFILLER_4_733 VPWR VGND sg13g2_decap_8
XFILLER_20_9 VPWR VGND sg13g2_fill_2
XFILLER_48_976 VPWR VGND sg13g2_decap_8
XFILLER_19_155 VPWR VGND sg13g2_fill_2
XFILLER_35_604 VPWR VGND sg13g2_decap_8
XFILLER_47_486 VPWR VGND sg13g2_decap_8
XFILLER_16_851 VPWR VGND sg13g2_decap_8
XFILLER_43_670 VPWR VGND sg13g2_decap_8
X_2950_ VGND VPWR _0511_ _0512_ _0513_ _2007_ sg13g2_a21oi_1
X_2881_ _0446_ net750 sap_3_inst.alu.tmp\[4\] _0340_ VPWR VGND sg13g2_and3_1
XFILLER_31_876 VPWR VGND sg13g2_decap_8
X_3502_ net24 net16 _0838_ _1031_ VPWR VGND sg13g2_mux2_1
X_3433_ _0961_ _0962_ net610 _0964_ VPWR VGND _0963_ sg13g2_nand4_1
X_3364_ _0896_ _0897_ _0898_ VPWR VGND sg13g2_and2_1
X_2315_ net689 _1717_ net732 _1736_ VPWR VGND sg13g2_nand3_1
X_3295_ _0797_ _0828_ net614 _0831_ VPWR VGND sg13g2_mux2_1
X_2246_ _1654_ _1660_ _1663_ _1666_ _1667_ VPWR VGND sg13g2_nor4_1
XFILLER_39_943 VPWR VGND sg13g2_decap_8
XFILLER_26_604 VPWR VGND sg13g2_decap_8
X_2177_ _1598_ _1516_ _1561_ VPWR VGND sg13g2_nand2_1
XFILLER_22_876 VPWR VGND sg13g2_decap_8
Xoutput25 net25 uo_out[0] VPWR VGND sg13g2_buf_1
Xoutput14 net14 uio_oe[5] VPWR VGND sg13g2_buf_1
XFILLER_1_758 VPWR VGND sg13g2_decap_8
XFILLER_44_423 VPWR VGND sg13g2_decap_8
XFILLER_17_626 VPWR VGND sg13g2_decap_8
XFILLER_29_475 VPWR VGND sg13g2_decap_8
XFILLER_45_968 VPWR VGND sg13g2_decap_8
XFILLER_13_810 VPWR VGND sg13g2_decap_8
XFILLER_31_106 VPWR VGND sg13g2_fill_2
XFILLER_25_681 VPWR VGND sg13g2_decap_8
XFILLER_40_662 VPWR VGND sg13g2_decap_8
XFILLER_9_803 VPWR VGND sg13g2_decap_8
XFILLER_13_887 VPWR VGND sg13g2_decap_8
XFILLER_4_530 VPWR VGND sg13g2_decap_8
Xclkbuf_5_26__f_sap_3_inst.alu.clk_regs clknet_4_13_0_sap_3_inst.alu.clk_regs clknet_5_26__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2100_ VGND VPWR _1521_ net728 net726 sg13g2_or2_1
X_3080_ net687 VPWR _0616_ VGND _1587_ _1592_ sg13g2_o21ai_1
XFILLER_48_773 VPWR VGND sg13g2_decap_8
X_2031_ _1454_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] VPWR VGND
+ sg13g2_inv_2
XFILLER_36_913 VPWR VGND sg13g2_decap_8
X_3982_ _1402_ sap_3_inst.alu.act\[4\] net548 _0182_ VPWR VGND sg13g2_mux2_1
XFILLER_44_990 VPWR VGND sg13g2_decap_8
X_2933_ VGND VPWR net543 _0491_ _0497_ _0314_ sg13g2_a21oi_1
X_2864_ _0423_ _0429_ _0430_ VPWR VGND sg13g2_nor2_1
XFILLER_31_673 VPWR VGND sg13g2_decap_8
X_2795_ VPWR VGND _0322_ _0362_ _0358_ net563 _0363_ _0354_ sg13g2_a221oi_1
XFILLER_7_60 VPWR VGND sg13g2_decap_8
XFILLER_11_1026 VPWR VGND sg13g2_fill_2
X_3416_ _0946_ _0947_ net610 _0948_ VPWR VGND sg13g2_mux2_1
X_3347_ _0882_ net553 _0825_ _0881_ VPWR VGND sg13g2_and3_2
X_3278_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] _0813_
+ net656 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] _0814_ net608 sg13g2_a221oi_1
XFILLER_39_740 VPWR VGND sg13g2_decap_8
X_2229_ _1650_ _1587_ _1649_ VPWR VGND sg13g2_nand2_1
XFILLER_26_401 VPWR VGND sg13g2_decap_8
XFILLER_27_935 VPWR VGND sg13g2_decap_8
XFILLER_42_916 VPWR VGND sg13g2_decap_8
XFILLER_13_106 VPWR VGND sg13g2_fill_1
XFILLER_14_607 VPWR VGND sg13g2_decap_8
XFILLER_26_478 VPWR VGND sg13g2_decap_8
XFILLER_22_673 VPWR VGND sg13g2_decap_8
XFILLER_6_806 VPWR VGND sg13g2_decap_8
XFILLER_10_846 VPWR VGND sg13g2_decap_8
XFILLER_1_555 VPWR VGND sg13g2_decap_8
XFILLER_18_957 VPWR VGND sg13g2_decap_8
XFILLER_45_765 VPWR VGND sg13g2_decap_8
XFILLER_33_949 VPWR VGND sg13g2_decap_8
XFILLER_9_600 VPWR VGND sg13g2_decap_8
XFILLER_13_684 VPWR VGND sg13g2_decap_8
XFILLER_34_1026 VPWR VGND sg13g2_fill_2
XFILLER_9_677 VPWR VGND sg13g2_decap_8
X_2580_ _1991_ _1989_ _1990_ VPWR VGND sg13g2_nand2_1
XFILLER_5_894 VPWR VGND sg13g2_decap_8
X_3201_ _0691_ _0694_ _0711_ _0728_ _0737_ VPWR VGND sg13g2_and4_1
X_4181_ net799 VGND VPWR net64 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_2
X_3132_ _0661_ VPWR _0668_ VGND _1675_ _0667_ sg13g2_o21ai_1
XFILLER_48_570 VPWR VGND sg13g2_decap_8
X_3063_ net706 VPWR _0599_ VGND _1577_ _1638_ sg13g2_o21ai_1
XFILLER_36_710 VPWR VGND sg13g2_decap_8
X_2014_ _1437_ net732 VPWR VGND sg13g2_inv_2
XFILLER_36_787 VPWR VGND sg13g2_decap_8
XFILLER_17_990 VPWR VGND sg13g2_decap_8
X_3965_ _0299_ _0301_ net683 _1390_ VPWR VGND sg13g2_nand3_1
X_2916_ _0480_ _0479_ _0333_ _0477_ _0340_ VPWR VGND sg13g2_a22oi_1
X_3896_ net764 net53 _1335_ _0163_ VPWR VGND sg13g2_a21o_1
X_2847_ VGND VPWR _0399_ _0403_ _0413_ _0411_ sg13g2_a21oi_1
X_2778_ VPWR VGND net757 net670 net572 _0337_ _0347_ net573 sg13g2_a221oi_1
Xfanout612 net613 net612 VPWR VGND sg13g2_buf_8
Xfanout601 _0724_ net601 VPWR VGND sg13g2_buf_1
Xfanout623 net624 net623 VPWR VGND sg13g2_buf_8
Xfanout667 net668 net667 VPWR VGND sg13g2_buf_8
Xfanout645 _0733_ net645 VPWR VGND sg13g2_buf_8
Xfanout656 net658 net656 VPWR VGND sg13g2_buf_8
Xfanout634 _1796_ net634 VPWR VGND sg13g2_buf_8
XFILLER_46_507 VPWR VGND sg13g2_decap_8
Xfanout689 _1552_ net689 VPWR VGND sg13g2_buf_8
Xfanout678 net679 net678 VPWR VGND sg13g2_buf_1
XFILLER_27_732 VPWR VGND sg13g2_decap_8
XFILLER_42_713 VPWR VGND sg13g2_decap_8
XFILLER_15_927 VPWR VGND sg13g2_decap_8
XFILLER_14_415 VPWR VGND sg13g2_fill_1
XFILLER_22_470 VPWR VGND sg13g2_decap_8
XFILLER_6_603 VPWR VGND sg13g2_decap_8
XFILLER_10_643 VPWR VGND sg13g2_decap_8
XFILLER_5_113 VPWR VGND sg13g2_fill_2
XFILLER_5_168 VPWR VGND sg13g2_fill_1
XFILLER_5_157 VPWR VGND sg13g2_fill_2
XFILLER_2_875 VPWR VGND sg13g2_decap_8
XFILLER_49_367 VPWR VGND sg13g2_decap_8
XFILLER_18_754 VPWR VGND sg13g2_decap_8
XFILLER_45_562 VPWR VGND sg13g2_decap_8
XFILLER_33_746 VPWR VGND sg13g2_decap_8
XFILLER_21_919 VPWR VGND sg13g2_decap_8
XFILLER_14_971 VPWR VGND sg13g2_decap_8
XFILLER_32_289 VPWR VGND sg13g2_fill_1
X_3750_ VGND VPWR _1220_ _1221_ _1222_ _1218_ sg13g2_a21oi_1
X_2701_ net565 _1887_ net14 VPWR VGND sg13g2_nor2b_2
X_3681_ _1027_ _1177_ _1178_ VPWR VGND sg13g2_nor2_1
X_2632_ _0227_ VPWR _0228_ VGND _1858_ net32 sg13g2_o21ai_1
X_2563_ VPWR net20 net546 VGND sg13g2_inv_1
XFILLER_5_691 VPWR VGND sg13g2_decap_8
X_2494_ _1909_ _1828_ sap_3_inst.alu.flags\[4\] _1827_ net751 VPWR VGND sg13g2_a22oi_1
XFILLER_4_94 VPWR VGND sg13g2_fill_1
XFILLER_4_72 VPWR VGND sg13g2_fill_2
X_4164_ net794 VGND VPWR _0142_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\]
+ clknet_5_28__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3115_ _1515_ VPWR _0651_ VGND net682 _0650_ sg13g2_o21ai_1
X_4095_ net780 VGND VPWR _0073_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[6\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
X_3046_ net24 sap_3_inst.alu.tmp\[7\] net668 _0058_ VPWR VGND sg13g2_mux2_1
XFILLER_36_584 VPWR VGND sg13g2_decap_8
XFILLER_24_757 VPWR VGND sg13g2_decap_8
X_3948_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] _1381_
+ net721 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] _1382_ _1308_ sg13g2_a221oi_1
X_3879_ _1320_ _1311_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] _1302_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_996 VPWR VGND sg13g2_decap_8
XFILLER_42_510 VPWR VGND sg13g2_decap_8
XFILLER_15_724 VPWR VGND sg13g2_decap_8
XFILLER_42_587 VPWR VGND sg13g2_decap_8
XFILLER_30_738 VPWR VGND sg13g2_decap_8
XFILLER_7_923 VPWR VGND sg13g2_decap_8
XFILLER_11_963 VPWR VGND sg13g2_decap_8
XFILLER_2_672 VPWR VGND sg13g2_decap_8
XFILLER_38_816 VPWR VGND sg13g2_decap_8
XFILLER_46_871 VPWR VGND sg13g2_decap_8
XFILLER_18_551 VPWR VGND sg13g2_decap_8
XFILLER_33_543 VPWR VGND sg13g2_decap_8
XFILLER_21_716 VPWR VGND sg13g2_decap_8
X_3802_ net608 _1038_ _1258_ VPWR VGND sg13g2_nor2_1
X_3733_ net556 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] _1212_ _0123_
+ VPWR VGND sg13g2_a21o_1
X_3664_ net14 net568 _1163_ VPWR VGND sg13g2_nor2_1
X_2615_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] _0211_
+ net634 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] _0212_ net679 sg13g2_a221oi_1
X_3595_ VGND VPWR _1110_ _1109_ net578 sg13g2_or2_1
XFILLER_47_1025 VPWR VGND sg13g2_decap_4
X_2546_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] net637
+ net624 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\] _1959_ net678 sg13g2_a221oi_1
X_2477_ _1894_ net625 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] net633
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4216_ net797 VGND VPWR _0193_ sap_3_inst.reg_file.array_serializer_inst.word_index\[3\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_2
Xclkbuf_5_0__f_sap_3_inst.alu.clk_regs clknet_4_0_0_sap_3_inst.alu.clk_regs clknet_5_0__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_4147_ net793 VGND VPWR _0125_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\]
+ clknet_5_25__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_44_808 VPWR VGND sg13g2_decap_8
X_4078_ net791 VGND VPWR _0056_ sap_3_inst.alu.tmp\[5\] clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3029_ _0568_ _0573_ _0582_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_554 VPWR VGND sg13g2_decap_8
XFILLER_12_749 VPWR VGND sg13g2_decap_8
Xclkload2 clknet_3_2__leaf_clk clkload2/X VPWR VGND sg13g2_buf_1
XFILLER_20_793 VPWR VGND sg13g2_decap_8
XFILLER_4_915 VPWR VGND sg13g2_decap_8
XFILLER_3_458 VPWR VGND sg13g2_decap_8
XFILLER_47_668 VPWR VGND sg13g2_decap_8
XFILLER_15_521 VPWR VGND sg13g2_decap_8
XFILLER_43_852 VPWR VGND sg13g2_decap_8
XFILLER_42_351 VPWR VGND sg13g2_fill_1
XFILLER_42_395 VPWR VGND sg13g2_fill_2
XFILLER_15_598 VPWR VGND sg13g2_decap_8
XFILLER_30_535 VPWR VGND sg13g2_decap_8
XFILLER_11_760 VPWR VGND sg13g2_decap_8
XFILLER_7_720 VPWR VGND sg13g2_decap_8
XFILLER_7_797 VPWR VGND sg13g2_decap_8
X_2400_ net695 _1565_ _1821_ VPWR VGND sg13g2_nor2_1
X_3380_ _0913_ net645 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] net650
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2331_ net724 net698 net735 _1752_ VPWR VGND _1549_ sg13g2_nand4_1
X_2262_ _1682_ VPWR _1683_ VGND _1578_ _1616_ sg13g2_o21ai_1
X_4001_ _1414_ VPWR _1417_ VGND u_ser.bit_pos\[1\] _1416_ sg13g2_o21ai_1
XFILLER_38_613 VPWR VGND sg13g2_decap_8
X_2193_ net731 net729 _1614_ VPWR VGND sg13g2_nor2b_2
XFILLER_25_318 VPWR VGND sg13g2_fill_1
XFILLER_34_830 VPWR VGND sg13g2_decap_8
XFILLER_21_513 VPWR VGND sg13g2_decap_8
XFILLER_14_1013 VPWR VGND sg13g2_decap_8
X_3716_ net645 VPWR _1202_ VGND net576 _0898_ sg13g2_o21ai_1
X_3647_ _0101_ _0901_ _1148_ net596 _1451_ VPWR VGND sg13g2_a22oi_1
X_3578_ _1095_ net546 net570 VPWR VGND sg13g2_nand2_1
X_2529_ _1551_ _1925_ net730 _1942_ VPWR VGND sg13g2_nand3_1
Xhold14 u_ser.shadow_reg\[1\] VPWR VGND net61 sg13g2_dlygate4sd3_1
Xhold25 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\] VPWR VGND net72 sg13g2_dlygate4sd3_1
XFILLER_21_1017 VPWR VGND sg13g2_decap_8
XFILLER_44_605 VPWR VGND sg13g2_decap_8
XFILLER_17_808 VPWR VGND sg13g2_decap_8
XFILLER_21_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_657 VPWR VGND sg13g2_decap_8
XFILLER_16_329 VPWR VGND sg13g2_fill_2
XFILLER_25_863 VPWR VGND sg13g2_decap_8
XFILLER_40_844 VPWR VGND sg13g2_decap_8
XFILLER_12_546 VPWR VGND sg13g2_decap_8
XFILLER_8_517 VPWR VGND sg13g2_decap_8
XFILLER_6_29 VPWR VGND sg13g2_fill_1
XFILLER_20_590 VPWR VGND sg13g2_decap_8
XFILLER_4_712 VPWR VGND sg13g2_decap_8
XFILLER_3_211 VPWR VGND sg13g2_fill_1
XFILLER_4_789 VPWR VGND sg13g2_decap_8
XFILLER_48_955 VPWR VGND sg13g2_decap_8
XFILLER_0_995 VPWR VGND sg13g2_decap_8
XFILLER_47_465 VPWR VGND sg13g2_decap_8
XFILLER_16_830 VPWR VGND sg13g2_decap_8
XFILLER_37_1024 VPWR VGND sg13g2_decap_4
X_2880_ _0443_ _0442_ _1937_ _0445_ VPWR VGND sg13g2_a21o_1
XFILLER_31_855 VPWR VGND sg13g2_decap_8
X_3501_ _1027_ net613 _1029_ _1030_ VPWR VGND sg13g2_a21o_1
XFILLER_7_594 VPWR VGND sg13g2_decap_8
X_3432_ _0963_ net646 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] net649
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] VPWR VGND sg13g2_a22oi_1
X_3363_ _0857_ _0872_ _0797_ _0897_ VPWR VGND _0895_ sg13g2_nand4_1
X_2314_ _1735_ _1734_ _1631_ _1724_ _1618_ VPWR VGND sg13g2_a22oi_1
X_3294_ _0830_ net666 VPWR VGND net660 sg13g2_nand2b_2
X_2245_ _1666_ _1665_ _1604_ _1636_ net694 VPWR VGND sg13g2_a22oi_1
XFILLER_39_922 VPWR VGND sg13g2_decap_8
X_2176_ net737 _1519_ _1562_ _1595_ _1597_ VPWR VGND sg13g2_or4_1
XFILLER_38_487 VPWR VGND sg13g2_decap_8
XFILLER_39_999 VPWR VGND sg13g2_decap_8
XFILLER_41_619 VPWR VGND sg13g2_decap_8
XFILLER_40_107 VPWR VGND sg13g2_fill_1
XFILLER_22_855 VPWR VGND sg13g2_decap_8
XFILLER_21_376 VPWR VGND sg13g2_fill_1
XFILLER_5_509 VPWR VGND sg13g2_decap_8
XFILLER_31_48 VPWR VGND sg13g2_fill_1
Xoutput15 net15 uio_oe[6] VPWR VGND sg13g2_buf_1
Xoutput26 net26 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_737 VPWR VGND sg13g2_decap_8
XFILLER_29_410 VPWR VGND sg13g2_fill_1
XFILLER_29_454 VPWR VGND sg13g2_decap_8
XFILLER_45_947 VPWR VGND sg13g2_decap_8
XFILLER_44_402 VPWR VGND sg13g2_decap_8
XFILLER_17_605 VPWR VGND sg13g2_decap_8
XFILLER_44_479 VPWR VGND sg13g2_decap_8
XFILLER_25_660 VPWR VGND sg13g2_decap_8
XFILLER_24_181 VPWR VGND sg13g2_fill_2
XFILLER_40_641 VPWR VGND sg13g2_decap_8
XFILLER_13_866 VPWR VGND sg13g2_decap_8
XFILLER_9_859 VPWR VGND sg13g2_decap_8
XFILLER_4_586 VPWR VGND sg13g2_decap_8
XFILLER_0_792 VPWR VGND sg13g2_decap_8
XFILLER_48_752 VPWR VGND sg13g2_decap_8
X_2030_ VPWR _1453_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_36_969 VPWR VGND sg13g2_decap_8
X_3981_ _0458_ net750 net663 _1402_ VPWR VGND sg13g2_mux2_1
XFILLER_23_619 VPWR VGND sg13g2_decap_8
XFILLER_35_457 VPWR VGND sg13g2_fill_2
XFILLER_15_170 VPWR VGND sg13g2_fill_1
X_2932_ _0494_ _0495_ _0475_ _0496_ VPWR VGND sg13g2_nand3_1
XFILLER_31_652 VPWR VGND sg13g2_decap_8
X_2863_ VGND VPWR net755 _1464_ _0429_ _0390_ sg13g2_a21oi_1
X_2794_ _0361_ VPWR _0362_ VGND net757 _0327_ sg13g2_o21ai_1
XFILLER_11_1005 VPWR VGND sg13g2_decap_8
XFILLER_8_881 VPWR VGND sg13g2_decap_8
X_3415_ _0947_ _0775_ _0823_ VPWR VGND sg13g2_xnor2_1
X_3346_ _0744_ _0871_ _0881_ VPWR VGND sg13g2_and2_1
X_3277_ _0810_ _0811_ _0809_ _0813_ VPWR VGND _0812_ sg13g2_nand4_1
X_2228_ _1649_ _1623_ _1648_ VPWR VGND sg13g2_nand2b_1
XFILLER_27_914 VPWR VGND sg13g2_decap_8
XFILLER_39_796 VPWR VGND sg13g2_decap_8
X_2159_ _1580_ net694 _1578_ VPWR VGND sg13g2_nand2_1
XFILLER_26_457 VPWR VGND sg13g2_decap_8
XFILLER_41_438 VPWR VGND sg13g2_fill_2
XFILLER_13_129 VPWR VGND sg13g2_fill_1
XFILLER_22_652 VPWR VGND sg13g2_decap_8
XFILLER_10_825 VPWR VGND sg13g2_decap_8
XFILLER_1_534 VPWR VGND sg13g2_decap_8
XFILLER_27_1012 VPWR VGND sg13g2_decap_8
XFILLER_49_549 VPWR VGND sg13g2_decap_8
XFILLER_18_936 VPWR VGND sg13g2_decap_8
XFILLER_29_251 VPWR VGND sg13g2_fill_1
XFILLER_45_744 VPWR VGND sg13g2_decap_8
XFILLER_44_210 VPWR VGND sg13g2_fill_2
XFILLER_33_928 VPWR VGND sg13g2_decap_8
XFILLER_34_1005 VPWR VGND sg13g2_decap_8
XFILLER_41_983 VPWR VGND sg13g2_decap_8
XFILLER_12_151 VPWR VGND sg13g2_fill_1
XFILLER_13_663 VPWR VGND sg13g2_decap_8
XFILLER_8_122 VPWR VGND sg13g2_fill_1
XFILLER_9_656 VPWR VGND sg13g2_decap_8
XFILLER_5_873 VPWR VGND sg13g2_decap_8
X_3200_ _0725_ _0730_ net610 _0736_ VPWR VGND _0735_ sg13g2_nand4_1
X_4180_ net799 VGND VPWR net73 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_2
X_3131_ _1594_ _1608_ _1609_ _0667_ VPWR VGND sg13g2_nor3_1
X_3062_ net696 _1716_ _1510_ _0598_ VPWR VGND sg13g2_nand3_1
X_2013_ net738 _1436_ VPWR VGND sg13g2_inv_4
XFILLER_36_766 VPWR VGND sg13g2_decap_8
XFILLER_23_438 VPWR VGND sg13g2_decap_8
XFILLER_24_939 VPWR VGND sg13g2_decap_8
X_3964_ net602 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] _1389_ _0177_
+ VPWR VGND sg13g2_a21o_1
X_2915_ _0477_ _0478_ _0479_ VPWR VGND sg13g2_nor2b_2
X_3895_ VPWR VGND _1334_ net765 _1328_ _1457_ _1335_ net762 sg13g2_a221oi_1
XFILLER_32_994 VPWR VGND sg13g2_decap_8
X_2846_ _0412_ net753 net672 VPWR VGND sg13g2_xnor2_1
X_2777_ _0346_ _0343_ _0344_ _0325_ net564 VPWR VGND sg13g2_a22oi_1
Xfanout602 net603 net602 VPWR VGND sg13g2_buf_8
Xfanout624 _1801_ net624 VPWR VGND sg13g2_buf_8
Xfanout613 net614 net613 VPWR VGND sg13g2_buf_2
Xfanout646 net648 net646 VPWR VGND sg13g2_buf_8
Xfanout657 net658 net657 VPWR VGND sg13g2_buf_1
Xfanout635 net636 net635 VPWR VGND sg13g2_buf_8
Xfanout668 _0585_ net668 VPWR VGND sg13g2_buf_8
Xfanout679 _1753_ net679 VPWR VGND sg13g2_buf_8
X_3329_ _0864_ net656 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] net608
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_27_711 VPWR VGND sg13g2_decap_8
XFILLER_39_593 VPWR VGND sg13g2_decap_8
XFILLER_15_906 VPWR VGND sg13g2_decap_8
XFILLER_27_788 VPWR VGND sg13g2_decap_8
XFILLER_42_769 VPWR VGND sg13g2_decap_8
XFILLER_23_983 VPWR VGND sg13g2_decap_8
XFILLER_10_622 VPWR VGND sg13g2_decap_8
XFILLER_6_659 VPWR VGND sg13g2_decap_8
XFILLER_10_699 VPWR VGND sg13g2_decap_8
XFILLER_2_854 VPWR VGND sg13g2_decap_8
XFILLER_49_346 VPWR VGND sg13g2_decap_8
XFILLER_18_733 VPWR VGND sg13g2_decap_8
XFILLER_45_541 VPWR VGND sg13g2_decap_8
XFILLER_33_725 VPWR VGND sg13g2_decap_8
XFILLER_14_950 VPWR VGND sg13g2_decap_8
XFILLER_41_780 VPWR VGND sg13g2_decap_8
X_2700_ net565 _1908_ net13 VPWR VGND sg13g2_nor2b_2
X_3680_ net585 VPWR _1177_ VGND net651 _1028_ sg13g2_o21ai_1
X_2631_ _1940_ _0204_ _0226_ _0227_ VPWR VGND sg13g2_nor3_1
X_2562_ _1975_ _1964_ _1965_ _1974_ VPWR VGND sg13g2_and3_2
XFILLER_5_670 VPWR VGND sg13g2_decap_8
X_2493_ _1908_ _1903_ _1907_ net638 _1468_ VPWR VGND sg13g2_a22oi_1
XFILLER_4_62 VPWR VGND sg13g2_fill_1
X_4163_ net786 VGND VPWR _0141_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4094_ net778 VGND VPWR _0072_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[5\]
+ clknet_5_10__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
X_3114_ VGND VPWR _0598_ _0623_ _0650_ _1437_ sg13g2_a21oi_1
XFILLER_28_519 VPWR VGND sg13g2_decap_8
X_3045_ _0590_ VPWR _0057_ VGND net547 net667 sg13g2_o21ai_1
XFILLER_36_563 VPWR VGND sg13g2_decap_8
XFILLER_24_736 VPWR VGND sg13g2_decap_8
X_3947_ _1377_ _1378_ _1376_ _1381_ VPWR VGND _1380_ sg13g2_nand4_1
XFILLER_17_1011 VPWR VGND sg13g2_decap_8
XFILLER_32_791 VPWR VGND sg13g2_decap_8
XFILLER_20_975 VPWR VGND sg13g2_decap_8
X_3878_ _1319_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] _1306_
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2829_ VPWR VGND _2008_ _0395_ _0393_ _0324_ _0396_ _0388_ sg13g2_a221oi_1
XFILLER_15_703 VPWR VGND sg13g2_decap_8
XFILLER_27_585 VPWR VGND sg13g2_decap_8
XFILLER_14_246 VPWR VGND sg13g2_fill_2
XFILLER_42_566 VPWR VGND sg13g2_decap_8
XFILLER_30_717 VPWR VGND sg13g2_decap_8
XFILLER_11_942 VPWR VGND sg13g2_decap_8
XFILLER_23_780 VPWR VGND sg13g2_decap_8
XFILLER_7_902 VPWR VGND sg13g2_decap_8
XFILLER_10_441 VPWR VGND sg13g2_fill_1
XFILLER_7_979 VPWR VGND sg13g2_decap_8
XFILLER_2_651 VPWR VGND sg13g2_decap_8
XFILLER_36_8 VPWR VGND sg13g2_fill_1
XFILLER_49_187 VPWR VGND sg13g2_fill_2
XFILLER_46_850 VPWR VGND sg13g2_decap_8
XFILLER_18_530 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_33_522 VPWR VGND sg13g2_decap_8
X_3801_ VGND VPWR _1492_ net598 _0146_ _1257_ sg13g2_a21oi_1
XFILLER_33_599 VPWR VGND sg13g2_decap_8
X_3732_ _1040_ _1041_ net556 _1212_ VPWR VGND sg13g2_nor3_1
Xclkload20 VPWR clkload20/Y clknet_5_29__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_3663_ VPWR VGND net596 net583 _0975_ _0971_ _1162_ _0972_ sg13g2_a221oi_1
X_2614_ _0208_ _0210_ _0207_ _0211_ VPWR VGND sg13g2_nand3_1
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
X_3594_ VGND VPWR _0766_ _0853_ _1109_ _1108_ sg13g2_a21oi_1
X_2545_ _1956_ _1957_ _1958_ VPWR VGND sg13g2_and2_1
X_2476_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] net621
+ net629 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] _1893_ net677 sg13g2_a221oi_1
X_4215_ net797 VGND VPWR _0192_ sap_3_inst.reg_file.array_serializer_inst.word_index\[2\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_2
X_4146_ net773 VGND VPWR _0124_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\]
+ clknet_5_6__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_839 VPWR VGND sg13g2_decap_8
X_4077_ net790 VGND VPWR _0055_ sap_3_inst.alu.tmp\[4\] clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3028_ _0566_ _0579_ _0580_ _0581_ VPWR VGND sg13g2_nor3_1
XFILLER_24_533 VPWR VGND sg13g2_decap_8
XFILLER_12_728 VPWR VGND sg13g2_decap_8
Xclkload3 VPWR clkload3/Y clknet_3_3__leaf_clk VGND sg13g2_inv_1
XFILLER_20_772 VPWR VGND sg13g2_decap_8
XFILLER_47_647 VPWR VGND sg13g2_decap_8
XFILLER_28_883 VPWR VGND sg13g2_decap_8
XFILLER_43_831 VPWR VGND sg13g2_decap_8
XFILLER_15_577 VPWR VGND sg13g2_decap_8
XFILLER_30_514 VPWR VGND sg13g2_decap_8
XFILLER_7_776 VPWR VGND sg13g2_decap_8
X_2330_ net733 _1750_ _1751_ VPWR VGND sg13g2_nor2_1
X_2261_ net684 VPWR _1682_ VGND net706 _1655_ sg13g2_o21ai_1
X_4000_ _1415_ VPWR _1416_ VGND u_ser.bit_pos\[0\] u_ser.shadow_reg\[5\] sg13g2_o21ai_1
X_2192_ _1590_ _1610_ _1554_ _1613_ VPWR VGND _1612_ sg13g2_nand4_1
XFILLER_37_102 VPWR VGND sg13g2_fill_2
X_2077__2 VPWR net36 clknet_leaf_2_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_38_669 VPWR VGND sg13g2_decap_8
XFILLER_19_894 VPWR VGND sg13g2_decap_8
XFILLER_34_886 VPWR VGND sg13g2_decap_8
XFILLER_21_569 VPWR VGND sg13g2_decap_8
X_3715_ net19 net580 _1200_ _1201_ VPWR VGND sg13g2_nor3_1
X_3646_ net596 _1147_ _1148_ VPWR VGND sg13g2_nor2_1
X_3577_ _1094_ net590 _0935_ VPWR VGND sg13g2_nand2_1
XFILLER_1_919 VPWR VGND sg13g2_decap_8
X_2528_ net725 _1508_ net729 _1941_ VPWR VGND net688 sg13g2_nand4_1
Xhold15 u_ser.shadow_reg\[2\] VPWR VGND net62 sg13g2_dlygate4sd3_1
X_2459_ VGND VPWR _1877_ _1878_ _1866_ _1723_ sg13g2_a21oi_2
Xhold26 _0158_ VPWR VGND net73 sg13g2_dlygate4sd3_1
XFILLER_29_636 VPWR VGND sg13g2_decap_8
XFILLER_28_157 VPWR VGND sg13g2_fill_1
X_4129_ net796 VGND VPWR _0107_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\]
+ clknet_5_31__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_43_105 VPWR VGND sg13g2_fill_1
XFILLER_25_842 VPWR VGND sg13g2_decap_8
XFILLER_40_823 VPWR VGND sg13g2_decap_8
XFILLER_12_525 VPWR VGND sg13g2_decap_8
XFILLER_4_768 VPWR VGND sg13g2_decap_8
XFILLER_0_974 VPWR VGND sg13g2_decap_8
XFILLER_48_934 VPWR VGND sg13g2_decap_8
XFILLER_47_444 VPWR VGND sg13g2_decap_8
XFILLER_35_639 VPWR VGND sg13g2_decap_8
XFILLER_28_680 VPWR VGND sg13g2_decap_8
XFILLER_16_886 VPWR VGND sg13g2_decap_8
XFILLER_37_1003 VPWR VGND sg13g2_decap_8
XFILLER_31_834 VPWR VGND sg13g2_decap_8
XFILLER_30_377 VPWR VGND sg13g2_decap_4
X_3500_ net585 VPWR _1029_ VGND net612 _1028_ sg13g2_o21ai_1
XFILLER_7_573 VPWR VGND sg13g2_decap_8
X_3431_ _0962_ net643 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] net651
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] VPWR VGND sg13g2_a22oi_1
X_3362_ _0894_ VPWR _0896_ VGND net560 _0873_ sg13g2_o21ai_1
XFILLER_44_1018 VPWR VGND sg13g2_decap_8
X_2313_ _1685_ _1726_ _1731_ _1733_ _1734_ VPWR VGND sg13g2_and4_1
X_3293_ net660 _0633_ _0829_ VPWR VGND sg13g2_nor2_1
XFILLER_39_901 VPWR VGND sg13g2_decap_8
X_2244_ _1665_ net696 _1553_ VPWR VGND sg13g2_nand2_1
X_2175_ net738 _1519_ _1562_ _1596_ VGND VPWR _1595_ sg13g2_nor4_2
XFILLER_18_0 VPWR VGND sg13g2_fill_1
XFILLER_39_978 VPWR VGND sg13g2_decap_8
XFILLER_26_639 VPWR VGND sg13g2_decap_8
XFILLER_19_691 VPWR VGND sg13g2_decap_8
XFILLER_22_834 VPWR VGND sg13g2_decap_8
XFILLER_34_683 VPWR VGND sg13g2_decap_8
XFILLER_21_355 VPWR VGND sg13g2_fill_1
X_3629_ net550 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] _1135_ _0096_
+ VPWR VGND sg13g2_a21o_1
Xoutput27 net27 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_716 VPWR VGND sg13g2_decap_8
Xoutput16 net16 uio_oe[7] VPWR VGND sg13g2_buf_1
XFILLER_45_926 VPWR VGND sg13g2_decap_8
XFILLER_16_127 VPWR VGND sg13g2_fill_1
XFILLER_16_138 VPWR VGND sg13g2_fill_2
XFILLER_44_458 VPWR VGND sg13g2_decap_8
XFILLER_32_609 VPWR VGND sg13g2_decap_8
XFILLER_40_620 VPWR VGND sg13g2_decap_8
XFILLER_13_845 VPWR VGND sg13g2_decap_8
XFILLER_40_697 VPWR VGND sg13g2_decap_8
XFILLER_9_838 VPWR VGND sg13g2_decap_8
XFILLER_12_366 VPWR VGND sg13g2_fill_2
XFILLER_4_565 VPWR VGND sg13g2_decap_8
XFILLER_0_771 VPWR VGND sg13g2_decap_8
XFILLER_48_731 VPWR VGND sg13g2_decap_8
XFILLER_36_948 VPWR VGND sg13g2_decap_8
X_3980_ _1401_ VPWR _0181_ VGND net548 _1400_ sg13g2_o21ai_1
X_2931_ _0495_ _0493_ _0324_ _0489_ _0488_ VPWR VGND sg13g2_a22oi_1
XFILLER_16_683 VPWR VGND sg13g2_decap_8
XFILLER_22_108 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_30_130 VPWR VGND sg13g2_fill_1
XFILLER_31_631 VPWR VGND sg13g2_decap_8
X_2862_ _0426_ _0427_ _0324_ _0428_ VPWR VGND sg13g2_nand3_1
X_2793_ _2008_ VPWR _0361_ VGND _0359_ _0360_ sg13g2_o21ai_1
XFILLER_8_860 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
X_3414_ _0946_ _0931_ _0945_ VPWR VGND sg13g2_xnor2_1
X_3345_ _0880_ _0820_ _0844_ VPWR VGND sg13g2_nand2_1
X_3276_ _0657_ _0670_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] _0812_
+ VPWR VGND _0710_ sg13g2_nand4_1
X_2227_ _1648_ _1578_ _1647_ VPWR VGND sg13g2_nand2_1
Xclkbuf_4_0_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_0_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_39_775 VPWR VGND sg13g2_decap_8
X_2158_ _1579_ _1533_ net710 _1527_ _1499_ VPWR VGND sg13g2_a22oi_1
XFILLER_26_436 VPWR VGND sg13g2_decap_8
X_2089_ net725 net727 _1510_ VPWR VGND sg13g2_nor2b_2
XFILLER_22_631 VPWR VGND sg13g2_decap_8
XFILLER_42_48 VPWR VGND sg13g2_fill_2
XFILLER_10_804 VPWR VGND sg13g2_decap_8
XFILLER_1_513 VPWR VGND sg13g2_decap_8
XFILLER_49_528 VPWR VGND sg13g2_decap_8
XFILLER_18_915 VPWR VGND sg13g2_decap_8
XFILLER_45_723 VPWR VGND sg13g2_decap_8
XFILLER_33_907 VPWR VGND sg13g2_decap_8
XFILLER_41_962 VPWR VGND sg13g2_decap_8
XFILLER_13_642 VPWR VGND sg13g2_decap_8
XFILLER_8_101 VPWR VGND sg13g2_decap_8
XFILLER_9_635 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_494 VPWR VGND sg13g2_decap_8
XFILLER_5_852 VPWR VGND sg13g2_decap_8
X_3130_ _1587_ _1592_ _1605_ _0666_ VPWR VGND sg13g2_nor3_1
X_3061_ VGND VPWR _1439_ net692 _0066_ _0597_ sg13g2_a21oi_1
X_2012_ VPWR _1435_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\] VGND sg13g2_inv_1
XFILLER_36_745 VPWR VGND sg13g2_decap_8
XFILLER_24_918 VPWR VGND sg13g2_decap_8
XFILLER_23_417 VPWR VGND sg13g2_decap_8
X_3963_ net602 _1025_ _1075_ _1389_ VPWR VGND sg13g2_nor3_1
X_2914_ VGND VPWR _0478_ sap_3_inst.alu.tmp\[5\] net747 sg13g2_or2_1
X_3894_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] _1333_
+ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] _1334_ _1306_ sg13g2_a221oi_1
XFILLER_32_973 VPWR VGND sg13g2_decap_8
X_2845_ net754 net672 _0411_ VPWR VGND sg13g2_nor2_1
X_2776_ _0345_ net720 _0321_ VPWR VGND sg13g2_nand2_1
Xfanout603 _0722_ net603 VPWR VGND sg13g2_buf_8
Xfanout614 net615 net614 VPWR VGND sg13g2_buf_8
Xfanout658 _0723_ net658 VPWR VGND sg13g2_buf_8
X_3328_ _1457_ _0717_ _0863_ VPWR VGND sg13g2_nor2_1
Xfanout647 net648 net647 VPWR VGND sg13g2_buf_1
Xfanout625 net626 net625 VPWR VGND sg13g2_buf_8
Xfanout636 _1795_ net636 VPWR VGND sg13g2_buf_8
Xfanout669 net670 net669 VPWR VGND sg13g2_buf_8
X_3259_ _0795_ _0789_ _0790_ _0791_ VPWR VGND sg13g2_and3_1
XFILLER_2_1015 VPWR VGND sg13g2_decap_8
XFILLER_39_572 VPWR VGND sg13g2_decap_8
XFILLER_27_767 VPWR VGND sg13g2_decap_8
XFILLER_42_748 VPWR VGND sg13g2_decap_8
XFILLER_10_601 VPWR VGND sg13g2_decap_8
XFILLER_23_962 VPWR VGND sg13g2_decap_8
XFILLER_10_678 VPWR VGND sg13g2_decap_8
XFILLER_6_638 VPWR VGND sg13g2_decap_8
XFILLER_5_126 VPWR VGND sg13g2_fill_1
XFILLER_5_159 VPWR VGND sg13g2_fill_1
XFILLER_2_833 VPWR VGND sg13g2_decap_8
XFILLER_49_325 VPWR VGND sg13g2_decap_8
XFILLER_45_520 VPWR VGND sg13g2_decap_8
XFILLER_17_200 VPWR VGND sg13g2_fill_1
XFILLER_18_712 VPWR VGND sg13g2_decap_8
XFILLER_17_222 VPWR VGND sg13g2_fill_2
XFILLER_17_244 VPWR VGND sg13g2_fill_2
XFILLER_27_81 VPWR VGND sg13g2_fill_1
XFILLER_33_704 VPWR VGND sg13g2_decap_8
XFILLER_45_597 VPWR VGND sg13g2_decap_8
XFILLER_18_789 VPWR VGND sg13g2_decap_8
XFILLER_40_291 VPWR VGND sg13g2_fill_1
X_2630_ sap_3_inst.alu.carry net675 _0226_ VPWR VGND sg13g2_nor2_1
X_2561_ VGND VPWR _1723_ _1963_ _1974_ _1973_ sg13g2_a21oi_1
X_2492_ _1907_ _1904_ _1905_ _1906_ VPWR VGND sg13g2_and3_1
X_4162_ net786 VGND VPWR _0140_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3113_ _0642_ _0646_ _0647_ _0648_ _0649_ VPWR VGND sg13g2_and4_1
X_4093_ net774 VGND VPWR _0071_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[4\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
XFILLER_49_892 VPWR VGND sg13g2_decap_8
X_3044_ _0590_ sap_3_inst.alu.tmp\[6\] net668 VPWR VGND sg13g2_nand2_1
XFILLER_36_542 VPWR VGND sg13g2_decap_8
XFILLER_24_715 VPWR VGND sg13g2_decap_8
X_3946_ _1380_ _1311_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] _1302_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_32_770 VPWR VGND sg13g2_decap_8
XFILLER_23_39 VPWR VGND sg13g2_fill_2
XFILLER_20_954 VPWR VGND sg13g2_decap_8
X_3877_ _1318_ _1308_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] _1305_
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2828_ _0394_ VPWR _0395_ VGND net755 _0327_ sg13g2_o21ai_1
XFILLER_3_619 VPWR VGND sg13g2_decap_8
X_2759_ VGND VPWR _0202_ _0316_ _0328_ _1936_ sg13g2_a21oi_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_24_1016 VPWR VGND sg13g2_decap_8
XFILLER_24_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_829 VPWR VGND sg13g2_decap_8
XFILLER_19_509 VPWR VGND sg13g2_decap_8
XFILLER_27_564 VPWR VGND sg13g2_decap_8
XFILLER_42_545 VPWR VGND sg13g2_decap_8
XFILLER_15_759 VPWR VGND sg13g2_decap_8
XFILLER_11_921 VPWR VGND sg13g2_decap_8
XFILLER_31_1009 VPWR VGND sg13g2_decap_8
XFILLER_7_958 VPWR VGND sg13g2_decap_8
XFILLER_11_998 VPWR VGND sg13g2_decap_8
XFILLER_2_630 VPWR VGND sg13g2_decap_8
XFILLER_18_586 VPWR VGND sg13g2_decap_8
XFILLER_33_501 VPWR VGND sg13g2_decap_8
XFILLER_45_394 VPWR VGND sg13g2_decap_8
X_3800_ net598 _1033_ _1195_ _1257_ VPWR VGND sg13g2_nor3_1
XFILLER_33_578 VPWR VGND sg13g2_decap_8
X_3731_ net556 _1211_ VPWR VGND sg13g2_inv_4
XFILLER_13_291 VPWR VGND sg13g2_fill_2
X_3662_ _1161_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] net596 VPWR
+ VGND sg13g2_nand2_1
Xclkload10 VPWR clkload10/Y clknet_5_5__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_2613_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] net636
+ _0210_ net637 sg13g2_a21oi_1
X_3593_ _1108_ _0844_ _0854_ VPWR VGND sg13g2_nand2_1
X_2544_ _1957_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] net634
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_2475_ _1890_ _1891_ _1892_ VPWR VGND sg13g2_and2_1
X_4214_ net797 VGND VPWR _0191_ sap_3_inst.reg_file.array_serializer_inst.word_index\[1\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_2
XFILLER_29_818 VPWR VGND sg13g2_decap_8
X_4145_ net796 VGND VPWR _0123_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\]
+ clknet_5_29__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4076_ net789 VGND VPWR _0054_ sap_3_inst.alu.tmp\[3\] clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3027_ _0568_ VPWR _0580_ VGND _0323_ _0565_ sg13g2_o21ai_1
XFILLER_24_512 VPWR VGND sg13g2_decap_8
XFILLER_37_884 VPWR VGND sg13g2_decap_8
XFILLER_12_707 VPWR VGND sg13g2_decap_8
XFILLER_24_589 VPWR VGND sg13g2_decap_8
X_3929_ _1362_ _1363_ _1361_ _1365_ VPWR VGND _1364_ sg13g2_nand4_1
XFILLER_20_751 VPWR VGND sg13g2_decap_8
Xclkload4 VPWR clkload4/Y clknet_3_5__leaf_clk VGND sg13g2_inv_1
XFILLER_8_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_626 VPWR VGND sg13g2_decap_8
XFILLER_43_810 VPWR VGND sg13g2_decap_8
XFILLER_28_862 VPWR VGND sg13g2_decap_8
XFILLER_43_887 VPWR VGND sg13g2_decap_8
XFILLER_15_556 VPWR VGND sg13g2_decap_8
XFILLER_10_261 VPWR VGND sg13g2_fill_2
XFILLER_7_755 VPWR VGND sg13g2_decap_8
XFILLER_11_795 VPWR VGND sg13g2_decap_8
XFILLER_3_983 VPWR VGND sg13g2_decap_8
X_2260_ _1648_ VPWR _1681_ VGND _1592_ _1679_ sg13g2_o21ai_1
X_2191_ VGND VPWR _1612_ _1595_ _1524_ sg13g2_or2_1
XFILLER_37_125 VPWR VGND sg13g2_fill_1
XFILLER_38_648 VPWR VGND sg13g2_decap_8
XFILLER_19_873 VPWR VGND sg13g2_decap_8
XFILLER_34_865 VPWR VGND sg13g2_decap_8
Xclkbuf_5_5__f_sap_3_inst.alu.clk_regs clknet_4_2_0_sap_3_inst.alu.clk_regs clknet_5_5__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_21_548 VPWR VGND sg13g2_decap_8
X_3714_ _1199_ _0850_ _1048_ _1200_ VPWR VGND sg13g2_a21o_1
X_3645_ net11 net19 _0836_ _1147_ VPWR VGND sg13g2_mux2_1
X_3576_ _0085_ _1092_ _1093_ net589 _1453_ VPWR VGND sg13g2_a22oi_1
X_2527_ _1940_ _1939_ VPWR VGND sg13g2_inv_2
X_2458_ _1868_ VPWR _1877_ VGND net565 _1876_ sg13g2_o21ai_1
Xhold27 u_ser.shadow_reg\[4\] VPWR VGND net74 sg13g2_dlygate4sd3_1
Xhold16 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\] VPWR VGND net63 sg13g2_dlygate4sd3_1
X_2389_ _1810_ _1804_ _1809_ net638 _1490_ VPWR VGND sg13g2_a22oi_1
XFILLER_29_615 VPWR VGND sg13g2_decap_8
X_4128_ net775 VGND VPWR _0106_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\]
+ clknet_5_3__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4059_ net789 VGND VPWR _0037_ sap_3_inst.alu.acc\[3\] clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_43_128 VPWR VGND sg13g2_fill_2
XFILLER_25_821 VPWR VGND sg13g2_decap_8
XFILLER_37_681 VPWR VGND sg13g2_decap_8
XFILLER_40_802 VPWR VGND sg13g2_decap_8
XFILLER_12_504 VPWR VGND sg13g2_decap_8
XFILLER_24_386 VPWR VGND sg13g2_decap_8
XFILLER_25_898 VPWR VGND sg13g2_decap_8
XFILLER_40_879 VPWR VGND sg13g2_decap_8
XFILLER_4_747 VPWR VGND sg13g2_decap_8
XFILLER_48_913 VPWR VGND sg13g2_decap_8
XFILLER_0_953 VPWR VGND sg13g2_decap_8
XFILLER_47_423 VPWR VGND sg13g2_decap_8
XFILLER_35_618 VPWR VGND sg13g2_decap_8
XFILLER_34_117 VPWR VGND sg13g2_fill_1
XFILLER_16_865 VPWR VGND sg13g2_decap_8
XFILLER_43_684 VPWR VGND sg13g2_decap_8
XFILLER_31_813 VPWR VGND sg13g2_decap_8
Xclkbuf_5_12__f_sap_3_inst.alu.clk_regs clknet_4_6_0_sap_3_inst.alu.clk_regs clknet_5_12__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_11_592 VPWR VGND sg13g2_decap_8
XFILLER_7_552 VPWR VGND sg13g2_decap_8
X_3430_ _0961_ net655 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] net606
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] VPWR VGND sg13g2_a22oi_1
X_3361_ VPWR _0895_ _0894_ VGND sg13g2_inv_1
X_2312_ _1660_ _1732_ _1733_ VPWR VGND sg13g2_nor2_1
XFILLER_3_780 VPWR VGND sg13g2_decap_8
X_3292_ _0828_ _0744_ _0826_ VPWR VGND sg13g2_xnor2_1
X_2243_ net694 _1554_ _1664_ VPWR VGND sg13g2_nor2_1
X_2174_ net741 net736 _1595_ VPWR VGND net739 sg13g2_nand3b_1
XFILLER_39_957 VPWR VGND sg13g2_decap_8
XFILLER_26_618 VPWR VGND sg13g2_decap_8
XFILLER_47_990 VPWR VGND sg13g2_decap_8
XFILLER_19_670 VPWR VGND sg13g2_decap_8
XFILLER_34_662 VPWR VGND sg13g2_decap_8
XFILLER_22_813 VPWR VGND sg13g2_decap_8
X_3628_ net550 _1133_ _1134_ _1135_ VPWR VGND sg13g2_nor3_1
Xoutput28 net28 uo_out[3] VPWR VGND sg13g2_buf_1
Xoutput17 net31 uio_out[0] VPWR VGND sg13g2_buf_1
X_3559_ _1079_ net31 _1077_ VPWR VGND sg13g2_nand2_1
XFILLER_5_1013 VPWR VGND sg13g2_decap_8
XFILLER_45_905 VPWR VGND sg13g2_decap_8
XFILLER_29_489 VPWR VGND sg13g2_decap_8
XFILLER_44_437 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_sap_3_inst.alu.clk clknet_0_sap_3_inst.alu.clk clknet_1_1__leaf_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_13_824 VPWR VGND sg13g2_decap_8
XFILLER_25_695 VPWR VGND sg13g2_decap_8
XFILLER_9_817 VPWR VGND sg13g2_decap_8
XFILLER_40_676 VPWR VGND sg13g2_decap_8
XFILLER_4_544 VPWR VGND sg13g2_decap_8
XFILLER_0_750 VPWR VGND sg13g2_decap_8
XFILLER_48_710 VPWR VGND sg13g2_decap_8
XFILLER_48_787 VPWR VGND sg13g2_decap_8
XFILLER_36_927 VPWR VGND sg13g2_decap_8
XFILLER_35_459 VPWR VGND sg13g2_fill_1
X_2930_ net544 _0481_ _0484_ _0494_ VPWR VGND sg13g2_nor3_1
XFILLER_16_662 VPWR VGND sg13g2_decap_8
XFILLER_31_610 VPWR VGND sg13g2_decap_8
XFILLER_43_481 VPWR VGND sg13g2_decap_8
X_2861_ _0425_ VPWR _0427_ VGND _0366_ _0387_ sg13g2_o21ai_1
XFILLER_31_687 VPWR VGND sg13g2_decap_8
X_2792_ _0343_ _0358_ _0360_ VPWR VGND sg13g2_and2_1
XFILLER_7_41 VPWR VGND sg13g2_fill_1
X_3413_ VPWR _0945_ net552 VGND sg13g2_inv_1
X_3344_ _0878_ VPWR _0879_ VGND net32 _0838_ sg13g2_o21ai_1
XFILLER_30_0 VPWR VGND sg13g2_fill_2
X_3275_ _0658_ net665 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] _0811_
+ VPWR VGND _0710_ sg13g2_nand4_1
X_2226_ _1647_ net714 net705 VPWR VGND sg13g2_nand2_2
XFILLER_39_754 VPWR VGND sg13g2_decap_8
X_2157_ _1578_ _1533_ net710 VPWR VGND sg13g2_nand2_2
XFILLER_26_415 VPWR VGND sg13g2_decap_8
XFILLER_27_949 VPWR VGND sg13g2_decap_8
X_2088_ net737 net740 _1509_ VPWR VGND net742 sg13g2_nand3b_1
XFILLER_41_418 VPWR VGND sg13g2_decap_4
XFILLER_22_610 VPWR VGND sg13g2_decap_8
XFILLER_35_982 VPWR VGND sg13g2_decap_8
XFILLER_42_38 VPWR VGND sg13g2_fill_2
XFILLER_22_687 VPWR VGND sg13g2_decap_8
XFILLER_1_569 VPWR VGND sg13g2_decap_8
XFILLER_49_507 VPWR VGND sg13g2_decap_8
XFILLER_45_702 VPWR VGND sg13g2_decap_8
XFILLER_45_779 VPWR VGND sg13g2_decap_8
XFILLER_26_982 VPWR VGND sg13g2_decap_8
XFILLER_41_941 VPWR VGND sg13g2_decap_8
XFILLER_13_621 VPWR VGND sg13g2_decap_8
XFILLER_25_492 VPWR VGND sg13g2_decap_8
XFILLER_9_614 VPWR VGND sg13g2_decap_8
XFILLER_40_473 VPWR VGND sg13g2_decap_8
XFILLER_13_698 VPWR VGND sg13g2_decap_8
XFILLER_5_831 VPWR VGND sg13g2_decap_8
X_3060_ net692 net24 _0597_ VPWR VGND sg13g2_nor2_1
X_2011_ VPWR _1434_ u_ser.bit_pos\[2\] VGND sg13g2_inv_1
XFILLER_48_584 VPWR VGND sg13g2_decap_8
XFILLER_36_724 VPWR VGND sg13g2_decap_8
XFILLER_35_245 VPWR VGND sg13g2_fill_2
XFILLER_23_407 VPWR VGND sg13g2_decap_4
XFILLER_32_952 VPWR VGND sg13g2_decap_8
X_3962_ VGND VPWR _1480_ net605 _0176_ _1388_ sg13g2_a21oi_1
X_2913_ net747 sap_3_inst.alu.tmp\[5\] _0477_ VPWR VGND sg13g2_and2_1
X_3893_ _1330_ _1331_ _1329_ _1333_ VPWR VGND _1332_ sg13g2_nand4_1
X_2844_ _0410_ _0399_ _0403_ VPWR VGND sg13g2_nand2_1
XFILLER_31_484 VPWR VGND sg13g2_decap_8
X_2775_ _0344_ _0321_ net720 VPWR VGND sg13g2_nand2b_1
Xfanout615 _0714_ net615 VPWR VGND sg13g2_buf_8
Xfanout604 _0722_ net604 VPWR VGND sg13g2_buf_8
Xfanout648 _0732_ net648 VPWR VGND sg13g2_buf_8
Xfanout637 _1794_ net637 VPWR VGND sg13g2_buf_8
Xfanout626 _1800_ net626 VPWR VGND sg13g2_buf_8
X_3327_ _0718_ VPWR _0067_ VGND _0848_ _0862_ sg13g2_o21ai_1
Xfanout659 _0712_ net659 VPWR VGND sg13g2_buf_8
X_3258_ _0794_ net657 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] net609
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_551 VPWR VGND sg13g2_decap_8
X_2209_ VGND VPWR _1579_ _1627_ _1630_ _1597_ sg13g2_a21oi_1
X_3189_ _0725_ net657 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] net609
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_27_746 VPWR VGND sg13g2_decap_8
XFILLER_42_727 VPWR VGND sg13g2_decap_8
XFILLER_14_407 VPWR VGND sg13g2_fill_1
XFILLER_23_941 VPWR VGND sg13g2_decap_8
XFILLER_22_484 VPWR VGND sg13g2_decap_8
XFILLER_6_617 VPWR VGND sg13g2_decap_8
XFILLER_10_657 VPWR VGND sg13g2_decap_8
XFILLER_5_149 VPWR VGND sg13g2_fill_2
XFILLER_2_812 VPWR VGND sg13g2_decap_8
XFILLER_2_889 VPWR VGND sg13g2_decap_8
XFILLER_18_768 VPWR VGND sg13g2_decap_8
XFILLER_45_576 VPWR VGND sg13g2_decap_8
XFILLER_14_985 VPWR VGND sg13g2_decap_8
XFILLER_32_259 VPWR VGND sg13g2_fill_2
XFILLER_9_488 VPWR VGND sg13g2_decap_8
X_2560_ VGND VPWR _1968_ _1972_ _1973_ net566 sg13g2_a21oi_1
X_2491_ _1906_ net625 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] net677
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4161_ net796 VGND VPWR _0139_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\]
+ clknet_5_26__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3112_ _1730_ _0636_ _0637_ _0643_ _0648_ VPWR VGND sg13g2_and4_1
X_4092_ net782 VGND VPWR _0070_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[3\]
+ clknet_5_6__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
XFILLER_49_871 VPWR VGND sg13g2_decap_8
X_3043_ _0589_ VPWR _0056_ VGND _1899_ net667 sg13g2_o21ai_1
XFILLER_36_521 VPWR VGND sg13g2_decap_8
XFILLER_48_381 VPWR VGND sg13g2_decap_8
XFILLER_36_598 VPWR VGND sg13g2_decap_8
X_3945_ _1379_ _1313_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] _1305_
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_933 VPWR VGND sg13g2_decap_8
X_3876_ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\] net768 _1300_ _1317_
+ VPWR VGND sg13g2_nor3_2
XFILLER_31_281 VPWR VGND sg13g2_fill_1
X_2827_ net563 VPWR _0394_ VGND net755 sap_3_inst.alu.tmp\[2\] sg13g2_o21ai_1
X_2758_ _0327_ _0202_ _0316_ VPWR VGND sg13g2_nand2_2
X_2689_ _1526_ _0279_ _0280_ _0281_ VPWR VGND sg13g2_nor3_1
XFILLER_47_808 VPWR VGND sg13g2_decap_8
XFILLER_27_543 VPWR VGND sg13g2_decap_8
XFILLER_42_524 VPWR VGND sg13g2_decap_8
XFILLER_15_738 VPWR VGND sg13g2_decap_8
XFILLER_11_900 VPWR VGND sg13g2_decap_8
XFILLER_14_248 VPWR VGND sg13g2_fill_1
XFILLER_11_977 VPWR VGND sg13g2_decap_8
XFILLER_7_937 VPWR VGND sg13g2_decap_8
XFILLER_2_686 VPWR VGND sg13g2_decap_8
XFILLER_1_185 VPWR VGND sg13g2_fill_2
XFILLER_46_885 VPWR VGND sg13g2_decap_8
XFILLER_18_565 VPWR VGND sg13g2_decap_8
XFILLER_45_373 VPWR VGND sg13g2_decap_8
XFILLER_33_557 VPWR VGND sg13g2_decap_8
XFILLER_14_782 VPWR VGND sg13g2_decap_8
X_3730_ net650 _1209_ _1210_ VPWR VGND sg13g2_nor2_2
X_3661_ _0103_ _1102_ _1160_ net596 _1473_ VPWR VGND sg13g2_a22oi_1
X_3592_ VGND VPWR _1899_ net570 _1107_ _1106_ sg13g2_a21oi_1
X_2612_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] _0206_
+ net626 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] _0209_ net630 sg13g2_a221oi_1
Xclkload11 clknet_5_6__leaf_sap_3_inst.alu.clk_regs clkload11/X VPWR VGND sg13g2_buf_1
XFILLER_6_981 VPWR VGND sg13g2_decap_8
X_2543_ _1956_ net622 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] net636
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2474_ _1891_ net623 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] net638
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4213_ net797 VGND VPWR _0190_ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_2
X_4144_ net777 VGND VPWR _0122_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\]
+ clknet_5_11__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4075_ net789 VGND VPWR _0053_ sap_3_inst.alu.tmp\[2\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3026_ _0577_ _0578_ _0575_ _0579_ VPWR VGND sg13g2_nand3_1
XFILLER_37_863 VPWR VGND sg13g2_decap_8
XFILLER_24_568 VPWR VGND sg13g2_decap_8
X_3928_ _1364_ _1305_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] _1302_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_730 VPWR VGND sg13g2_decap_8
Xclkload5 VPWR clkload5/Y clknet_3_6__leaf_clk VGND sg13g2_inv_1
X_3859_ _1300_ sap_3_inst.reg_file.array_serializer_inst.word_index\[3\] VPWR VGND
+ sap_3_inst.reg_file.array_serializer_inst.word_index\[2\] sg13g2_nand2b_2
XFILLER_4_929 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_fill_2
XFILLER_8_1000 VPWR VGND sg13g2_decap_8
XFILLER_47_605 VPWR VGND sg13g2_decap_8
XFILLER_46_137 VPWR VGND sg13g2_fill_1
XFILLER_28_841 VPWR VGND sg13g2_decap_8
XFILLER_15_535 VPWR VGND sg13g2_decap_8
XFILLER_43_866 VPWR VGND sg13g2_decap_8
XFILLER_30_549 VPWR VGND sg13g2_decap_8
XFILLER_7_734 VPWR VGND sg13g2_decap_8
XFILLER_11_774 VPWR VGND sg13g2_decap_8
XFILLER_3_962 VPWR VGND sg13g2_decap_8
XFILLER_2_483 VPWR VGND sg13g2_decap_8
X_2190_ net722 _1595_ _1611_ VPWR VGND sg13g2_nor2_1
XFILLER_38_627 VPWR VGND sg13g2_decap_8
XFILLER_1_54 VPWR VGND sg13g2_decap_4
XFILLER_1_43 VPWR VGND sg13g2_fill_1
XFILLER_19_852 VPWR VGND sg13g2_decap_8
XFILLER_18_340 VPWR VGND sg13g2_fill_2
XFILLER_46_682 VPWR VGND sg13g2_decap_8
XFILLER_34_844 VPWR VGND sg13g2_decap_8
XFILLER_21_527 VPWR VGND sg13g2_decap_8
XFILLER_14_1027 VPWR VGND sg13g2_fill_2
X_3713_ VGND VPWR _0808_ _0820_ _1199_ _0845_ sg13g2_a21oi_1
X_3644_ VGND VPWR _1459_ net596 _0100_ _1146_ sg13g2_a21oi_1
X_3575_ VGND VPWR net577 _0898_ _1093_ net589 sg13g2_a21oi_1
X_2526_ _1858_ VPWR _1939_ VGND _1922_ _1935_ sg13g2_o21ai_1
X_2457_ _1871_ _1875_ _1876_ VPWR VGND sg13g2_nor2_1
Xhold28 sap_3_inst.reg_file.array_serializer_inst.state\[1\] VPWR VGND net75 sg13g2_dlygate4sd3_1
Xhold17 _0159_ VPWR VGND net64 sg13g2_dlygate4sd3_1
X_2388_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] _1808_
+ net621 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] _1809_ net631 sg13g2_a221oi_1
X_4127_ net780 VGND VPWR _0105_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_44_619 VPWR VGND sg13g2_decap_8
X_4058_ net790 VGND VPWR _0036_ sap_3_inst.alu.acc\[2\] clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_25_800 VPWR VGND sg13g2_decap_8
XFILLER_37_660 VPWR VGND sg13g2_decap_8
X_3009_ _0562_ _1938_ _0204_ VPWR VGND sg13g2_nand2b_1
XFILLER_25_877 VPWR VGND sg13g2_decap_8
XFILLER_40_858 VPWR VGND sg13g2_decap_8
XFILLER_4_726 VPWR VGND sg13g2_decap_8
XFILLER_0_932 VPWR VGND sg13g2_decap_8
XFILLER_47_402 VPWR VGND sg13g2_decap_8
XFILLER_48_969 VPWR VGND sg13g2_decap_8
XFILLER_47_479 VPWR VGND sg13g2_decap_8
XFILLER_16_844 VPWR VGND sg13g2_decap_8
XFILLER_43_663 VPWR VGND sg13g2_decap_8
XFILLER_27_192 VPWR VGND sg13g2_fill_2
XFILLER_31_869 VPWR VGND sg13g2_decap_8
XFILLER_7_531 VPWR VGND sg13g2_decap_8
XFILLER_11_571 VPWR VGND sg13g2_decap_8
X_3360_ _0893_ VPWR _0894_ VGND sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[2\]
+ net610 sg13g2_o21ai_1
X_2311_ VGND VPWR _1604_ _1606_ _1732_ _1642_ sg13g2_a21oi_1
X_3291_ net553 _0825_ _0744_ _0827_ VPWR VGND sg13g2_nand3_1
X_2242_ VGND VPWR _1579_ _1627_ _1663_ _1662_ sg13g2_a21oi_1
XFILLER_39_936 VPWR VGND sg13g2_decap_8
X_2173_ _1590_ _1593_ _1588_ _1594_ VPWR VGND sg13g2_nand3_1
XFILLER_38_468 VPWR VGND sg13g2_fill_2
XFILLER_34_641 VPWR VGND sg13g2_decap_8
XFILLER_21_313 VPWR VGND sg13g2_fill_1
XFILLER_21_324 VPWR VGND sg13g2_fill_1
XFILLER_22_869 VPWR VGND sg13g2_decap_8
X_3627_ net579 _0987_ _1134_ VPWR VGND sg13g2_and2_1
Xoutput18 net32 uio_out[1] VPWR VGND sg13g2_buf_1
Xoutput29 net29 uo_out[4] VPWR VGND sg13g2_buf_1
X_3558_ net570 _1078_ VPWR VGND sg13g2_inv_4
X_2509_ VGND VPWR _1540_ net688 _1922_ net682 sg13g2_a21oi_1
X_3489_ _1018_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] net640 VPWR
+ VGND sg13g2_nand2_1
XFILLER_17_619 VPWR VGND sg13g2_decap_8
XFILLER_29_468 VPWR VGND sg13g2_decap_8
XFILLER_44_416 VPWR VGND sg13g2_decap_8
XFILLER_38_991 VPWR VGND sg13g2_decap_8
XFILLER_13_803 VPWR VGND sg13g2_decap_8
XFILLER_25_674 VPWR VGND sg13g2_decap_8
XFILLER_40_655 VPWR VGND sg13g2_decap_8
XFILLER_21_891 VPWR VGND sg13g2_decap_8
XFILLER_4_523 VPWR VGND sg13g2_decap_8
XFILLER_43_1020 VPWR VGND sg13g2_decap_8
XFILLER_48_766 VPWR VGND sg13g2_decap_8
XFILLER_36_906 VPWR VGND sg13g2_decap_8
XFILLER_16_641 VPWR VGND sg13g2_decap_8
XFILLER_44_983 VPWR VGND sg13g2_decap_8
XFILLER_43_460 VPWR VGND sg13g2_decap_8
X_2860_ _0366_ _0387_ _0425_ _0426_ VPWR VGND sg13g2_or3_1
XFILLER_31_666 VPWR VGND sg13g2_decap_8
X_2791_ _0343_ _0358_ _0359_ VPWR VGND sg13g2_nor2_1
XFILLER_7_53 VPWR VGND sg13g2_decap_8
XFILLER_11_1019 VPWR VGND sg13g2_decap_8
XFILLER_8_895 VPWR VGND sg13g2_decap_8
X_3412_ _0943_ VPWR _0944_ VGND _0940_ _0942_ sg13g2_o21ai_1
X_3343_ _0878_ _0838_ net10 VPWR VGND sg13g2_nand2b_1
X_3274_ _0710_ _0728_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] _0810_
+ VPWR VGND sg13g2_nand3_1
X_2225_ net714 net704 _1646_ VPWR VGND sg13g2_and2_1
XFILLER_39_733 VPWR VGND sg13g2_decap_8
XFILLER_27_928 VPWR VGND sg13g2_decap_8
X_2156_ _1533_ _1556_ _1577_ VPWR VGND sg13g2_and2_1
XFILLER_26_29 VPWR VGND sg13g2_fill_2
XFILLER_42_909 VPWR VGND sg13g2_decap_8
X_2087_ _1436_ _1507_ _1508_ VPWR VGND sg13g2_nor2_2
XFILLER_35_961 VPWR VGND sg13g2_decap_8
XFILLER_34_460 VPWR VGND sg13g2_fill_2
XFILLER_34_471 VPWR VGND sg13g2_fill_1
XFILLER_21_132 VPWR VGND sg13g2_fill_1
XFILLER_22_666 VPWR VGND sg13g2_decap_8
XFILLER_10_839 VPWR VGND sg13g2_decap_8
X_2989_ _0506_ VPWR _0551_ VGND _0505_ _0515_ sg13g2_o21ai_1
XFILLER_1_548 VPWR VGND sg13g2_decap_8
XFILLER_27_1026 VPWR VGND sg13g2_fill_2
XFILLER_17_405 VPWR VGND sg13g2_fill_2
XFILLER_45_758 VPWR VGND sg13g2_decap_8
XFILLER_44_246 VPWR VGND sg13g2_fill_2
XFILLER_13_600 VPWR VGND sg13g2_decap_8
XFILLER_26_961 VPWR VGND sg13g2_decap_8
XFILLER_41_920 VPWR VGND sg13g2_decap_8
XFILLER_25_471 VPWR VGND sg13g2_decap_8
XFILLER_40_441 VPWR VGND sg13g2_fill_2
XFILLER_13_677 VPWR VGND sg13g2_decap_8
XFILLER_34_1019 VPWR VGND sg13g2_decap_8
XFILLER_41_997 VPWR VGND sg13g2_decap_8
XFILLER_5_810 VPWR VGND sg13g2_decap_8
XFILLER_5_887 VPWR VGND sg13g2_decap_8
XFILLER_48_563 VPWR VGND sg13g2_decap_8
X_2010_ VPWR _1433_ u_ser.state\[1\] VGND sg13g2_inv_1
XFILLER_36_703 VPWR VGND sg13g2_decap_8
XFILLER_17_983 VPWR VGND sg13g2_decap_8
X_3961_ net604 _1002_ _1068_ _1388_ VPWR VGND sg13g2_nor3_1
XFILLER_44_780 VPWR VGND sg13g2_decap_8
X_2912_ _0476_ _0339_ net746 _0338_ net752 VPWR VGND sg13g2_a22oi_1
XFILLER_32_931 VPWR VGND sg13g2_decap_8
X_3892_ _1332_ net761 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] _1302_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2843_ net554 sap_3_inst.alu.acc\[2\] _0409_ _0036_ VPWR VGND sg13g2_a21o_1
X_2774_ _0343_ net720 _0321_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_692 VPWR VGND sg13g2_decap_8
Xfanout605 _0722_ net605 VPWR VGND sg13g2_buf_1
Xfanout638 net639 net638 VPWR VGND sg13g2_buf_8
Xfanout616 net617 net616 VPWR VGND sg13g2_buf_8
X_3326_ _0717_ VPWR _0862_ VGND _0843_ _0860_ sg13g2_o21ai_1
Xfanout649 net650 net649 VPWR VGND sg13g2_buf_8
Xfanout627 net628 net627 VPWR VGND sg13g2_buf_8
X_3257_ _0793_ net588 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] net615
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_530 VPWR VGND sg13g2_decap_8
X_2208_ VGND VPWR _1623_ _1628_ _1629_ _1600_ sg13g2_a21oi_1
XFILLER_27_725 VPWR VGND sg13g2_decap_8
X_3188_ _0724_ _0672_ _0695_ VPWR VGND sg13g2_nand2_2
X_2139_ _1555_ VPWR _1560_ VGND net699 _1558_ sg13g2_o21ai_1
XFILLER_42_706 VPWR VGND sg13g2_decap_8
XFILLER_23_920 VPWR VGND sg13g2_decap_8
XFILLER_10_636 VPWR VGND sg13g2_decap_8
XFILLER_22_463 VPWR VGND sg13g2_decap_8
XFILLER_23_997 VPWR VGND sg13g2_decap_8
XFILLER_2_868 VPWR VGND sg13g2_decap_8
XFILLER_40_1012 VPWR VGND sg13g2_decap_8
XFILLER_45_555 VPWR VGND sg13g2_decap_8
XFILLER_18_747 VPWR VGND sg13g2_decap_8
XFILLER_33_739 VPWR VGND sg13g2_decap_8
XFILLER_14_964 VPWR VGND sg13g2_decap_8
XFILLER_41_794 VPWR VGND sg13g2_decap_8
X_2490_ _1905_ net627 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] net635
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_684 VPWR VGND sg13g2_decap_8
X_4160_ net775 VGND VPWR _0138_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\]
+ clknet_5_11__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3111_ _1715_ _1818_ _0603_ _0647_ VPWR VGND sg13g2_nor3_1
XFILLER_4_87 VPWR VGND sg13g2_decap_8
XFILLER_49_850 VPWR VGND sg13g2_decap_8
X_4091_ net774 VGND VPWR _0069_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[2\]
+ clknet_5_1__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_48_360 VPWR VGND sg13g2_decap_8
X_3042_ _0589_ sap_3_inst.alu.tmp\[5\] net667 VPWR VGND sg13g2_nand2_1
XFILLER_36_500 VPWR VGND sg13g2_decap_8
XFILLER_36_577 VPWR VGND sg13g2_decap_8
XFILLER_17_780 VPWR VGND sg13g2_decap_8
X_3944_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] _1317_
+ _1378_ net763 sg13g2_a21oi_1
X_3875_ _1303_ _1307_ _1316_ VPWR VGND sg13g2_nor2_2
XFILLER_17_1025 VPWR VGND sg13g2_decap_4
XFILLER_20_912 VPWR VGND sg13g2_decap_8
X_2826_ _0391_ _0359_ _0393_ VPWR VGND sg13g2_xor2_1
XFILLER_20_989 VPWR VGND sg13g2_decap_8
X_2757_ _0322_ _0324_ _0326_ VPWR VGND sg13g2_nor2_1
X_2688_ VGND VPWR net703 _1515_ _0280_ _1675_ sg13g2_a21oi_1
X_3309_ _0845_ net661 net666 VPWR VGND sg13g2_nand2_1
XFILLER_27_522 VPWR VGND sg13g2_decap_8
XFILLER_42_503 VPWR VGND sg13g2_decap_8
XFILLER_15_717 VPWR VGND sg13g2_decap_8
XFILLER_27_599 VPWR VGND sg13g2_decap_8
Xfanout31 net17 net31 VPWR VGND sg13g2_buf_2
XFILLER_23_794 VPWR VGND sg13g2_decap_8
XFILLER_7_916 VPWR VGND sg13g2_decap_8
XFILLER_11_956 VPWR VGND sg13g2_decap_8
XFILLER_2_665 VPWR VGND sg13g2_decap_8
XFILLER_38_809 VPWR VGND sg13g2_decap_8
XFILLER_18_544 VPWR VGND sg13g2_decap_8
XFILLER_46_864 VPWR VGND sg13g2_decap_8
XFILLER_33_536 VPWR VGND sg13g2_decap_8
XFILLER_21_709 VPWR VGND sg13g2_decap_8
XFILLER_14_761 VPWR VGND sg13g2_decap_8
XFILLER_41_591 VPWR VGND sg13g2_decap_8
XFILLER_9_220 VPWR VGND sg13g2_fill_1
XFILLER_13_271 VPWR VGND sg13g2_fill_2
XFILLER_13_293 VPWR VGND sg13g2_fill_1
X_3660_ net596 _1159_ _1160_ VPWR VGND sg13g2_nor2_1
Xclkload12 VPWR clkload12/Y clknet_5_9__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_3591_ net14 net570 _1106_ VPWR VGND sg13g2_nor2_1
X_2611_ _0208_ net620 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\] net622
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_960 VPWR VGND sg13g2_decap_8
X_2542_ VGND VPWR _1945_ _1953_ _1955_ _1940_ sg13g2_a21oi_1
XFILLER_47_1018 VPWR VGND sg13g2_decap_8
XFILLER_5_481 VPWR VGND sg13g2_decap_8
X_2473_ _1890_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] net635
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4212_ net783 VGND VPWR net69 sap_3_outputReg_start_sync clknet_3_0__leaf_clk sg13g2_dfrbpq_1
X_4143_ net780 VGND VPWR _0121_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4074_ net785 VGND VPWR _0052_ sap_3_inst.alu.tmp\[1\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3025_ _0578_ net572 net760 net573 net744 VPWR VGND sg13g2_a22oi_1
XFILLER_37_842 VPWR VGND sg13g2_decap_8
XFILLER_24_547 VPWR VGND sg13g2_decap_8
X_3927_ _1363_ _1313_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] _1311_
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_786 VPWR VGND sg13g2_decap_8
Xclkload6 VPWR clkload6/Y clknet_3_7__leaf_clk VGND sg13g2_inv_1
X_3858_ VGND VPWR _1298_ _1299_ _0161_ _1290_ sg13g2_a21oi_1
X_2809_ VGND VPWR net544 _0368_ _0377_ net670 sg13g2_a21oi_1
XFILLER_4_908 VPWR VGND sg13g2_decap_8
X_3789_ net600 _1050_ _1200_ _1251_ VPWR VGND sg13g2_nor3_1
XFILLER_30_1011 VPWR VGND sg13g2_decap_8
Xclkbuf_5_20__f_sap_3_inst.alu.clk_regs clknet_4_10_0_sap_3_inst.alu.clk_regs clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_46_127 VPWR VGND sg13g2_fill_1
XFILLER_28_820 VPWR VGND sg13g2_decap_8
XFILLER_43_845 VPWR VGND sg13g2_decap_8
XFILLER_15_514 VPWR VGND sg13g2_decap_8
XFILLER_28_897 VPWR VGND sg13g2_decap_8
XFILLER_30_528 VPWR VGND sg13g2_decap_8
XFILLER_23_591 VPWR VGND sg13g2_decap_8
XFILLER_7_713 VPWR VGND sg13g2_decap_8
XFILLER_11_753 VPWR VGND sg13g2_decap_8
XFILLER_3_941 VPWR VGND sg13g2_decap_8
XFILLER_2_462 VPWR VGND sg13g2_decap_8
XFILLER_38_606 VPWR VGND sg13g2_decap_8
XFILLER_1_33 VPWR VGND sg13g2_fill_2
XFILLER_19_831 VPWR VGND sg13g2_decap_8
XFILLER_46_661 VPWR VGND sg13g2_decap_8
XFILLER_1_66 VPWR VGND sg13g2_fill_1
XFILLER_34_823 VPWR VGND sg13g2_decap_8
XFILLER_21_506 VPWR VGND sg13g2_decap_8
XFILLER_14_1006 VPWR VGND sg13g2_decap_8
X_3712_ _1198_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] net595 VPWR
+ VGND sg13g2_nand2_1
X_3643_ net596 _0885_ _1144_ _1145_ _1146_ VPWR VGND sg13g2_nor4_1
X_3574_ net660 _1090_ _1091_ _1092_ VPWR VGND sg13g2_or3_1
X_2525_ _1922_ _1935_ _1938_ VPWR VGND sg13g2_nor2_1
X_2456_ _1873_ _1874_ _1872_ _1875_ VPWR VGND sg13g2_nand3_1
Xhold18 u_ser.shadow_reg\[5\] VPWR VGND net65 sg13g2_dlygate4sd3_1
Xhold29 _0160_ VPWR VGND net76 sg13g2_dlygate4sd3_1
X_2387_ _1806_ _1807_ _1805_ _1808_ VPWR VGND sg13g2_nand3_1
X_4126_ net777 VGND VPWR _0104_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4057_ net784 VGND VPWR _0035_ sap_3_inst.alu.acc\[1\] clknet_5_18__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3008_ net744 sap_3_inst.out\[7\] net673 _0049_ VPWR VGND sg13g2_mux2_1
XFILLER_25_856 VPWR VGND sg13g2_decap_8
XFILLER_40_837 VPWR VGND sg13g2_decap_8
XFILLER_12_539 VPWR VGND sg13g2_decap_8
XFILLER_20_583 VPWR VGND sg13g2_decap_8
XFILLER_4_705 VPWR VGND sg13g2_decap_8
XFILLER_10_64 VPWR VGND sg13g2_fill_1
XFILLER_0_911 VPWR VGND sg13g2_decap_8
XFILLER_0_988 VPWR VGND sg13g2_decap_8
XFILLER_48_948 VPWR VGND sg13g2_decap_8
XFILLER_47_458 VPWR VGND sg13g2_decap_8
XFILLER_16_823 VPWR VGND sg13g2_decap_8
XFILLER_28_694 VPWR VGND sg13g2_decap_8
XFILLER_43_642 VPWR VGND sg13g2_decap_8
XFILLER_37_1017 VPWR VGND sg13g2_decap_8
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_31_848 VPWR VGND sg13g2_decap_8
XFILLER_11_550 VPWR VGND sg13g2_decap_8
XFILLER_7_510 VPWR VGND sg13g2_decap_8
XFILLER_7_587 VPWR VGND sg13g2_decap_8
X_2310_ _1730_ _1729_ _1437_ _1731_ VPWR VGND sg13g2_a21o_1
X_3290_ _0826_ net553 _0825_ VPWR VGND sg13g2_nand2_1
X_2241_ _1506_ _1523_ _1504_ _1662_ VPWR VGND sg13g2_nand3_1
XFILLER_25_4 VPWR VGND sg13g2_fill_1
XFILLER_39_915 VPWR VGND sg13g2_decap_8
X_2172_ _1522_ _1561_ _1518_ _1593_ VPWR VGND _1563_ sg13g2_nand4_1
XFILLER_20_1010 VPWR VGND sg13g2_decap_8
XFILLER_38_458 VPWR VGND sg13g2_fill_1
XFILLER_34_620 VPWR VGND sg13g2_decap_8
XFILLER_22_848 VPWR VGND sg13g2_decap_8
XFILLER_34_697 VPWR VGND sg13g2_decap_8
XFILLER_30_892 VPWR VGND sg13g2_decap_8
X_3626_ net22 _1063_ _1110_ _1133_ VPWR VGND sg13g2_nor3_2
Xoutput19 net19 uio_out[2] VPWR VGND sg13g2_buf_1
X_3557_ _1077_ net592 VPWR VGND _0836_ sg13g2_nand2b_2
X_2508_ VGND VPWR net676 _1920_ _0030_ _1921_ sg13g2_a21oi_1
X_3488_ _1014_ _1015_ net610 _1017_ VPWR VGND _1016_ sg13g2_nand4_1
X_2439_ sap_3_inst.alu.flags\[7\] net542 net675 _0033_ VPWR VGND sg13g2_mux2_1
XFILLER_29_403 VPWR VGND sg13g2_decap_8
XFILLER_29_447 VPWR VGND sg13g2_decap_8
X_4109_ net774 VGND VPWR _0087_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\]
+ clknet_5_3__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_38_970 VPWR VGND sg13g2_decap_8
XFILLER_25_653 VPWR VGND sg13g2_decap_8
XFILLER_40_634 VPWR VGND sg13g2_decap_8
XFILLER_12_325 VPWR VGND sg13g2_fill_2
XFILLER_13_859 VPWR VGND sg13g2_decap_8
XFILLER_21_870 VPWR VGND sg13g2_decap_8
XFILLER_4_502 VPWR VGND sg13g2_decap_8
XFILLER_4_579 VPWR VGND sg13g2_decap_8
Xclkbuf_5_17__f_sap_3_inst.alu.clk_regs clknet_4_8_0_sap_3_inst.alu.clk_regs clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_48_745 VPWR VGND sg13g2_decap_8
XFILLER_0_785 VPWR VGND sg13g2_decap_8
XFILLER_16_620 VPWR VGND sg13g2_decap_8
XFILLER_28_491 VPWR VGND sg13g2_decap_8
XFILLER_44_962 VPWR VGND sg13g2_decap_8
XFILLER_16_697 VPWR VGND sg13g2_decap_8
XFILLER_31_645 VPWR VGND sg13g2_decap_8
X_2790_ _0358_ _0355_ _0356_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_874 VPWR VGND sg13g2_decap_8
X_3411_ _0943_ _1468_ net612 VPWR VGND sg13g2_nand2_1
X_3342_ VGND VPWR net582 _0874_ _0877_ net562 sg13g2_a21oi_1
X_3273_ _0658_ _0670_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] _0809_
+ VPWR VGND _0710_ sg13g2_nand4_1
X_2224_ _1645_ _1605_ _1644_ VPWR VGND sg13g2_nand2_1
XFILLER_39_712 VPWR VGND sg13g2_decap_8
X_2155_ _1561_ _1573_ _1522_ _1576_ VPWR VGND sg13g2_nand3_1
XFILLER_27_907 VPWR VGND sg13g2_decap_8
XFILLER_39_789 VPWR VGND sg13g2_decap_8
X_2086_ _1507_ net739 VPWR VGND net742 sg13g2_nand2b_2
XFILLER_35_940 VPWR VGND sg13g2_decap_8
XFILLER_34_494 VPWR VGND sg13g2_decap_8
XFILLER_10_818 VPWR VGND sg13g2_decap_8
XFILLER_22_645 VPWR VGND sg13g2_decap_8
X_2988_ _0549_ VPWR _0550_ VGND _0323_ _0542_ sg13g2_o21ai_1
X_3609_ VGND VPWR net16 _1078_ _1122_ _0632_ sg13g2_a21oi_1
XFILLER_1_527 VPWR VGND sg13g2_decap_8
XFILLER_27_1005 VPWR VGND sg13g2_decap_8
XFILLER_29_200 VPWR VGND sg13g2_fill_1
XFILLER_45_737 VPWR VGND sg13g2_decap_8
XFILLER_18_929 VPWR VGND sg13g2_decap_8
XFILLER_26_940 VPWR VGND sg13g2_decap_8
XFILLER_25_450 VPWR VGND sg13g2_decap_8
XFILLER_16_85 VPWR VGND sg13g2_fill_2
XFILLER_41_976 VPWR VGND sg13g2_decap_8
XFILLER_40_453 VPWR VGND sg13g2_fill_2
XFILLER_13_656 VPWR VGND sg13g2_decap_8
XFILLER_9_649 VPWR VGND sg13g2_decap_8
XFILLER_32_84 VPWR VGND sg13g2_fill_1
XFILLER_5_866 VPWR VGND sg13g2_decap_8
XFILLER_0_582 VPWR VGND sg13g2_decap_8
XFILLER_48_542 VPWR VGND sg13g2_decap_8
XFILLER_35_247 VPWR VGND sg13g2_fill_1
XFILLER_36_759 VPWR VGND sg13g2_decap_8
X_3960_ _1387_ VPWR _0175_ VGND net603 _1190_ sg13g2_o21ai_1
XFILLER_17_962 VPWR VGND sg13g2_decap_8
XFILLER_32_910 VPWR VGND sg13g2_decap_8
X_2911_ _0474_ VPWR _0475_ VGND _0471_ _0473_ sg13g2_o21ai_1
X_3891_ _1331_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] net721
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_31_442 VPWR VGND sg13g2_fill_2
X_2842_ net554 _0381_ _0408_ _0409_ VPWR VGND sg13g2_nor3_1
XFILLER_32_987 VPWR VGND sg13g2_decap_8
X_2773_ net760 _0328_ _0342_ VPWR VGND sg13g2_nor2_1
XFILLER_8_671 VPWR VGND sg13g2_decap_8
XFILLER_7_181 VPWR VGND sg13g2_fill_2
Xfanout606 net607 net606 VPWR VGND sg13g2_buf_8
Xfanout617 _0310_ net617 VPWR VGND sg13g2_buf_8
Xfanout639 _1794_ net639 VPWR VGND sg13g2_buf_8
Xfanout628 _1799_ net628 VPWR VGND sg13g2_buf_8
X_3325_ net575 _0860_ _0861_ VPWR VGND sg13g2_nor2_1
X_3256_ _0792_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] net593 VPWR
+ VGND sg13g2_nand2_1
X_2207_ _1577_ _1626_ _1628_ VPWR VGND sg13g2_nor2_1
X_3187_ VPWR VGND _0694_ net665 _0691_ _0653_ _0723_ _0656_ sg13g2_a221oi_1
XFILLER_27_704 VPWR VGND sg13g2_decap_8
XFILLER_39_586 VPWR VGND sg13g2_decap_8
X_2138_ _1559_ net711 net710 VPWR VGND sg13g2_nand2_2
X_2069_ VPWR _1492_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_23_976 VPWR VGND sg13g2_decap_8
XFILLER_10_615 VPWR VGND sg13g2_decap_8
XFILLER_2_847 VPWR VGND sg13g2_decap_8
XFILLER_49_339 VPWR VGND sg13g2_decap_8
XFILLER_1_379 VPWR VGND sg13g2_fill_1
XFILLER_18_726 VPWR VGND sg13g2_decap_8
XFILLER_45_534 VPWR VGND sg13g2_decap_8
XFILLER_33_718 VPWR VGND sg13g2_decap_8
XFILLER_14_943 VPWR VGND sg13g2_decap_8
XFILLER_41_773 VPWR VGND sg13g2_decap_8
XFILLER_5_663 VPWR VGND sg13g2_decap_8
XFILLER_4_55 VPWR VGND sg13g2_decap_8
X_3110_ _0646_ _0645_ _1594_ _0644_ _1601_ VPWR VGND sg13g2_a22oi_1
XFILLER_1_891 VPWR VGND sg13g2_decap_8
X_4090_ net778 VGND VPWR _0068_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[1\]
+ clknet_5_1__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
X_3041_ _0588_ VPWR _0055_ VGND _1920_ net667 sg13g2_o21ai_1
XFILLER_36_556 VPWR VGND sg13g2_decap_8
XFILLER_24_729 VPWR VGND sg13g2_decap_8
X_3943_ _1377_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] _1312_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_17_1004 VPWR VGND sg13g2_decap_8
X_3874_ _1497_ _1498_ sap_3_inst.reg_file.array_serializer_inst.word_index\[3\] sap_3_inst.reg_file.array_serializer_inst.word_index\[2\]
+ _1315_ VPWR VGND sg13g2_nor4_1
XFILLER_32_784 VPWR VGND sg13g2_decap_8
X_2825_ _0392_ _0359_ _0391_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_20_968 VPWR VGND sg13g2_decap_8
X_2756_ _0325_ _0200_ _0316_ VPWR VGND sg13g2_nand2_1
X_2687_ net713 net712 _0277_ _0278_ _0279_ VPWR VGND sg13g2_nor4_1
X_3308_ net660 net666 _0844_ VPWR VGND sg13g2_and2_1
X_3239_ _0770_ _0772_ _0773_ _0774_ _0775_ VPWR VGND sg13g2_and4_1
XFILLER_27_501 VPWR VGND sg13g2_decap_8
XFILLER_39_361 VPWR VGND sg13g2_fill_1
XFILLER_27_578 VPWR VGND sg13g2_decap_8
XFILLER_42_559 VPWR VGND sg13g2_decap_8
Xfanout32 net18 net32 VPWR VGND sg13g2_buf_2
XFILLER_23_773 VPWR VGND sg13g2_decap_8
XFILLER_11_935 VPWR VGND sg13g2_decap_8
XFILLER_13_64 VPWR VGND sg13g2_fill_2
XFILLER_2_644 VPWR VGND sg13g2_decap_8
XFILLER_46_843 VPWR VGND sg13g2_decap_8
XFILLER_18_523 VPWR VGND sg13g2_decap_8
XFILLER_45_342 VPWR VGND sg13g2_decap_8
XFILLER_33_515 VPWR VGND sg13g2_decap_8
XFILLER_14_740 VPWR VGND sg13g2_decap_8
XFILLER_41_570 VPWR VGND sg13g2_decap_8
Xclkload13 clknet_5_10__leaf_sap_3_inst.alu.clk_regs clkload13/X VPWR VGND sg13g2_buf_1
XFILLER_9_298 VPWR VGND sg13g2_fill_2
X_2610_ _0207_ net628 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] net632
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] VPWR VGND sg13g2_a22oi_1
X_3590_ VPWR VGND net589 net583 _0975_ _0971_ _1105_ _0972_ sg13g2_a221oi_1
X_2541_ _1954_ _1945_ _1953_ VPWR VGND sg13g2_nand2_1
XFILLER_5_460 VPWR VGND sg13g2_decap_8
X_2472_ _1889_ net6 _1847_ VPWR VGND sg13g2_nand2_1
X_4211_ net783 VGND VPWR _0188_ sap_3_outputReg_serial clknet_3_1__leaf_clk sg13g2_dfrbpq_1
X_4142_ net776 VGND VPWR _0120_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\]
+ clknet_5_9__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4073_ net785 VGND VPWR _0051_ sap_3_inst.alu.tmp\[0\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3024_ _0202_ _0576_ _1950_ _0577_ VPWR VGND sg13g2_nand3_1
XFILLER_37_821 VPWR VGND sg13g2_decap_8
XFILLER_24_526 VPWR VGND sg13g2_decap_8
XFILLER_37_898 VPWR VGND sg13g2_decap_8
X_3926_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] net761
+ _1362_ net763 sg13g2_a21oi_1
XFILLER_32_581 VPWR VGND sg13g2_decap_8
Xclkload7 clknet_1_0__leaf_clk_div_out clkload7/X VPWR VGND sg13g2_buf_1
XFILLER_20_765 VPWR VGND sg13g2_decap_8
X_3857_ _1284_ VPWR _1299_ VGND net48 _1281_ sg13g2_o21ai_1
X_2808_ _0365_ _0375_ _0363_ _0376_ VPWR VGND sg13g2_nand3_1
X_3788_ net600 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[1\] _1250_ _0140_
+ VPWR VGND sg13g2_a21o_1
X_2739_ net683 _1845_ _0307_ _0308_ VPWR VGND sg13g2_nor3_1
XFILLER_1_9 VPWR VGND sg13g2_fill_1
XFILLER_28_876 VPWR VGND sg13g2_decap_8
XFILLER_43_824 VPWR VGND sg13g2_decap_8
XFILLER_30_507 VPWR VGND sg13g2_decap_8
XFILLER_11_732 VPWR VGND sg13g2_decap_8
XFILLER_23_570 VPWR VGND sg13g2_decap_8
XFILLER_7_769 VPWR VGND sg13g2_decap_8
XFILLER_3_920 VPWR VGND sg13g2_decap_8
XFILLER_2_441 VPWR VGND sg13g2_decap_8
XFILLER_3_997 VPWR VGND sg13g2_decap_8
XFILLER_19_810 VPWR VGND sg13g2_decap_8
XFILLER_46_640 VPWR VGND sg13g2_decap_8
XFILLER_1_78 VPWR VGND sg13g2_fill_2
XFILLER_34_802 VPWR VGND sg13g2_decap_8
XFILLER_19_887 VPWR VGND sg13g2_decap_8
XFILLER_34_879 VPWR VGND sg13g2_decap_8
X_3711_ VGND VPWR _1458_ net594 _0116_ _1197_ sg13g2_a21oi_1
X_3642_ net10 net32 net568 _1145_ VPWR VGND sg13g2_mux2_1
X_3573_ _0633_ _0900_ _1091_ VPWR VGND sg13g2_nor2_1
XFILLER_46_0 VPWR VGND sg13g2_fill_2
X_2524_ VPWR _1937_ _1936_ VGND sg13g2_inv_1
X_2455_ _1874_ net626 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] net630
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2386_ _1807_ net629 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] net677
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\] VPWR VGND sg13g2_a22oi_1
Xhold19 regFile_serial VPWR VGND net66 sg13g2_dlygate4sd3_1
XFILLER_29_629 VPWR VGND sg13g2_decap_8
X_4125_ net774 VGND VPWR _0103_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4056_ net785 VGND VPWR _0034_ sap_3_inst.alu.acc\[0\] clknet_5_18__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3007_ net746 sap_3_inst.out\[6\] net674 _0048_ VPWR VGND sg13g2_mux2_1
XFILLER_25_835 VPWR VGND sg13g2_decap_8
XFILLER_36_150 VPWR VGND sg13g2_fill_2
XFILLER_37_695 VPWR VGND sg13g2_decap_8
XFILLER_40_816 VPWR VGND sg13g2_decap_8
XFILLER_12_518 VPWR VGND sg13g2_decap_8
X_3909_ _1347_ net761 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] net721
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_562 VPWR VGND sg13g2_decap_8
XFILLER_10_32 VPWR VGND sg13g2_fill_1
XFILLER_48_927 VPWR VGND sg13g2_decap_8
XFILLER_0_967 VPWR VGND sg13g2_decap_8
XFILLER_47_437 VPWR VGND sg13g2_decap_8
XFILLER_16_802 VPWR VGND sg13g2_decap_8
XFILLER_28_673 VPWR VGND sg13g2_decap_8
XFILLER_43_621 VPWR VGND sg13g2_decap_8
XFILLER_42_131 VPWR VGND sg13g2_fill_1
XFILLER_16_879 VPWR VGND sg13g2_decap_8
XFILLER_31_827 VPWR VGND sg13g2_decap_8
XFILLER_43_698 VPWR VGND sg13g2_decap_8
XFILLER_24_890 VPWR VGND sg13g2_decap_8
XFILLER_7_566 VPWR VGND sg13g2_decap_8
X_2240_ net723 _1507_ net722 _1661_ VPWR VGND sg13g2_nor3_1
XFILLER_3_794 VPWR VGND sg13g2_decap_8
X_2171_ _1518_ _1522_ _1561_ _1563_ _1592_ VPWR VGND sg13g2_and4_1
XFILLER_19_684 VPWR VGND sg13g2_decap_8
XFILLER_22_827 VPWR VGND sg13g2_decap_8
XFILLER_33_131 VPWR VGND sg13g2_fill_1
XFILLER_34_676 VPWR VGND sg13g2_decap_8
XFILLER_33_175 VPWR VGND sg13g2_fill_1
XFILLER_30_871 VPWR VGND sg13g2_decap_8
X_3625_ _1131_ VPWR _0095_ VGND _1060_ _1132_ sg13g2_o21ai_1
X_3556_ net558 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] _1076_ _0082_
+ VPWR VGND sg13g2_a21o_1
XFILLER_1_709 VPWR VGND sg13g2_decap_8
X_2507_ sap_3_inst.alu.flags\[4\] net676 _1921_ VPWR VGND sg13g2_nor2_1
X_3487_ _1016_ net658 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] net606
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2438_ _1858_ net675 VPWR VGND sg13g2_inv_2
XFILLER_5_1027 VPWR VGND sg13g2_fill_2
X_2369_ _1502_ _1526_ _1788_ _1790_ VGND VPWR _1789_ sg13g2_nor4_2
XFILLER_45_919 VPWR VGND sg13g2_decap_8
X_4108_ net782 VGND VPWR _0086_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\]
+ clknet_5_6__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4039_ net784 VGND VPWR _0021_ u_ser.shadow_reg\[3\] clknet_3_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_25_632 VPWR VGND sg13g2_decap_8
XFILLER_40_613 VPWR VGND sg13g2_decap_8
XFILLER_13_838 VPWR VGND sg13g2_decap_8
XFILLER_4_558 VPWR VGND sg13g2_decap_8
XFILLER_0_764 VPWR VGND sg13g2_decap_8
XFILLER_48_724 VPWR VGND sg13g2_decap_8
XFILLER_29_993 VPWR VGND sg13g2_decap_8
XFILLER_44_941 VPWR VGND sg13g2_decap_8
XFILLER_28_470 VPWR VGND sg13g2_decap_8
XFILLER_16_676 VPWR VGND sg13g2_decap_8
XFILLER_43_495 VPWR VGND sg13g2_decap_8
XFILLER_15_186 VPWR VGND sg13g2_fill_1
XFILLER_31_624 VPWR VGND sg13g2_decap_8
XFILLER_12_882 VPWR VGND sg13g2_decap_8
XFILLER_8_853 VPWR VGND sg13g2_decap_8
X_3410_ _0941_ VPWR _0942_ VGND _1474_ net589 sg13g2_o21ai_1
Xclkbuf_4_11_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_11_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3341_ _0821_ _0875_ _0876_ VPWR VGND sg13g2_and2_1
XFILLER_3_591 VPWR VGND sg13g2_decap_8
X_3272_ _0802_ _0807_ _0808_ VPWR VGND sg13g2_and2_1
X_2223_ _1623_ _1636_ _1578_ _1644_ VPWR VGND _1642_ sg13g2_nand4_1
X_2154_ net735 net737 _1562_ _1575_ VGND VPWR _1574_ sg13g2_nor4_2
XFILLER_39_768 VPWR VGND sg13g2_decap_8
XFILLER_26_429 VPWR VGND sg13g2_decap_8
X_2085_ net742 net739 _1506_ VPWR VGND sg13g2_nor2b_2
XFILLER_22_624 VPWR VGND sg13g2_decap_8
XFILLER_35_996 VPWR VGND sg13g2_decap_8
X_2987_ _0545_ _0546_ _0547_ _0548_ _0549_ VPWR VGND sg13g2_and4_1
X_3608_ _1121_ net24 net570 VPWR VGND sg13g2_nand2_1
XFILLER_1_506 VPWR VGND sg13g2_decap_8
X_3539_ _1058_ VPWR _0079_ VGND _1060_ _1062_ sg13g2_o21ai_1
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
XFILLER_18_908 VPWR VGND sg13g2_decap_8
XFILLER_45_716 VPWR VGND sg13g2_decap_8
XFILLER_44_226 VPWR VGND sg13g2_fill_2
XFILLER_13_635 VPWR VGND sg13g2_decap_8
XFILLER_26_996 VPWR VGND sg13g2_decap_8
XFILLER_41_955 VPWR VGND sg13g2_decap_8
XFILLER_12_123 VPWR VGND sg13g2_fill_2
XFILLER_40_487 VPWR VGND sg13g2_decap_8
XFILLER_8_116 VPWR VGND sg13g2_fill_1
XFILLER_9_628 VPWR VGND sg13g2_decap_8
XFILLER_5_845 VPWR VGND sg13g2_decap_8
XFILLER_10_1021 VPWR VGND sg13g2_decap_8
XFILLER_0_561 VPWR VGND sg13g2_decap_8
XFILLER_48_521 VPWR VGND sg13g2_decap_8
XFILLER_48_598 VPWR VGND sg13g2_decap_8
XFILLER_17_941 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_3_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_29_790 VPWR VGND sg13g2_decap_8
XFILLER_36_738 VPWR VGND sg13g2_decap_8
XFILLER_16_440 VPWR VGND sg13g2_fill_2
X_2910_ VGND VPWR _0471_ _0473_ _0474_ _1937_ sg13g2_a21oi_1
X_3890_ _1330_ _1312_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] _1311_
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_32_966 VPWR VGND sg13g2_decap_8
X_2841_ VPWR VGND _0407_ net616 _0406_ sap_3_inst.alu.act\[2\] _0408_ net669 sg13g2_a221oi_1
X_2772_ _0341_ _0340_ _0320_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_498 VPWR VGND sg13g2_decap_8
XFILLER_8_650 VPWR VGND sg13g2_decap_8
Xfanout618 _1949_ net618 VPWR VGND sg13g2_buf_8
Xfanout607 _0721_ net607 VPWR VGND sg13g2_buf_8
X_3324_ _0860_ _0744_ _0858_ VPWR VGND sg13g2_xnor2_1
Xfanout629 net630 net629 VPWR VGND sg13g2_buf_8
X_3255_ _0791_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] net642 VPWR
+ VGND sg13g2_nand2_1
X_2206_ _1627_ net711 net704 VPWR VGND sg13g2_nand2_2
XFILLER_2_1008 VPWR VGND sg13g2_decap_8
X_3186_ _0722_ _0695_ _0719_ VPWR VGND sg13g2_nand2_2
XFILLER_39_565 VPWR VGND sg13g2_decap_8
X_2137_ net711 net710 _1558_ VPWR VGND sg13g2_and2_1
XFILLER_26_226 VPWR VGND sg13g2_fill_2
X_2068_ VPWR _1491_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_35_793 VPWR VGND sg13g2_decap_8
XFILLER_22_443 VPWR VGND sg13g2_fill_2
XFILLER_23_955 VPWR VGND sg13g2_decap_8
XFILLER_22_498 VPWR VGND sg13g2_decap_8
XFILLER_2_826 VPWR VGND sg13g2_decap_8
XFILLER_49_318 VPWR VGND sg13g2_decap_8
XFILLER_18_705 VPWR VGND sg13g2_decap_8
XFILLER_45_513 VPWR VGND sg13g2_decap_8
XFILLER_14_922 VPWR VGND sg13g2_decap_8
XFILLER_26_793 VPWR VGND sg13g2_decap_8
XFILLER_41_752 VPWR VGND sg13g2_decap_8
XFILLER_14_999 VPWR VGND sg13g2_decap_8
XFILLER_5_642 VPWR VGND sg13g2_decap_8
XFILLER_4_34 VPWR VGND sg13g2_fill_1
XFILLER_4_67 VPWR VGND sg13g2_fill_1
XFILLER_1_870 VPWR VGND sg13g2_decap_8
XFILLER_49_885 VPWR VGND sg13g2_decap_8
X_3040_ _0588_ sap_3_inst.alu.tmp\[4\] net667 VPWR VGND sg13g2_nand2_1
XFILLER_48_395 VPWR VGND sg13g2_decap_8
XFILLER_36_535 VPWR VGND sg13g2_decap_8
XFILLER_24_708 VPWR VGND sg13g2_decap_8
X_3942_ _1376_ net761 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] _1306_
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3873_ _1498_ _1304_ _1314_ VPWR VGND sg13g2_nor2_1
XFILLER_32_763 VPWR VGND sg13g2_decap_8
X_2824_ _0391_ _0382_ _0389_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_947 VPWR VGND sg13g2_decap_8
X_2755_ _0200_ _0316_ _0324_ VPWR VGND sg13g2_and2_1
XFILLER_9_992 VPWR VGND sg13g2_decap_8
X_2686_ VGND VPWR net698 _1713_ _0278_ _1823_ sg13g2_a21oi_1
XFILLER_24_1009 VPWR VGND sg13g2_decap_8
X_3307_ _0843_ net660 _0633_ VPWR VGND sg13g2_nand2_2
X_3238_ _0774_ _0768_ _0769_ _0771_ VPWR VGND sg13g2_and3_1
X_3169_ _1730_ _0599_ net682 _0705_ VPWR VGND _0704_ sg13g2_nand4_1
XFILLER_27_557 VPWR VGND sg13g2_decap_8
XFILLER_42_538 VPWR VGND sg13g2_decap_8
XFILLER_35_590 VPWR VGND sg13g2_decap_8
XFILLER_11_914 VPWR VGND sg13g2_decap_8
XFILLER_23_752 VPWR VGND sg13g2_decap_8
XFILLER_2_623 VPWR VGND sg13g2_decap_8
XFILLER_1_155 VPWR VGND sg13g2_decap_8
XFILLER_18_502 VPWR VGND sg13g2_decap_8
XFILLER_46_822 VPWR VGND sg13g2_decap_8
XFILLER_46_899 VPWR VGND sg13g2_decap_8
XFILLER_45_387 VPWR VGND sg13g2_decap_8
XFILLER_18_579 VPWR VGND sg13g2_decap_8
XFILLER_26_590 VPWR VGND sg13g2_decap_8
XFILLER_14_796 VPWR VGND sg13g2_decap_8
Xclkload14 VPWR clkload14/Y clknet_5_13__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_2540_ _1953_ _1946_ _1952_ VPWR VGND sg13g2_nand2_1
XFILLER_6_995 VPWR VGND sg13g2_decap_8
X_2471_ _1888_ _1828_ sap_3_inst.alu.flags\[5\] _1827_ net747 VPWR VGND sg13g2_a22oi_1
X_4210_ net783 VGND VPWR _0187_ u_ser.state\[1\] clknet_3_1__leaf_clk sg13g2_dfrbpq_2
X_4141_ net774 VGND VPWR _0119_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4072_ net787 VGND VPWR _0050_ sap_3_inst.alu.carry clknet_5_18__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_37_800 VPWR VGND sg13g2_decap_8
XFILLER_49_682 VPWR VGND sg13g2_decap_8
X_3023_ _0576_ sap_3_inst.alu.flags\[1\] net618 VPWR VGND sg13g2_nand2_1
XFILLER_37_877 VPWR VGND sg13g2_decap_8
XFILLER_24_505 VPWR VGND sg13g2_decap_8
XFILLER_36_398 VPWR VGND sg13g2_fill_1
X_3925_ _1361_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] net721
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_32_560 VPWR VGND sg13g2_decap_8
XFILLER_20_744 VPWR VGND sg13g2_decap_8
Xclkload8 VPWR clkload8/Y clknet_5_1__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_3856_ _1297_ VPWR _1298_ VGND sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\]
+ _1292_ sg13g2_o21ai_1
X_2807_ VPWR VGND _0369_ _0374_ _0366_ net756 _0375_ net572 sg13g2_a221oi_1
X_3787_ net600 _1184_ _1185_ _1250_ VPWR VGND sg13g2_nor3_1
X_2738_ _1511_ net695 _1716_ _0307_ VPWR VGND sg13g2_nor3_1
X_2669_ _1646_ VPWR _0261_ VGND _1575_ _1583_ sg13g2_o21ai_1
XFILLER_8_1014 VPWR VGND sg13g2_decap_8
XFILLER_47_619 VPWR VGND sg13g2_decap_8
XFILLER_43_803 VPWR VGND sg13g2_decap_8
XFILLER_28_855 VPWR VGND sg13g2_decap_8
XFILLER_15_549 VPWR VGND sg13g2_decap_8
XFILLER_11_711 VPWR VGND sg13g2_decap_8
XFILLER_7_748 VPWR VGND sg13g2_decap_8
XFILLER_11_788 VPWR VGND sg13g2_decap_8
XFILLER_3_976 VPWR VGND sg13g2_decap_8
XFILLER_2_497 VPWR VGND sg13g2_decap_8
Xfanout790 net791 net790 VPWR VGND sg13g2_buf_8
XFILLER_19_866 VPWR VGND sg13g2_decap_8
XFILLER_46_696 VPWR VGND sg13g2_decap_8
XFILLER_45_195 VPWR VGND sg13g2_fill_1
XFILLER_33_313 VPWR VGND sg13g2_fill_1
XFILLER_34_858 VPWR VGND sg13g2_decap_8
XFILLER_14_593 VPWR VGND sg13g2_decap_8
X_3710_ net32 net594 _1144_ _1197_ VPWR VGND sg13g2_nor3_1
X_3641_ net576 _0874_ _1144_ VPWR VGND sg13g2_nor2_1
X_3572_ VGND VPWR net11 _1078_ _1090_ _1089_ sg13g2_a21oi_1
X_2523_ _1922_ _1931_ _1936_ VPWR VGND sg13g2_nor2b_2
XFILLER_6_792 VPWR VGND sg13g2_decap_8
X_2454_ _1873_ _1803_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\] net639
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2385_ _1806_ net619 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] net633
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_0 VPWR VGND sg13g2_fill_1
X_4124_ net782 VGND VPWR _0102_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\]
+ clknet_5_26__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_608 VPWR VGND sg13g2_decap_8
XFILLER_28_129 VPWR VGND sg13g2_fill_1
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
X_4055_ net799 VGND VPWR _0033_ sap_3_inst.alu.flags\[7\] net47 sg13g2_dfrbpq_1
X_3006_ net749 sap_3_inst.out\[5\] net674 _0047_ VPWR VGND sg13g2_mux2_1
XFILLER_25_814 VPWR VGND sg13g2_decap_8
XFILLER_37_674 VPWR VGND sg13g2_decap_8
Xclkbuf_5_25__f_sap_3_inst.alu.clk_regs clknet_4_12_0_sap_3_inst.alu.clk_regs clknet_5_25__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_20_541 VPWR VGND sg13g2_decap_8
X_3908_ _1346_ _1313_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] _1311_
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] VPWR VGND sg13g2_a22oi_1
X_3839_ net769 _1282_ _1285_ VPWR VGND sg13g2_nor2_1
XFILLER_0_946 VPWR VGND sg13g2_decap_8
XFILLER_48_906 VPWR VGND sg13g2_decap_8
XFILLER_47_416 VPWR VGND sg13g2_decap_8
XFILLER_28_652 VPWR VGND sg13g2_decap_8
XFILLER_43_600 VPWR VGND sg13g2_decap_8
XFILLER_16_858 VPWR VGND sg13g2_decap_8
XFILLER_43_677 VPWR VGND sg13g2_decap_8
XFILLER_31_806 VPWR VGND sg13g2_decap_8
XFILLER_30_338 VPWR VGND sg13g2_fill_1
XFILLER_11_585 VPWR VGND sg13g2_decap_8
XFILLER_7_545 VPWR VGND sg13g2_decap_8
XFILLER_3_773 VPWR VGND sg13g2_decap_8
X_2170_ _1522_ _1563_ _1591_ VPWR VGND sg13g2_and2_1
XFILLER_47_983 VPWR VGND sg13g2_decap_8
XFILLER_19_663 VPWR VGND sg13g2_decap_8
XFILLER_46_493 VPWR VGND sg13g2_decap_8
XFILLER_22_806 VPWR VGND sg13g2_decap_8
XFILLER_34_655 VPWR VGND sg13g2_decap_8
XFILLER_30_850 VPWR VGND sg13g2_decap_8
X_3624_ _1061_ VPWR _1132_ VGND net642 _1078_ sg13g2_o21ai_1
X_3555_ _1025_ net558 _1075_ _1076_ VPWR VGND sg13g2_nor3_1
X_3486_ _1015_ net643 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] net651
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2506_ net21 _1920_ VPWR VGND sg13g2_inv_2
X_2437_ net724 _1576_ _1675_ _1857_ VPWR VGND sg13g2_nor3_2
XFILLER_5_1006 VPWR VGND sg13g2_decap_8
X_2368_ VGND VPWR net684 _1774_ _1789_ _1538_ sg13g2_a21oi_1
X_2299_ _1720_ _1510_ net698 net709 VPWR VGND sg13g2_and3_1
X_4107_ net771 VGND VPWR _0085_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\]
+ clknet_5_4__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4038_ net784 VGND VPWR _0020_ u_ser.shadow_reg\[2\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_24_110 VPWR VGND sg13g2_fill_2
XFILLER_25_611 VPWR VGND sg13g2_decap_8
XFILLER_13_817 VPWR VGND sg13g2_decap_8
XFILLER_12_327 VPWR VGND sg13g2_fill_1
XFILLER_25_688 VPWR VGND sg13g2_decap_8
XFILLER_40_669 VPWR VGND sg13g2_decap_8
XFILLER_4_537 VPWR VGND sg13g2_decap_8
XFILLER_48_703 VPWR VGND sg13g2_decap_8
XFILLER_0_743 VPWR VGND sg13g2_decap_8
XFILLER_47_279 VPWR VGND sg13g2_fill_2
XFILLER_29_972 VPWR VGND sg13g2_decap_8
XFILLER_44_920 VPWR VGND sg13g2_decap_8
XFILLER_16_655 VPWR VGND sg13g2_decap_8
XFILLER_44_997 VPWR VGND sg13g2_decap_8
XFILLER_43_474 VPWR VGND sg13g2_decap_8
XFILLER_31_603 VPWR VGND sg13g2_decap_8
XFILLER_8_832 VPWR VGND sg13g2_decap_8
XFILLER_12_861 VPWR VGND sg13g2_decap_8
XFILLER_7_67 VPWR VGND sg13g2_decap_4
X_3340_ VGND VPWR _0875_ _0820_ net561 sg13g2_or2_1
XFILLER_3_570 VPWR VGND sg13g2_decap_8
X_3271_ _0803_ _0804_ _0805_ _0806_ _0807_ VPWR VGND sg13g2_nor4_1
X_2222_ _1643_ _1578_ _1642_ VPWR VGND sg13g2_nand2_1
X_2153_ _1574_ net741 VPWR VGND net740 sg13g2_nand2b_2
XFILLER_39_747 VPWR VGND sg13g2_decap_8
XFILLER_26_408 VPWR VGND sg13g2_decap_8
XFILLER_47_780 VPWR VGND sg13g2_decap_8
X_2084_ _1505_ sap_3_inst.controller.opcode\[4\] net730 VPWR VGND sg13g2_nand2_1
XFILLER_35_975 VPWR VGND sg13g2_decap_8
XFILLER_22_603 VPWR VGND sg13g2_decap_8
X_2986_ VGND VPWR _0548_ _0327_ net744 sg13g2_or2_1
X_3607_ _0089_ _1115_ _1120_ net590 _1488_ VPWR VGND sg13g2_a22oi_1
X_3538_ _1062_ _1061_ net558 VPWR VGND sg13g2_nand2b_1
X_3469_ VGND VPWR _0998_ _0999_ _0995_ _0982_ sg13g2_a21oi_2
XFILLER_26_975 VPWR VGND sg13g2_decap_8
XFILLER_41_934 VPWR VGND sg13g2_decap_8
XFILLER_13_614 VPWR VGND sg13g2_decap_8
XFILLER_25_485 VPWR VGND sg13g2_decap_8
XFILLER_9_607 VPWR VGND sg13g2_decap_8
XFILLER_40_466 VPWR VGND sg13g2_decap_8
XFILLER_5_824 VPWR VGND sg13g2_decap_8
XFILLER_10_1000 VPWR VGND sg13g2_decap_8
XFILLER_32_75 VPWR VGND sg13g2_fill_1
XFILLER_0_540 VPWR VGND sg13g2_decap_8
XFILLER_48_500 VPWR VGND sg13g2_decap_8
XFILLER_48_577 VPWR VGND sg13g2_decap_8
XFILLER_36_717 VPWR VGND sg13g2_decap_8
XFILLER_17_920 VPWR VGND sg13g2_decap_8
XFILLER_44_794 VPWR VGND sg13g2_decap_8
XFILLER_17_997 VPWR VGND sg13g2_decap_8
X_2840_ VGND VPWR net543 _0387_ _0407_ net669 sg13g2_a21oi_1
XFILLER_32_945 VPWR VGND sg13g2_decap_8
X_2771_ _1949_ _0197_ _0340_ VPWR VGND sg13g2_nor2_2
XFILLER_7_183 VPWR VGND sg13g2_fill_1
Xfanout608 net609 net608 VPWR VGND sg13g2_buf_8
Xfanout619 net620 net619 VPWR VGND sg13g2_buf_8
X_3323_ _0859_ _0797_ _0857_ VPWR VGND sg13g2_nand2_1
XFILLER_21_0 VPWR VGND sg13g2_fill_2
X_3254_ _0790_ net647 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] net650
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2205_ net711 net704 _1626_ VPWR VGND sg13g2_and2_1
XFILLER_39_544 VPWR VGND sg13g2_decap_8
X_3185_ _0695_ _0719_ _0721_ VPWR VGND sg13g2_and2_1
X_2136_ _1557_ net717 VPWR VGND sap_3_inst.controller.stage\[3\] sg13g2_nand2b_2
XFILLER_27_739 VPWR VGND sg13g2_decap_8
X_2067_ _1490_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[7\] VPWR VGND
+ sg13g2_inv_2
XFILLER_23_934 VPWR VGND sg13g2_decap_8
XFILLER_35_772 VPWR VGND sg13g2_decap_8
XFILLER_22_477 VPWR VGND sg13g2_decap_8
X_2969_ VPWR VGND _0531_ net554 _0530_ net547 _0532_ _0310_ sg13g2_a221oi_1
XFILLER_5_109 VPWR VGND sg13g2_decap_4
XFILLER_2_805 VPWR VGND sg13g2_decap_8
XFILLER_40_1026 VPWR VGND sg13g2_fill_2
XFILLER_45_569 VPWR VGND sg13g2_decap_8
XFILLER_14_901 VPWR VGND sg13g2_decap_8
XFILLER_26_772 VPWR VGND sg13g2_decap_8
XFILLER_41_731 VPWR VGND sg13g2_decap_8
XFILLER_9_415 VPWR VGND sg13g2_fill_1
XFILLER_14_978 VPWR VGND sg13g2_decap_8
XFILLER_5_621 VPWR VGND sg13g2_decap_8
XFILLER_5_698 VPWR VGND sg13g2_decap_8
XFILLER_4_79 VPWR VGND sg13g2_fill_2
XFILLER_49_864 VPWR VGND sg13g2_decap_8
XFILLER_48_374 VPWR VGND sg13g2_decap_8
XFILLER_36_514 VPWR VGND sg13g2_decap_8
XFILLER_23_219 VPWR VGND sg13g2_decap_4
XFILLER_44_591 VPWR VGND sg13g2_decap_8
X_3941_ _1280_ net50 _1375_ _0168_ VPWR VGND sg13g2_a21o_1
XFILLER_17_794 VPWR VGND sg13g2_decap_8
XFILLER_32_742 VPWR VGND sg13g2_decap_8
X_3872_ _1498_ _1301_ _1313_ VPWR VGND sg13g2_nor2_2
XFILLER_20_926 VPWR VGND sg13g2_decap_8
X_2823_ _0383_ _0389_ _0390_ VPWR VGND sg13g2_nor2_1
XFILLER_9_971 VPWR VGND sg13g2_decap_8
X_2754_ _0323_ _0200_ _0201_ VPWR VGND sg13g2_nand2_2
X_2685_ VPWR VGND _0276_ _1930_ _0274_ net690 _0277_ net688 sg13g2_a221oi_1
X_3306_ net660 _0633_ _0842_ VPWR VGND sg13g2_and2_1
X_3237_ _0773_ net658 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] net606
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3168_ _1549_ net687 net729 _0704_ VPWR VGND sg13g2_nand3_1
XFILLER_27_536 VPWR VGND sg13g2_decap_8
X_2119_ net723 _1517_ _1521_ _1540_ VGND VPWR _1539_ sg13g2_nor4_2
XFILLER_42_517 VPWR VGND sg13g2_decap_8
X_3099_ _0610_ _0634_ _0635_ VPWR VGND sg13g2_and2_1
XFILLER_23_731 VPWR VGND sg13g2_decap_8
XFILLER_13_44 VPWR VGND sg13g2_fill_2
XFILLER_2_602 VPWR VGND sg13g2_decap_8
XFILLER_1_134 VPWR VGND sg13g2_decap_4
XFILLER_2_679 VPWR VGND sg13g2_decap_8
XFILLER_46_801 VPWR VGND sg13g2_decap_8
XFILLER_46_878 VPWR VGND sg13g2_decap_8
XFILLER_45_322 VPWR VGND sg13g2_fill_2
XFILLER_18_558 VPWR VGND sg13g2_decap_8
XFILLER_14_775 VPWR VGND sg13g2_decap_8
XFILLER_9_212 VPWR VGND sg13g2_fill_2
Xclkload15 VPWR clkload15/Y clknet_5_17__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_2470_ _1887_ _1881_ _1886_ net639 _1475_ VPWR VGND sg13g2_a22oi_1
XFILLER_6_974 VPWR VGND sg13g2_decap_8
XFILLER_5_495 VPWR VGND sg13g2_decap_8
X_4140_ net795 VGND VPWR _0118_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\]
+ clknet_5_25__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_49_661 VPWR VGND sg13g2_decap_8
X_4071_ net788 VGND VPWR _0049_ sap_3_inst.out\[7\] clknet_5_18__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3022_ _0575_ _0324_ _0574_ VPWR VGND sg13g2_nand2_1
XFILLER_37_856 VPWR VGND sg13g2_decap_8
XFILLER_17_591 VPWR VGND sg13g2_decap_8
X_3924_ _1360_ _1308_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] _1306_
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_723 VPWR VGND sg13g2_decap_8
Xclkload9 VPWR clkload9/Y clknet_5_3__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
X_3855_ _1296_ _1282_ _1297_ VPWR VGND sg13g2_nor2b_1
X_2806_ VGND VPWR net759 _0372_ _0374_ _0373_ sg13g2_a21oi_1
XFILLER_30_1025 VPWR VGND sg13g2_decap_4
X_3786_ net600 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[0\] _1249_ _0139_
+ VPWR VGND sg13g2_a21o_1
X_2737_ VGND VPWR _0299_ _0305_ _0306_ _1715_ sg13g2_a21oi_1
X_2668_ _1561_ _1591_ net700 _0260_ VPWR VGND _1620_ sg13g2_nand4_1
X_2599_ VPWR _2008_ net564 VGND sg13g2_inv_1
XFILLER_27_300 VPWR VGND sg13g2_fill_1
XFILLER_28_834 VPWR VGND sg13g2_decap_8
XFILLER_43_859 VPWR VGND sg13g2_decap_8
XFILLER_15_528 VPWR VGND sg13g2_decap_8
XFILLER_11_767 VPWR VGND sg13g2_decap_8
XFILLER_7_727 VPWR VGND sg13g2_decap_8
XFILLER_3_955 VPWR VGND sg13g2_decap_8
XFILLER_2_476 VPWR VGND sg13g2_decap_8
Xfanout780 net781 net780 VPWR VGND sg13g2_buf_8
Xfanout791 net792 net791 VPWR VGND sg13g2_buf_8
XFILLER_19_845 VPWR VGND sg13g2_decap_8
XFILLER_46_675 VPWR VGND sg13g2_decap_8
XFILLER_34_837 VPWR VGND sg13g2_decap_8
XFILLER_42_881 VPWR VGND sg13g2_decap_8
XFILLER_14_572 VPWR VGND sg13g2_decap_8
X_3640_ net597 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] _1143_ _0099_
+ VPWR VGND sg13g2_a21o_1
X_3571_ net570 net19 net666 _1089_ VPWR VGND sg13g2_a21o_1
XFILLER_6_771 VPWR VGND sg13g2_decap_8
X_2522_ _1928_ _1931_ _1934_ _1935_ VPWR VGND sg13g2_nor3_1
XFILLER_46_2 VPWR VGND sg13g2_fill_1
X_2453_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\] net621
+ net627 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] _1872_ net677 sg13g2_a221oi_1
X_2384_ _1805_ net627 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] net635
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4123_ net771 VGND VPWR _0101_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\]
+ clknet_5_4__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4054_ net793 VGND VPWR _0032_ sap_3_inst.alu.flags\[6\] net46 sg13g2_dfrbpq_1
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
X_3005_ net752 sap_3_inst.out\[4\] net674 _0046_ VPWR VGND sg13g2_mux2_1
XFILLER_37_653 VPWR VGND sg13g2_decap_8
XFILLER_20_520 VPWR VGND sg13g2_decap_8
X_3907_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] _1316_
+ _1345_ net762 sg13g2_a21oi_1
X_3838_ _0156_ _1281_ _1284_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_3_sap_3_inst.alu.clk clknet_1_0__leaf_sap_3_inst.alu.clk clknet_leaf_3_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_20_597 VPWR VGND sg13g2_decap_8
X_3769_ net13 net599 _1236_ _1237_ VPWR VGND sg13g2_nor3_1
XFILLER_4_719 VPWR VGND sg13g2_decap_8
XFILLER_0_925 VPWR VGND sg13g2_decap_8
XFILLER_19_76 VPWR VGND sg13g2_fill_2
XFILLER_28_631 VPWR VGND sg13g2_decap_8
XFILLER_15_303 VPWR VGND sg13g2_fill_2
XFILLER_15_314 VPWR VGND sg13g2_fill_2
XFILLER_16_837 VPWR VGND sg13g2_decap_8
XFILLER_43_656 VPWR VGND sg13g2_decap_8
XFILLER_15_347 VPWR VGND sg13g2_fill_1
XFILLER_42_155 VPWR VGND sg13g2_fill_2
XFILLER_7_524 VPWR VGND sg13g2_decap_8
XFILLER_11_564 VPWR VGND sg13g2_decap_8
XFILLER_13_1020 VPWR VGND sg13g2_decap_8
XFILLER_3_752 VPWR VGND sg13g2_decap_8
XFILLER_2_284 VPWR VGND sg13g2_fill_1
XFILLER_39_929 VPWR VGND sg13g2_decap_8
XFILLER_19_642 VPWR VGND sg13g2_decap_8
XFILLER_47_962 VPWR VGND sg13g2_decap_8
XFILLER_20_1024 VPWR VGND sg13g2_decap_4
XFILLER_46_472 VPWR VGND sg13g2_decap_8
XFILLER_34_634 VPWR VGND sg13g2_decap_8
XFILLER_15_892 VPWR VGND sg13g2_decap_8
X_3623_ _1131_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] net550 VPWR
+ VGND sg13g2_nand2_1
X_3554_ net24 net578 _1033_ _1074_ _1075_ VPWR VGND sg13g2_nor4_1
X_3485_ _1014_ net646 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] net649
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2505_ _1920_ _1909_ _1910_ _1919_ VPWR VGND sg13g2_and3_2
X_2436_ _1811_ _1849_ _1856_ net542 VPWR VGND sg13g2_or3_1
X_2367_ VGND VPWR _1775_ _1787_ _1788_ net712 sg13g2_a21oi_1
X_2298_ VPWR VGND _1547_ _1715_ _1718_ _1697_ _1719_ _1711_ sg13g2_a221oi_1
X_4106_ net770 VGND VPWR _0084_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_44_409 VPWR VGND sg13g2_decap_8
X_4037_ net784 VGND VPWR _0019_ u_ser.shadow_reg\[1\] clknet_3_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_38_984 VPWR VGND sg13g2_decap_8
XFILLER_25_667 VPWR VGND sg13g2_decap_8
XFILLER_40_648 VPWR VGND sg13g2_decap_8
XFILLER_24_188 VPWR VGND sg13g2_decap_4
XFILLER_21_884 VPWR VGND sg13g2_decap_8
XFILLER_4_516 VPWR VGND sg13g2_decap_8
XFILLER_0_722 VPWR VGND sg13g2_decap_8
XFILLER_43_1013 VPWR VGND sg13g2_decap_8
XFILLER_0_799 VPWR VGND sg13g2_decap_8
XFILLER_48_759 VPWR VGND sg13g2_decap_8
XFILLER_29_951 VPWR VGND sg13g2_decap_8
XFILLER_16_634 VPWR VGND sg13g2_decap_8
XFILLER_44_976 VPWR VGND sg13g2_decap_8
XFILLER_43_453 VPWR VGND sg13g2_decap_8
XFILLER_12_840 VPWR VGND sg13g2_decap_8
XFILLER_31_659 VPWR VGND sg13g2_decap_8
XFILLER_8_811 VPWR VGND sg13g2_decap_8
XFILLER_8_888 VPWR VGND sg13g2_decap_8
X_3270_ _1452_ _0713_ _0720_ _0806_ VPWR VGND sg13g2_nor3_1
X_2221_ _1642_ _1633_ net711 net704 _1533_ VPWR VGND sg13g2_a22oi_1
XFILLER_23_4 VPWR VGND sg13g2_fill_1
XFILLER_39_726 VPWR VGND sg13g2_decap_8
X_2152_ net740 net741 _1573_ VPWR VGND sg13g2_nor2b_2
X_2083_ net731 net729 _1504_ VPWR VGND sg13g2_and2_1
XFILLER_19_461 VPWR VGND sg13g2_fill_1
XFILLER_35_954 VPWR VGND sg13g2_decap_8
XFILLER_22_659 VPWR VGND sg13g2_decap_8
X_2985_ _0547_ _0330_ _0538_ VPWR VGND sg13g2_nand2_1
X_3606_ VPWR VGND _1119_ _1070_ _1118_ _1116_ _1120_ _1117_ sg13g2_a221oi_1
X_3537_ net579 VPWR _1061_ VGND net587 _0959_ sg13g2_o21ai_1
XFILLER_27_1019 VPWR VGND sg13g2_decap_8
X_3468_ net559 _0918_ _0944_ _0996_ _0998_ VPWR VGND sg13g2_nor4_1
X_2419_ _1607_ _1662_ _1840_ VPWR VGND _1838_ sg13g2_nand3b_1
X_3399_ _0894_ _0882_ _0916_ _0932_ VPWR VGND sg13g2_a21o_1
XFILLER_38_781 VPWR VGND sg13g2_decap_8
XFILLER_26_954 VPWR VGND sg13g2_decap_8
XFILLER_41_913 VPWR VGND sg13g2_decap_8
XFILLER_25_464 VPWR VGND sg13g2_decap_8
XFILLER_12_125 VPWR VGND sg13g2_fill_1
X_4026__4 VPWR net38 clknet_leaf_2_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_21_681 VPWR VGND sg13g2_decap_8
XFILLER_5_803 VPWR VGND sg13g2_decap_8
XFILLER_0_596 VPWR VGND sg13g2_decap_8
XFILLER_48_556 VPWR VGND sg13g2_decap_8
XFILLER_16_442 VPWR VGND sg13g2_fill_1
XFILLER_44_773 VPWR VGND sg13g2_decap_8
XFILLER_16_464 VPWR VGND sg13g2_fill_2
XFILLER_17_976 VPWR VGND sg13g2_decap_8
XFILLER_32_924 VPWR VGND sg13g2_decap_8
X_2770_ _0198_ _1949_ _0339_ VPWR VGND sg13g2_nor2b_2
XFILLER_8_685 VPWR VGND sg13g2_decap_8
XFILLER_7_162 VPWR VGND sg13g2_fill_2
XFILLER_4_880 VPWR VGND sg13g2_decap_8
Xfanout609 _0721_ net609 VPWR VGND sg13g2_buf_8
X_3322_ net559 _0856_ _0858_ VPWR VGND sg13g2_nor2_1
X_3253_ _0789_ net644 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] net654
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2204_ _1625_ net716 net717 VPWR VGND sg13g2_nand2b_1
X_3184_ _0720_ _0657_ _0670_ VPWR VGND sg13g2_nand2_1
XFILLER_39_523 VPWR VGND sg13g2_decap_8
X_2135_ sap_3_inst.controller.stage\[3\] net717 _1556_ VPWR VGND sg13g2_nor2b_2
XFILLER_27_718 VPWR VGND sg13g2_decap_8
XFILLER_26_228 VPWR VGND sg13g2_fill_1
XFILLER_35_751 VPWR VGND sg13g2_decap_8
X_2066_ VPWR _1489_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_23_913 VPWR VGND sg13g2_decap_8
XFILLER_34_283 VPWR VGND sg13g2_fill_1
XFILLER_10_629 VPWR VGND sg13g2_decap_8
X_2968_ VGND VPWR sap_3_inst.alu.act\[6\] net669 _0531_ net616 sg13g2_a21oi_1
XFILLER_33_1012 VPWR VGND sg13g2_decap_8
X_2899_ _0455_ VPWR _0464_ VGND net564 _0463_ sg13g2_o21ai_1
XFILLER_40_1005 VPWR VGND sg13g2_decap_8
XFILLER_45_548 VPWR VGND sg13g2_decap_8
XFILLER_41_710 VPWR VGND sg13g2_decap_8
XFILLER_26_751 VPWR VGND sg13g2_decap_8
XFILLER_14_957 VPWR VGND sg13g2_decap_8
XFILLER_13_467 VPWR VGND sg13g2_fill_1
XFILLER_41_787 VPWR VGND sg13g2_decap_8
XFILLER_40_297 VPWR VGND sg13g2_decap_4
XFILLER_5_600 VPWR VGND sg13g2_decap_8
XFILLER_4_121 VPWR VGND sg13g2_decap_8
XFILLER_5_677 VPWR VGND sg13g2_decap_8
XFILLER_49_843 VPWR VGND sg13g2_decap_8
XFILLER_48_353 VPWR VGND sg13g2_decap_8
XFILLER_1_1010 VPWR VGND sg13g2_decap_8
XFILLER_17_773 VPWR VGND sg13g2_decap_8
X_3940_ VPWR VGND _1374_ net765 _1369_ _1479_ _1375_ _1310_ sg13g2_a221oi_1
XFILLER_44_570 VPWR VGND sg13g2_decap_8
XFILLER_32_721 VPWR VGND sg13g2_decap_8
X_3871_ sap_3_inst.reg_file.array_serializer_inst.word_index\[3\] sap_3_inst.reg_file.array_serializer_inst.word_index\[2\]
+ _1307_ _1312_ VPWR VGND sg13g2_nor3_2
XFILLER_17_1018 VPWR VGND sg13g2_decap_8
XFILLER_20_905 VPWR VGND sg13g2_decap_8
X_2822_ VGND VPWR net758 _1463_ _0389_ _0357_ sg13g2_a21oi_1
XFILLER_32_798 VPWR VGND sg13g2_decap_8
XFILLER_9_950 VPWR VGND sg13g2_decap_8
X_2753_ _0200_ _0201_ _0322_ VPWR VGND sg13g2_and2_1
XFILLER_8_460 VPWR VGND sg13g2_fill_1
X_2684_ VGND VPWR _1926_ _0275_ _0276_ net690 sg13g2_a21oi_1
X_3305_ _0841_ _0839_ _0840_ _0831_ net586 VPWR VGND sg13g2_a22oi_1
X_3236_ _0772_ net587 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] net592
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3167_ _0643_ VPWR _0703_ VGND _1616_ _0702_ sg13g2_o21ai_1
XFILLER_27_515 VPWR VGND sg13g2_decap_8
X_2118_ _1539_ net737 net736 VPWR VGND sg13g2_nand2b_1
X_3098_ net660 net666 _0634_ VPWR VGND sg13g2_nor2_1
XFILLER_39_397 VPWR VGND sg13g2_fill_2
X_2049_ VPWR _1472_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_23_710 VPWR VGND sg13g2_decap_8
XFILLER_11_949 VPWR VGND sg13g2_decap_8
XFILLER_23_787 VPWR VGND sg13g2_decap_8
XFILLER_7_909 VPWR VGND sg13g2_decap_8
XFILLER_2_658 VPWR VGND sg13g2_decap_8
XFILLER_38_86 VPWR VGND sg13g2_fill_2
XFILLER_46_857 VPWR VGND sg13g2_decap_8
XFILLER_18_537 VPWR VGND sg13g2_decap_8
XFILLER_33_529 VPWR VGND sg13g2_decap_8
XFILLER_14_754 VPWR VGND sg13g2_decap_8
XFILLER_41_584 VPWR VGND sg13g2_decap_8
Xclkload16 clknet_5_18__leaf_sap_3_inst.alu.clk_regs clkload16/X VPWR VGND sg13g2_buf_1
XFILLER_6_953 VPWR VGND sg13g2_decap_8
XFILLER_10_993 VPWR VGND sg13g2_decap_8
XFILLER_5_474 VPWR VGND sg13g2_decap_8
XFILLER_49_640 VPWR VGND sg13g2_decap_8
X_4070_ net789 VGND VPWR _0048_ sap_3_inst.out\[6\] clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_23_1011 VPWR VGND sg13g2_decap_8
X_3021_ _0573_ VPWR _0574_ VGND _0426_ _0570_ sg13g2_o21ai_1
XFILLER_37_835 VPWR VGND sg13g2_decap_8
XFILLER_36_312 VPWR VGND sg13g2_fill_2
XFILLER_17_570 VPWR VGND sg13g2_decap_8
X_3923_ net764 net49 _1359_ _0166_ VPWR VGND sg13g2_a21o_1
X_3854_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[7\] _1291_
+ _1296_ _1295_ sg13g2_a21oi_1
XFILLER_20_702 VPWR VGND sg13g2_decap_8
X_2805_ _1936_ VPWR _0373_ VGND net760 _0372_ sg13g2_o21ai_1
XFILLER_32_595 VPWR VGND sg13g2_decap_8
XFILLER_20_779 VPWR VGND sg13g2_decap_8
XFILLER_30_1004 VPWR VGND sg13g2_decap_8
X_3785_ net600 _1040_ _1041_ _1249_ VPWR VGND sg13g2_nor3_1
X_2736_ _0303_ _0304_ _0300_ _0305_ VPWR VGND sg13g2_nand3_1
X_2667_ VGND VPWR _1812_ _0259_ mem_ram_we _1526_ sg13g2_a21oi_1
X_2598_ VGND VPWR _2007_ _1952_ _1945_ sg13g2_or2_1
XFILLER_28_813 VPWR VGND sg13g2_decap_8
X_3219_ _0755_ net588 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] net657
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_161 VPWR VGND sg13g2_fill_2
X_4199_ net775 VGND VPWR _0177_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\]
+ clknet_5_11__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_15_507 VPWR VGND sg13g2_decap_8
XFILLER_43_838 VPWR VGND sg13g2_decap_8
XFILLER_42_337 VPWR VGND sg13g2_fill_1
XFILLER_23_584 VPWR VGND sg13g2_decap_8
XFILLER_7_706 VPWR VGND sg13g2_decap_8
XFILLER_11_746 VPWR VGND sg13g2_decap_8
XFILLER_24_99 VPWR VGND sg13g2_fill_1
XFILLER_3_934 VPWR VGND sg13g2_decap_8
XFILLER_46_1011 VPWR VGND sg13g2_decap_8
XFILLER_2_455 VPWR VGND sg13g2_decap_8
Xfanout781 net782 net781 VPWR VGND sg13g2_buf_8
XFILLER_19_824 VPWR VGND sg13g2_decap_8
Xfanout770 net772 net770 VPWR VGND sg13g2_buf_8
Xfanout792 net801 net792 VPWR VGND sg13g2_buf_8
XFILLER_46_654 VPWR VGND sg13g2_decap_8
XFILLER_34_816 VPWR VGND sg13g2_decap_8
XFILLER_42_860 VPWR VGND sg13g2_decap_8
XFILLER_14_551 VPWR VGND sg13g2_decap_8
XFILLER_10_790 VPWR VGND sg13g2_decap_8
X_3570_ net589 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] _1088_ _0084_
+ VPWR VGND sg13g2_a21o_1
XFILLER_6_750 VPWR VGND sg13g2_decap_8
X_2521_ net690 _1933_ _1934_ VPWR VGND sg13g2_nor2_1
X_2452_ _1871_ _1869_ _1870_ VPWR VGND sg13g2_nand2_1
X_2383_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] net638
+ net623 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] _1804_ net625 sg13g2_a221oi_1
X_4122_ net773 VGND VPWR _0100_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\]
+ clknet_5_4__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4053_ net787 VGND VPWR _0031_ sap_3_inst.alu.flags\[5\] net45 sg13g2_dfrbpq_1
X_3004_ net754 sap_3_inst.out\[3\] net674 _0045_ VPWR VGND sg13g2_mux2_1
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_37_632 VPWR VGND sg13g2_decap_8
XFILLER_25_849 VPWR VGND sg13g2_decap_8
X_3906_ _1344_ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] _1312_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_893 VPWR VGND sg13g2_decap_8
XFILLER_20_576 VPWR VGND sg13g2_decap_8
X_3837_ _1284_ _1282_ _1283_ VPWR VGND sg13g2_nand2_1
X_3768_ net574 _0955_ _1235_ _1236_ VPWR VGND sg13g2_nor3_1
X_2719_ mem_mar_we _1503_ _0297_ VPWR VGND sg13g2_nand2_1
X_3699_ net22 _1063_ _1065_ _1190_ VPWR VGND sg13g2_nor3_1
XFILLER_0_904 VPWR VGND sg13g2_decap_8
XFILLER_28_610 VPWR VGND sg13g2_decap_8
XFILLER_16_816 VPWR VGND sg13g2_decap_8
XFILLER_43_635 VPWR VGND sg13g2_decap_8
XFILLER_28_687 VPWR VGND sg13g2_decap_8
XFILLER_7_503 VPWR VGND sg13g2_decap_8
XFILLER_11_543 VPWR VGND sg13g2_decap_8
XFILLER_3_731 VPWR VGND sg13g2_decap_8
XFILLER_39_908 VPWR VGND sg13g2_decap_8
XFILLER_47_941 VPWR VGND sg13g2_decap_8
XFILLER_19_621 VPWR VGND sg13g2_decap_8
XFILLER_20_1003 VPWR VGND sg13g2_decap_8
XFILLER_46_451 VPWR VGND sg13g2_decap_8
XFILLER_19_698 VPWR VGND sg13g2_decap_8
XFILLER_34_613 VPWR VGND sg13g2_decap_8
XFILLER_15_871 VPWR VGND sg13g2_decap_8
X_3622_ _1130_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] net551 _0094_
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_885 VPWR VGND sg13g2_decap_8
X_3553_ VPWR _1074_ _1073_ VGND sg13g2_inv_1
X_2504_ VGND VPWR _1723_ _1908_ _1919_ _1918_ sg13g2_a21oi_1
X_3484_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[6\] _1013_ _0717_ _0073_
+ VPWR VGND sg13g2_mux2_1
X_2435_ VGND VPWR _1851_ _1855_ _1856_ net565 sg13g2_a21oi_1
X_2366_ _1776_ _1779_ _1726_ _1787_ VPWR VGND _1785_ sg13g2_nand4_1
X_4105_ net795 VGND VPWR _0083_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\]
+ clknet_5_27__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2297_ _1551_ _1717_ _1718_ VPWR VGND sg13g2_nor2_1
XFILLER_2_80 VPWR VGND sg13g2_fill_1
XFILLER_2_91 VPWR VGND sg13g2_fill_1
X_4036_ net783 VGND VPWR _0018_ u_ser.shadow_reg\[0\] clknet_3_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_38_963 VPWR VGND sg13g2_decap_8
XFILLER_37_473 VPWR VGND sg13g2_decap_4
XFILLER_24_123 VPWR VGND sg13g2_fill_1
XFILLER_25_646 VPWR VGND sg13g2_decap_8
XFILLER_40_627 VPWR VGND sg13g2_decap_8
XFILLER_33_690 VPWR VGND sg13g2_decap_8
XFILLER_21_863 VPWR VGND sg13g2_decap_8
XFILLER_0_701 VPWR VGND sg13g2_decap_8
XFILLER_0_778 VPWR VGND sg13g2_decap_8
XFILLER_48_738 VPWR VGND sg13g2_decap_8
XFILLER_29_930 VPWR VGND sg13g2_decap_8
XFILLER_16_613 VPWR VGND sg13g2_decap_8
XFILLER_28_484 VPWR VGND sg13g2_decap_8
XFILLER_44_955 VPWR VGND sg13g2_decap_8
XFILLER_43_432 VPWR VGND sg13g2_decap_8
XFILLER_15_145 VPWR VGND sg13g2_fill_2
XFILLER_15_178 VPWR VGND sg13g2_fill_1
XFILLER_31_638 VPWR VGND sg13g2_decap_8
XFILLER_12_896 VPWR VGND sg13g2_decap_8
XFILLER_8_867 VPWR VGND sg13g2_decap_8
XFILLER_7_47 VPWR VGND sg13g2_fill_1
X_2220_ net711 _1633_ _1641_ VPWR VGND sg13g2_and2_1
XFILLER_39_705 VPWR VGND sg13g2_decap_8
X_2151_ _1551_ VPWR _1572_ VGND _1569_ _1571_ sg13g2_o21ai_1
X_2082_ _1503_ _1499_ net715 VPWR VGND sg13g2_nand2_1
XFILLER_35_933 VPWR VGND sg13g2_decap_8
XFILLER_19_495 VPWR VGND sg13g2_decap_8
X_2984_ _0546_ _0540_ _0333_ net573 net746 VPWR VGND sg13g2_a22oi_1
XFILLER_22_638 VPWR VGND sg13g2_decap_8
XFILLER_30_682 VPWR VGND sg13g2_decap_8
X_3605_ _1119_ _1078_ net15 VPWR VGND sg13g2_nand2b_1
X_3536_ _0953_ _1059_ _1060_ VPWR VGND sg13g2_nor2_1
X_3467_ _0918_ net552 _0996_ _0997_ VPWR VGND sg13g2_nor3_1
X_2418_ _1554_ _1675_ _1839_ VPWR VGND sg13g2_nor2_1
X_3398_ _0825_ _0881_ net553 _0931_ VPWR VGND _0930_ sg13g2_nand4_1
X_2349_ _1765_ _1769_ _1770_ VPWR VGND net681 sg13g2_nand3b_1
X_4019_ net767 _1410_ _1429_ VPWR VGND sg13g2_nor2_1
XFILLER_26_933 VPWR VGND sg13g2_decap_8
XFILLER_38_760 VPWR VGND sg13g2_decap_8
XFILLER_25_443 VPWR VGND sg13g2_decap_8
XFILLER_13_649 VPWR VGND sg13g2_decap_8
XFILLER_41_969 VPWR VGND sg13g2_decap_8
XFILLER_8_108 VPWR VGND sg13g2_fill_2
XFILLER_21_660 VPWR VGND sg13g2_decap_8
XFILLER_5_859 VPWR VGND sg13g2_decap_8
XFILLER_48_535 VPWR VGND sg13g2_decap_8
XFILLER_0_575 VPWR VGND sg13g2_decap_8
XFILLER_17_955 VPWR VGND sg13g2_decap_8
XFILLER_44_752 VPWR VGND sg13g2_decap_8
XFILLER_32_903 VPWR VGND sg13g2_decap_8
XFILLER_31_413 VPWR VGND sg13g2_fill_2
XFILLER_40_991 VPWR VGND sg13g2_decap_8
XFILLER_8_664 VPWR VGND sg13g2_decap_8
XFILLER_12_693 VPWR VGND sg13g2_decap_8
X_3321_ _0744_ net553 _0757_ _0857_ VGND VPWR _0854_ sg13g2_nor4_2
XFILLER_3_380 VPWR VGND sg13g2_fill_1
X_3252_ _0777_ _0778_ _0781_ _0786_ _0788_ VPWR VGND sg13g2_or4_1
XFILLER_39_502 VPWR VGND sg13g2_decap_8
X_2203_ net717 net716 _1624_ VPWR VGND sg13g2_nor2b_1
X_3183_ _0658_ net665 _0719_ VPWR VGND sg13g2_nor2_2
X_2134_ net735 net723 _1509_ _1555_ VGND VPWR _1521_ sg13g2_nor4_2
XFILLER_39_579 VPWR VGND sg13g2_decap_8
XFILLER_35_730 VPWR VGND sg13g2_decap_8
X_2065_ VPWR _1488_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_10_608 VPWR VGND sg13g2_decap_8
XFILLER_23_969 VPWR VGND sg13g2_decap_8
X_2967_ _0530_ _0528_ _0529_ VPWR VGND sg13g2_nand2_1
X_2898_ _0458_ _0432_ _0463_ VPWR VGND sg13g2_xor2_1
X_3519_ VGND VPWR _1046_ _1043_ net32 sg13g2_or2_1
XFILLER_40_1028 VPWR VGND sg13g2_fill_1
XFILLER_45_527 VPWR VGND sg13g2_decap_8
XFILLER_18_719 VPWR VGND sg13g2_decap_8
XFILLER_27_22 VPWR VGND sg13g2_fill_2
XFILLER_26_730 VPWR VGND sg13g2_decap_8
XFILLER_13_424 VPWR VGND sg13g2_fill_1
XFILLER_14_936 VPWR VGND sg13g2_decap_8
XFILLER_41_766 VPWR VGND sg13g2_decap_8
XFILLER_40_276 VPWR VGND sg13g2_fill_1
XFILLER_5_656 VPWR VGND sg13g2_decap_8
XFILLER_49_822 VPWR VGND sg13g2_decap_8
XFILLER_1_884 VPWR VGND sg13g2_decap_8
XFILLER_48_332 VPWR VGND sg13g2_decap_8
XFILLER_49_899 VPWR VGND sg13g2_decap_8
XFILLER_36_549 VPWR VGND sg13g2_decap_8
XFILLER_17_752 VPWR VGND sg13g2_decap_8
XFILLER_32_700 VPWR VGND sg13g2_decap_8
X_3870_ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\] net768 _1303_ _1311_
+ VPWR VGND sg13g2_nor3_2
X_2821_ _0388_ _0366_ _0386_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_777 VPWR VGND sg13g2_decap_8
X_2752_ sap_3_inst.alu.tmp\[0\] net759 _0321_ VPWR VGND sg13g2_xor2_1
X_2683_ VPWR VGND _1555_ _1569_ _1690_ net688 _0275_ _1568_ sg13g2_a221oi_1
X_3304_ VGND VPWR net9 _0838_ _0840_ net584 sg13g2_a21oi_1
X_3235_ _0771_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] net640 VPWR
+ VGND sg13g2_nand2_1
XFILLER_39_332 VPWR VGND sg13g2_fill_2
X_3166_ net734 VPWR _0702_ VGND _1638_ _1641_ sg13g2_o21ai_1
X_2117_ _1538_ net712 net694 VPWR VGND sg13g2_nand2_2
X_3097_ net666 _0633_ VPWR VGND sg13g2_inv_4
X_2048_ VPWR _1471_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_23_766 VPWR VGND sg13g2_decap_8
X_3999_ _1415_ net767 u_ser.shadow_reg\[6\] VPWR VGND sg13g2_nand2b_1
XFILLER_11_928 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_fill_1
XFILLER_22_298 VPWR VGND sg13g2_fill_2
XFILLER_2_637 VPWR VGND sg13g2_decap_8
Xclkbuf_5_4__f_sap_3_inst.alu.clk_regs clknet_4_2_0_sap_3_inst.alu.clk_regs clknet_5_4__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_18_516 VPWR VGND sg13g2_decap_8
XFILLER_38_65 VPWR VGND sg13g2_fill_2
XFILLER_38_76 VPWR VGND sg13g2_fill_2
XFILLER_46_836 VPWR VGND sg13g2_decap_8
XFILLER_33_508 VPWR VGND sg13g2_decap_8
XFILLER_14_733 VPWR VGND sg13g2_decap_8
XFILLER_41_563 VPWR VGND sg13g2_decap_8
XFILLER_9_214 VPWR VGND sg13g2_fill_1
XFILLER_9_203 VPWR VGND sg13g2_fill_2
Xclkload17 VPWR clkload17/Y clknet_5_21__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
XFILLER_10_972 VPWR VGND sg13g2_decap_8
XFILLER_6_932 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_1_681 VPWR VGND sg13g2_decap_8
X_3020_ VPWR VGND _0538_ _0571_ _0572_ _0449_ _0573_ _0569_ sg13g2_a221oi_1
XFILLER_37_814 VPWR VGND sg13g2_decap_8
XFILLER_49_696 VPWR VGND sg13g2_decap_8
XFILLER_24_519 VPWR VGND sg13g2_decap_8
XFILLER_36_368 VPWR VGND sg13g2_fill_2
XFILLER_45_891 VPWR VGND sg13g2_decap_8
X_3922_ VPWR VGND _1358_ net765 _1353_ _1468_ _1359_ net763 sg13g2_a221oi_1
X_3853_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\] VPWR _1295_ VGND sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\]
+ _1294_ sg13g2_o21ai_1
XFILLER_32_574 VPWR VGND sg13g2_decap_8
X_2804_ _0370_ _0371_ _0372_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_758 VPWR VGND sg13g2_decap_8
X_3784_ _0138_ _1247_ _1248_ net598 _1493_ VPWR VGND sg13g2_a22oi_1
X_2735_ _0301_ _1832_ _0304_ VPWR VGND sg13g2_nor2b_1
X_2666_ _1823_ VPWR _0259_ VGND _1816_ _0258_ sg13g2_o21ai_1
X_2597_ _1978_ VPWR _0028_ VGND _1998_ _2006_ sg13g2_o21ai_1
Xclkbuf_5_11__f_sap_3_inst.alu.clk_regs clknet_4_5_0_sap_3_inst.alu.clk_regs clknet_5_11__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
X_3218_ _0754_ net593 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] net641
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] VPWR VGND sg13g2_a22oi_1
X_4198_ net780 VGND VPWR _0176_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\]
+ clknet_5_30__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3149_ _1786_ _0684_ _0685_ VPWR VGND sg13g2_nor2_1
XFILLER_43_817 VPWR VGND sg13g2_decap_8
XFILLER_28_869 VPWR VGND sg13g2_decap_8
XFILLER_11_725 VPWR VGND sg13g2_decap_8
XFILLER_23_563 VPWR VGND sg13g2_decap_8
XFILLER_10_213 VPWR VGND sg13g2_fill_2
XFILLER_3_913 VPWR VGND sg13g2_decap_8
Xfanout760 sap_3_inst.alu.acc\[0\] net760 VPWR VGND sg13g2_buf_8
XFILLER_19_803 VPWR VGND sg13g2_decap_8
Xfanout771 net772 net771 VPWR VGND sg13g2_buf_2
Xfanout782 net801 net782 VPWR VGND sg13g2_buf_8
Xfanout793 net798 net793 VPWR VGND sg13g2_buf_8
XFILLER_46_633 VPWR VGND sg13g2_decap_8
XFILLER_33_305 VPWR VGND sg13g2_fill_1
XFILLER_14_530 VPWR VGND sg13g2_decap_8
X_2520_ VGND VPWR net706 _1932_ _1933_ _1715_ sg13g2_a21oi_1
X_2451_ _1870_ net623 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] _1795_
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2382_ net662 _1761_ _1773_ _1803_ VPWR VGND sg13g2_nor3_2
X_4121_ net795 VGND VPWR _0099_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\]
+ clknet_5_26__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4052_ net787 VGND VPWR _0030_ sap_3_inst.alu.flags\[4\] net44 sg13g2_dfrbpq_1
XFILLER_49_493 VPWR VGND sg13g2_decap_8
X_3003_ net756 sap_3_inst.out\[2\] net673 _0044_ VPWR VGND sg13g2_mux2_1
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
XFILLER_36_110 VPWR VGND sg13g2_fill_1
XFILLER_37_611 VPWR VGND sg13g2_decap_8
XFILLER_18_880 VPWR VGND sg13g2_decap_8
XFILLER_25_828 VPWR VGND sg13g2_decap_8
XFILLER_37_688 VPWR VGND sg13g2_decap_8
XFILLER_40_809 VPWR VGND sg13g2_decap_8
X_3905_ net764 net54 _1343_ _0164_ VPWR VGND sg13g2_a21o_1
XFILLER_33_872 VPWR VGND sg13g2_decap_8
X_4033__11 VPWR net45 clknet_leaf_1_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_20_555 VPWR VGND sg13g2_decap_8
X_3836_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\] net769 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[2\]
+ _1283_ VPWR VGND sg13g2_nand3_1
X_3767_ _0918_ net552 _1235_ VPWR VGND sg13g2_and2_1
X_2718_ _0297_ _1537_ _0296_ VPWR VGND sg13g2_nand2_1
X_3698_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] _1182_ _1189_ VPWR
+ VGND sg13g2_nor2_1
X_2649_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] _1802_
+ net633 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] _0244_ net635 sg13g2_a221oi_1
XFILLER_27_121 VPWR VGND sg13g2_fill_2
XFILLER_28_666 VPWR VGND sg13g2_decap_8
XFILLER_43_614 VPWR VGND sg13g2_decap_8
XFILLER_27_187 VPWR VGND sg13g2_fill_1
XFILLER_27_198 VPWR VGND sg13g2_fill_2
XFILLER_24_883 VPWR VGND sg13g2_decap_8
XFILLER_35_88 VPWR VGND sg13g2_fill_1
XFILLER_11_522 VPWR VGND sg13g2_decap_8
XFILLER_11_599 VPWR VGND sg13g2_decap_8
XFILLER_7_559 VPWR VGND sg13g2_decap_8
XFILLER_3_710 VPWR VGND sg13g2_decap_8
XFILLER_3_787 VPWR VGND sg13g2_decap_8
XFILLER_19_600 VPWR VGND sg13g2_decap_8
XFILLER_47_920 VPWR VGND sg13g2_decap_8
Xfanout590 net591 net590 VPWR VGND sg13g2_buf_8
XFILLER_46_430 VPWR VGND sg13g2_decap_8
XFILLER_47_997 VPWR VGND sg13g2_decap_8
XFILLER_19_677 VPWR VGND sg13g2_decap_8
XFILLER_34_669 VPWR VGND sg13g2_decap_8
XFILLER_15_850 VPWR VGND sg13g2_decap_8
Xclkbuf_1_0__f_sap_3_inst.alu.clk clknet_0_sap_3_inst.alu.clk clknet_1_0__leaf_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_33_168 VPWR VGND sg13g2_fill_2
XFILLER_30_864 VPWR VGND sg13g2_decap_8
X_3621_ _1129_ net546 _1130_ VPWR VGND _1052_ sg13g2_nand3b_1
X_3552_ _1073_ net585 _1028_ VPWR VGND sg13g2_nand2_1
X_2503_ VGND VPWR _1913_ _1917_ _1918_ net565 sg13g2_a21oi_1
X_3483_ _1010_ _1012_ _1004_ _1013_ VPWR VGND sg13g2_nand3_1
X_2434_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] _1854_
+ net623 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] _1855_ net629 sg13g2_a221oi_1
X_2365_ _1554_ _1559_ _1786_ VPWR VGND sg13g2_nor2_1
X_4104_ net775 VGND VPWR _0082_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\]
+ clknet_5_3__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2296_ net698 _1716_ _1717_ VPWR VGND sg13g2_and2_1
XFILLER_38_942 VPWR VGND sg13g2_decap_8
XFILLER_25_625 VPWR VGND sg13g2_decap_8
XFILLER_40_606 VPWR VGND sg13g2_decap_8
XFILLER_36_1011 VPWR VGND sg13g2_decap_8
XFILLER_21_842 VPWR VGND sg13g2_decap_8
X_3819_ _1270_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] net602 VPWR
+ VGND sg13g2_nand2_1
XFILLER_48_717 VPWR VGND sg13g2_decap_8
XFILLER_0_757 VPWR VGND sg13g2_decap_8
XFILLER_47_216 VPWR VGND sg13g2_fill_1
XFILLER_46_76 VPWR VGND sg13g2_fill_1
XFILLER_44_934 VPWR VGND sg13g2_decap_8
XFILLER_28_463 VPWR VGND sg13g2_decap_8
XFILLER_29_986 VPWR VGND sg13g2_decap_8
XFILLER_43_411 VPWR VGND sg13g2_decap_8
XFILLER_15_168 VPWR VGND sg13g2_fill_2
XFILLER_16_669 VPWR VGND sg13g2_decap_8
XFILLER_31_617 VPWR VGND sg13g2_decap_8
XFILLER_43_488 VPWR VGND sg13g2_decap_8
XFILLER_24_680 VPWR VGND sg13g2_decap_8
XFILLER_8_846 VPWR VGND sg13g2_decap_8
XFILLER_12_875 VPWR VGND sg13g2_decap_8
XFILLER_7_334 VPWR VGND sg13g2_fill_2
XFILLER_3_584 VPWR VGND sg13g2_decap_8
X_2150_ _1571_ _1560_ _1570_ VPWR VGND sg13g2_nand2_1
X_2081_ net718 _1500_ _1502_ VPWR VGND sg13g2_nor2_1
XFILLER_4_1020 VPWR VGND sg13g2_decap_8
XFILLER_35_912 VPWR VGND sg13g2_decap_8
XFILLER_47_794 VPWR VGND sg13g2_decap_8
XFILLER_22_617 VPWR VGND sg13g2_decap_8
XFILLER_35_989 VPWR VGND sg13g2_decap_8
X_2983_ _0545_ _0340_ _0539_ net572 _0337_ VPWR VGND sg13g2_a22oi_1
XFILLER_30_661 VPWR VGND sg13g2_decap_8
X_3604_ _1118_ net547 _1077_ VPWR VGND sg13g2_nand2_1
X_3535_ _0947_ net584 net21 _1059_ VPWR VGND sg13g2_a21o_2
X_3466_ _0996_ _0969_ _0994_ VPWR VGND sg13g2_nand2_1
X_2417_ _1576_ net686 _1838_ VPWR VGND sg13g2_nor2_1
X_3397_ _0894_ _0916_ _0930_ VPWR VGND sg13g2_and2_1
X_2348_ _1664_ _1732_ _1766_ _1768_ _1769_ VPWR VGND sg13g2_nor4_1
XFILLER_45_709 VPWR VGND sg13g2_decap_8
X_2279_ VPWR _1700_ _1699_ VGND sg13g2_inv_1
XFILLER_29_249 VPWR VGND sg13g2_fill_2
X_4018_ VPWR _0193_ _1428_ VGND sg13g2_inv_1
XFILLER_26_912 VPWR VGND sg13g2_decap_8
XFILLER_25_422 VPWR VGND sg13g2_decap_8
XFILLER_26_989 VPWR VGND sg13g2_decap_8
XFILLER_41_948 VPWR VGND sg13g2_decap_8
XFILLER_13_628 VPWR VGND sg13g2_decap_8
XFILLER_25_499 VPWR VGND sg13g2_decap_8
XFILLER_12_149 VPWR VGND sg13g2_fill_2
XFILLER_5_838 VPWR VGND sg13g2_decap_8
XFILLER_10_1014 VPWR VGND sg13g2_decap_8
XFILLER_4_337 VPWR VGND sg13g2_fill_1
XFILLER_0_554 VPWR VGND sg13g2_decap_8
Xclkbuf_4_14_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_14_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_48_514 VPWR VGND sg13g2_decap_8
XFILLER_29_783 VPWR VGND sg13g2_decap_8
XFILLER_44_731 VPWR VGND sg13g2_decap_8
XFILLER_17_934 VPWR VGND sg13g2_decap_8
XFILLER_32_959 VPWR VGND sg13g2_decap_8
XFILLER_40_970 VPWR VGND sg13g2_decap_8
XFILLER_12_672 VPWR VGND sg13g2_decap_8
XFILLER_8_643 VPWR VGND sg13g2_decap_8
XFILLER_11_182 VPWR VGND sg13g2_fill_1
XFILLER_7_164 VPWR VGND sg13g2_fill_1
X_3320_ VGND VPWR _0856_ _0855_ net553 sg13g2_or2_1
XFILLER_26_1010 VPWR VGND sg13g2_decap_8
X_3251_ _0777_ _0778_ _0781_ _0787_ VGND VPWR _0786_ sg13g2_nor4_2
X_2202_ _1623_ net700 _1622_ VPWR VGND sg13g2_nand2_2
X_3182_ _0718_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[0\] _0716_ VPWR
+ VGND sg13g2_nand2_1
X_2133_ _1554_ _1520_ VPWR VGND _1509_ sg13g2_nand2b_2
XFILLER_39_558 VPWR VGND sg13g2_decap_8
XFILLER_47_591 VPWR VGND sg13g2_decap_8
X_2064_ VPWR _1487_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_23_948 VPWR VGND sg13g2_decap_8
XFILLER_35_786 VPWR VGND sg13g2_decap_8
X_2966_ VGND VPWR _0504_ _0527_ _0529_ net670 sg13g2_a21oi_1
XFILLER_31_981 VPWR VGND sg13g2_decap_8
X_2897_ _0462_ _0460_ _0461_ VPWR VGND sg13g2_nand2_1
XFILLER_2_819 VPWR VGND sg13g2_decap_8
X_3518_ net660 _1044_ _1045_ VPWR VGND sg13g2_nor2b_1
X_3449_ net661 _0979_ _0980_ VPWR VGND sg13g2_nor2b_1
XFILLER_45_506 VPWR VGND sg13g2_decap_8
XFILLER_14_915 VPWR VGND sg13g2_decap_8
Xclkbuf_4_6_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_6_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_26_786 VPWR VGND sg13g2_decap_8
XFILLER_41_745 VPWR VGND sg13g2_decap_8
XFILLER_13_458 VPWR VGND sg13g2_fill_1
XFILLER_9_429 VPWR VGND sg13g2_fill_2
XFILLER_22_981 VPWR VGND sg13g2_decap_8
XFILLER_5_635 VPWR VGND sg13g2_decap_8
XFILLER_4_167 VPWR VGND sg13g2_fill_2
XFILLER_49_801 VPWR VGND sg13g2_decap_8
XFILLER_1_863 VPWR VGND sg13g2_decap_8
XFILLER_49_878 VPWR VGND sg13g2_decap_8
XFILLER_48_388 VPWR VGND sg13g2_decap_8
XFILLER_17_731 VPWR VGND sg13g2_decap_8
XFILLER_29_580 VPWR VGND sg13g2_decap_8
XFILLER_36_528 VPWR VGND sg13g2_decap_8
XFILLER_31_233 VPWR VGND sg13g2_fill_1
XFILLER_32_756 VPWR VGND sg13g2_decap_8
X_2820_ VPWR _0387_ _0386_ VGND sg13g2_inv_1
X_2751_ _0320_ net759 sap_3_inst.alu.tmp\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_13_992 VPWR VGND sg13g2_decap_8
X_2682_ _0264_ _0272_ _1815_ _0274_ VPWR VGND sg13g2_nand3_1
XFILLER_9_985 VPWR VGND sg13g2_decap_8
X_3303_ _0839_ net31 net571 VPWR VGND sg13g2_nand2_1
X_3234_ _0770_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] net613 VPWR
+ VGND sg13g2_nand2_1
X_3165_ _0699_ _0700_ _0698_ _0701_ VPWR VGND sg13g2_nand3_1
X_3096_ _0631_ VPWR _0632_ VGND _1651_ _0626_ sg13g2_o21ai_1
X_2116_ VPWR VGND _1499_ _1526_ _1536_ net713 _1537_ net694 sg13g2_a221oi_1
X_2047_ VPWR _1470_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_35_583 VPWR VGND sg13g2_decap_8
XFILLER_11_907 VPWR VGND sg13g2_decap_8
XFILLER_23_745 VPWR VGND sg13g2_decap_8
X_3998_ u_ser.shadow_reg\[7\] u_ser.bit_pos\[1\] _1414_ VPWR VGND net767 sg13g2_nand3b_1
X_2949_ VGND VPWR _0512_ _0510_ _0482_ sg13g2_or2_1
XFILLER_2_616 VPWR VGND sg13g2_decap_8
XFILLER_46_815 VPWR VGND sg13g2_decap_8
XFILLER_38_88 VPWR VGND sg13g2_fill_1
XFILLER_14_712 VPWR VGND sg13g2_decap_8
XFILLER_26_583 VPWR VGND sg13g2_decap_8
XFILLER_41_542 VPWR VGND sg13g2_decap_8
XFILLER_14_789 VPWR VGND sg13g2_decap_8
XFILLER_6_911 VPWR VGND sg13g2_decap_8
XFILLER_10_951 VPWR VGND sg13g2_decap_8
Xclkload18 clknet_5_23__leaf_sap_3_inst.alu.clk_regs clkload18/X VPWR VGND sg13g2_buf_1
XFILLER_6_988 VPWR VGND sg13g2_decap_8
XFILLER_1_660 VPWR VGND sg13g2_decap_8
XFILLER_49_675 VPWR VGND sg13g2_decap_8
XFILLER_45_870 VPWR VGND sg13g2_decap_8
XFILLER_44_380 VPWR VGND sg13g2_fill_2
X_3921_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] _1357_
+ _1313_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] _1358_ _1306_ sg13g2_a221oi_1
X_3852_ _1293_ VPWR _1294_ VGND net769 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[5\]
+ sg13g2_o21ai_1
XFILLER_32_553 VPWR VGND sg13g2_decap_8
X_2803_ _1455_ VPWR _0371_ VGND _1550_ _1747_ sg13g2_o21ai_1
XFILLER_20_737 VPWR VGND sg13g2_decap_8
X_3783_ net655 _1125_ _1248_ VPWR VGND sg13g2_and2_1
X_2734_ VGND VPWR _1690_ _0302_ _0303_ _1837_ sg13g2_a21oi_1
XFILLER_9_782 VPWR VGND sg13g2_decap_8
X_2665_ _1699_ net682 _1686_ _0258_ VPWR VGND _0257_ sg13g2_nand4_1
X_2596_ _1955_ VPWR _2006_ VGND net675 _2005_ sg13g2_o21ai_1
XFILLER_8_1007 VPWR VGND sg13g2_decap_8
X_4197_ net779 VGND VPWR _0175_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\]
+ clknet_5_14__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3217_ _0753_ net646 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] _0729_
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] VPWR VGND sg13g2_a22oi_1
X_3148_ VGND VPWR _1593_ _1662_ _0684_ _1703_ sg13g2_a21oi_1
XFILLER_28_848 VPWR VGND sg13g2_decap_8
XFILLER_42_317 VPWR VGND sg13g2_fill_2
X_3079_ _0615_ _1589_ _1932_ VPWR VGND sg13g2_nand2_1
XFILLER_39_1020 VPWR VGND sg13g2_decap_8
XFILLER_23_542 VPWR VGND sg13g2_decap_8
XFILLER_36_892 VPWR VGND sg13g2_decap_8
XFILLER_11_704 VPWR VGND sg13g2_decap_8
XFILLER_40_89 VPWR VGND sg13g2_fill_2
XFILLER_49_21 VPWR VGND sg13g2_fill_2
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_3_969 VPWR VGND sg13g2_decap_8
Xfanout750 net751 net750 VPWR VGND sg13g2_buf_8
Xfanout761 _1315_ net761 VPWR VGND sg13g2_buf_8
Xfanout783 net785 net783 VPWR VGND sg13g2_buf_8
Xfanout772 net773 net772 VPWR VGND sg13g2_buf_8
Xfanout794 net798 net794 VPWR VGND sg13g2_buf_1
XFILLER_46_612 VPWR VGND sg13g2_decap_8
XFILLER_1_39 VPWR VGND sg13g2_decap_4
XFILLER_19_859 VPWR VGND sg13g2_decap_8
XFILLER_46_689 VPWR VGND sg13g2_decap_8
XFILLER_26_380 VPWR VGND sg13g2_decap_8
XFILLER_42_895 VPWR VGND sg13g2_decap_8
XFILLER_14_586 VPWR VGND sg13g2_decap_8
XFILLER_6_785 VPWR VGND sg13g2_decap_8
X_2450_ _1869_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] _1796_
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2381_ _1802_ net662 _1761_ _1772_ VPWR VGND sg13g2_and3_2
X_4120_ net775 VGND VPWR _0098_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\]
+ clknet_5_11__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_2_980 VPWR VGND sg13g2_decap_8
X_4051_ net772 VGND VPWR _0005_ sap_3_inst.controller.stage\[3\] net43 sg13g2_dfrbpq_2
XFILLER_49_472 VPWR VGND sg13g2_decap_8
X_3002_ _0561_ VPWR _0043_ VGND _1455_ net673 sg13g2_o21ai_1
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
XFILLER_25_807 VPWR VGND sg13g2_decap_8
XFILLER_37_667 VPWR VGND sg13g2_decap_8
XFILLER_24_317 VPWR VGND sg13g2_fill_1
X_3904_ VPWR VGND _1342_ net765 _1336_ _1444_ _1343_ net762 sg13g2_a221oi_1
XFILLER_33_851 VPWR VGND sg13g2_decap_8
XFILLER_20_534 VPWR VGND sg13g2_decap_8
X_3835_ sap_3_inst.reg_file.array_serializer_inst.state\[0\] sap_3_inst.reg_file.array_serializer_inst.state\[1\]
+ _1282_ VPWR VGND sg13g2_nor2b_2
X_3766_ VGND VPWR _1441_ net600 _0134_ _1234_ sg13g2_a21oi_1
X_2717_ _0296_ net703 _0295_ VPWR VGND sg13g2_nand2_1
X_3697_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] _1188_ _1182_ _0111_
+ VPWR VGND sg13g2_mux2_1
XFILLER_10_48 VPWR VGND sg13g2_fill_1
X_2648_ _0243_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] net639
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_0_939 VPWR VGND sg13g2_decap_8
X_2579_ _1990_ net626 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] net630
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_47_409 VPWR VGND sg13g2_decap_8
XFILLER_28_645 VPWR VGND sg13g2_decap_8
XFILLER_24_862 VPWR VGND sg13g2_decap_8
XFILLER_11_501 VPWR VGND sg13g2_decap_8
XFILLER_23_383 VPWR VGND sg13g2_decap_4
XFILLER_7_538 VPWR VGND sg13g2_decap_8
XFILLER_11_578 VPWR VGND sg13g2_decap_8
XFILLER_3_766 VPWR VGND sg13g2_decap_8
Xfanout591 _0739_ net591 VPWR VGND sg13g2_buf_8
Xfanout580 net582 net580 VPWR VGND sg13g2_buf_8
XFILLER_47_976 VPWR VGND sg13g2_decap_8
XFILLER_18_133 VPWR VGND sg13g2_fill_1
XFILLER_19_656 VPWR VGND sg13g2_decap_8
XFILLER_46_486 VPWR VGND sg13g2_decap_8
XFILLER_34_648 VPWR VGND sg13g2_decap_8
XFILLER_42_692 VPWR VGND sg13g2_decap_8
XFILLER_30_843 VPWR VGND sg13g2_decap_8
X_3620_ _1129_ net580 _0924_ VPWR VGND sg13g2_nand2_1
X_3551_ VGND VPWR _1489_ net558 _0081_ _1072_ sg13g2_a21oi_1
X_2502_ _1917_ _1914_ _1915_ _1916_ VPWR VGND sg13g2_and3_1
XFILLER_6_582 VPWR VGND sg13g2_decap_8
X_3482_ _1011_ VPWR _1012_ VGND net15 net571 sg13g2_o21ai_1
X_2433_ _1852_ _1853_ _1850_ _1854_ VPWR VGND sg13g2_nand3_1
X_2364_ _1699_ net682 _1780_ _1784_ _1785_ VPWR VGND sg13g2_and4_1
X_4103_ net797 VGND VPWR _0081_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\]
+ clknet_5_31__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2295_ _1716_ net734 _1504_ VPWR VGND sg13g2_nand2_2
XFILLER_38_921 VPWR VGND sg13g2_decap_8
XFILLER_49_291 VPWR VGND sg13g2_decap_8
XFILLER_25_604 VPWR VGND sg13g2_decap_8
XFILLER_38_998 VPWR VGND sg13g2_decap_8
XFILLER_24_147 VPWR VGND sg13g2_fill_2
XFILLER_21_821 VPWR VGND sg13g2_decap_8
XFILLER_21_898 VPWR VGND sg13g2_decap_8
X_3818_ _0151_ _1103_ _1269_ net603 _1469_ VPWR VGND sg13g2_a22oi_1
X_3749_ net9 net581 _1039_ _1221_ VPWR VGND sg13g2_nor3_1
XFILLER_0_736 VPWR VGND sg13g2_decap_8
XFILLER_43_1027 VPWR VGND sg13g2_fill_2
XFILLER_28_442 VPWR VGND sg13g2_decap_8
XFILLER_29_965 VPWR VGND sg13g2_decap_8
XFILLER_44_913 VPWR VGND sg13g2_decap_8
XFILLER_16_648 VPWR VGND sg13g2_decap_8
XFILLER_43_467 VPWR VGND sg13g2_decap_8
XFILLER_15_147 VPWR VGND sg13g2_fill_1
XFILLER_30_128 VPWR VGND sg13g2_fill_2
XFILLER_12_854 VPWR VGND sg13g2_decap_8
XFILLER_8_825 VPWR VGND sg13g2_decap_8
XFILLER_7_16 VPWR VGND sg13g2_fill_2
XFILLER_3_563 VPWR VGND sg13g2_decap_8
X_2080_ net719 net718 _1501_ VPWR VGND sg13g2_nor2_1
XFILLER_47_773 VPWR VGND sg13g2_decap_8
XFILLER_35_968 VPWR VGND sg13g2_decap_8
X_2982_ _0544_ _0511_ _0542_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_640 VPWR VGND sg13g2_decap_8
X_3603_ net586 _1006_ _1117_ VPWR VGND sg13g2_and2_1
X_3534_ _1058_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] net558 VPWR
+ VGND sg13g2_nand2_1
X_3465_ VPWR _0995_ _0994_ VGND sg13g2_inv_1
X_2416_ _1837_ net736 _1655_ _1690_ VPWR VGND sg13g2_and3_1
X_3396_ _0928_ _0851_ net580 _0929_ VPWR VGND sg13g2_a21o_2
X_2347_ _1768_ _1658_ _1767_ _1606_ _1604_ VPWR VGND sg13g2_a22oi_1
X_2278_ _1699_ _1555_ _1577_ VPWR VGND sg13g2_nand2_2
X_4017_ _1428_ _1425_ net78 _1424_ net721 VPWR VGND sg13g2_a22oi_1
XFILLER_25_401 VPWR VGND sg13g2_decap_8
XFILLER_38_795 VPWR VGND sg13g2_decap_8
XFILLER_13_607 VPWR VGND sg13g2_decap_8
XFILLER_16_58 VPWR VGND sg13g2_fill_1
XFILLER_26_968 VPWR VGND sg13g2_decap_8
XFILLER_41_927 VPWR VGND sg13g2_decap_8
XFILLER_25_478 VPWR VGND sg13g2_decap_8
XFILLER_40_459 VPWR VGND sg13g2_decap_8
XFILLER_21_695 VPWR VGND sg13g2_decap_8
XFILLER_5_817 VPWR VGND sg13g2_decap_8
XFILLER_0_533 VPWR VGND sg13g2_decap_8
XFILLER_17_913 VPWR VGND sg13g2_decap_8
XFILLER_29_762 VPWR VGND sg13g2_decap_8
XFILLER_44_710 VPWR VGND sg13g2_decap_8
XFILLER_16_412 VPWR VGND sg13g2_fill_1
XFILLER_44_787 VPWR VGND sg13g2_decap_8
XFILLER_32_938 VPWR VGND sg13g2_decap_8
XFILLER_8_622 VPWR VGND sg13g2_decap_8
XFILLER_12_651 VPWR VGND sg13g2_decap_8
XFILLER_8_699 VPWR VGND sg13g2_decap_8
XFILLER_4_894 VPWR VGND sg13g2_decap_8
X_3250_ _0783_ _0784_ _0782_ _0786_ VPWR VGND _0785_ sg13g2_nand4_1
X_2201_ _1622_ net735 _1621_ VPWR VGND sg13g2_xnor2_1
X_3181_ _0716_ _0717_ VPWR VGND sg13g2_inv_4
X_2132_ _1509_ _1521_ _1553_ VPWR VGND sg13g2_nor2_2
XFILLER_39_537 VPWR VGND sg13g2_decap_8
XFILLER_47_570 VPWR VGND sg13g2_decap_8
X_2063_ VPWR _1486_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_34_242 VPWR VGND sg13g2_fill_2
XFILLER_35_765 VPWR VGND sg13g2_decap_8
XFILLER_23_927 VPWR VGND sg13g2_decap_8
X_2965_ _0528_ net543 _0516_ VPWR VGND sg13g2_nand2_1
XFILLER_31_960 VPWR VGND sg13g2_decap_8
XFILLER_33_1026 VPWR VGND sg13g2_fill_2
X_2896_ VPWR VGND _0333_ _0446_ _0447_ sap_3_inst.alu.acc\[3\] _0461_ net573 sg13g2_a221oi_1
X_3517_ net586 VPWR _1044_ VGND net655 _0876_ sg13g2_o21ai_1
X_3448_ _0978_ VPWR _0979_ VGND _1899_ _0838_ sg13g2_o21ai_1
X_3379_ _0912_ net648 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] net653
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_40_1019 VPWR VGND sg13g2_decap_8
XFILLER_38_592 VPWR VGND sg13g2_decap_8
XFILLER_26_765 VPWR VGND sg13g2_decap_8
XFILLER_27_79 VPWR VGND sg13g2_fill_2
XFILLER_41_724 VPWR VGND sg13g2_decap_8
XFILLER_22_960 VPWR VGND sg13g2_decap_8
XFILLER_5_614 VPWR VGND sg13g2_decap_8
XFILLER_21_492 VPWR VGND sg13g2_decap_8
XFILLER_49_1011 VPWR VGND sg13g2_decap_8
XFILLER_1_842 VPWR VGND sg13g2_decap_8
XFILLER_49_857 VPWR VGND sg13g2_decap_8
XFILLER_48_367 VPWR VGND sg13g2_decap_8
XFILLER_36_507 VPWR VGND sg13g2_decap_8
XFILLER_1_1024 VPWR VGND sg13g2_decap_4
XFILLER_17_710 VPWR VGND sg13g2_decap_8
XFILLER_44_584 VPWR VGND sg13g2_decap_8
XFILLER_17_787 VPWR VGND sg13g2_decap_8
XFILLER_32_735 VPWR VGND sg13g2_decap_8
XFILLER_13_971 VPWR VGND sg13g2_decap_8
XFILLER_20_919 VPWR VGND sg13g2_decap_8
XFILLER_31_256 VPWR VGND sg13g2_fill_2
X_2750_ _0319_ _0317_ _0318_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_441 VPWR VGND sg13g2_fill_1
X_2681_ VGND VPWR _1606_ _0273_ _1622_ net700 sg13g2_a21oi_2
XFILLER_9_964 VPWR VGND sg13g2_decap_8
XFILLER_4_691 VPWR VGND sg13g2_decap_8
X_3302_ net571 _0838_ VPWR VGND sg13g2_inv_4
X_3233_ _0769_ net649 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\] net651
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3164_ net684 _1782_ _1553_ _0700_ VPWR VGND sg13g2_nand3_1
XFILLER_39_367 VPWR VGND sg13g2_fill_2
X_3095_ _0617_ _0629_ _0630_ _0631_ VPWR VGND sg13g2_nor3_1
X_2115_ sap_3_inst.controller.stage\[1\] net719 _1536_ VPWR VGND sg13g2_xor2_1
XFILLER_27_529 VPWR VGND sg13g2_decap_8
X_2046_ VPWR _1469_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] VGND
+ sg13g2_inv_1
XFILLER_23_724 VPWR VGND sg13g2_decap_8
XFILLER_35_562 VPWR VGND sg13g2_decap_8
X_3997_ _1413_ VPWR _0187_ VGND _1432_ u_ser.state\[1\] sg13g2_o21ai_1
X_2948_ _0511_ _0482_ _0510_ VPWR VGND sg13g2_nand2_1
X_2879_ _0442_ _0443_ _0444_ VPWR VGND sg13g2_nor2_1
XFILLER_8_8 VPWR VGND sg13g2_fill_2
XFILLER_45_315 VPWR VGND sg13g2_decap_8
XFILLER_26_562 VPWR VGND sg13g2_decap_8
XFILLER_41_521 VPWR VGND sg13g2_decap_8
XFILLER_9_205 VPWR VGND sg13g2_fill_1
XFILLER_14_768 VPWR VGND sg13g2_decap_8
XFILLER_41_598 VPWR VGND sg13g2_decap_8
XFILLER_10_930 VPWR VGND sg13g2_decap_8
Xclkload19 VPWR clkload19/Y clknet_5_25__leaf_sap_3_inst.alu.clk_regs VGND sg13g2_inv_1
XFILLER_6_967 VPWR VGND sg13g2_decap_8
XFILLER_5_488 VPWR VGND sg13g2_decap_8
XFILLER_49_654 VPWR VGND sg13g2_decap_8
XFILLER_23_1025 VPWR VGND sg13g2_decap_4
XFILLER_37_849 VPWR VGND sg13g2_decap_8
X_3920_ _1354_ _1355_ _1352_ _1357_ VPWR VGND _1356_ sg13g2_nand4_1
XFILLER_17_584 VPWR VGND sg13g2_decap_8
XFILLER_32_532 VPWR VGND sg13g2_decap_8
X_3851_ _1293_ net769 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[6\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_20_716 VPWR VGND sg13g2_decap_8
X_3782_ VGND VPWR _1247_ _1246_ net579 sg13g2_or2_1
X_2802_ _1455_ _1550_ _1747_ _0370_ VPWR VGND sg13g2_nor3_1
X_2733_ _1612_ VPWR _0302_ VGND net723 _1576_ sg13g2_o21ai_1
XFILLER_9_761 VPWR VGND sg13g2_decap_8
XFILLER_30_1018 VPWR VGND sg13g2_decap_8
X_2664_ VGND VPWR _1604_ _1698_ _0257_ _1768_ sg13g2_a21oi_1
X_2595_ _2005_ _2001_ _2004_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_93 VPWR VGND sg13g2_fill_2
X_4196_ net781 VGND VPWR _0174_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\]
+ clknet_5_15__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3216_ _0752_ net644 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\] net653
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] VPWR VGND sg13g2_a22oi_1
X_3147_ _0681_ _0682_ _0679_ _0683_ VPWR VGND sg13g2_nand3_1
XFILLER_28_827 VPWR VGND sg13g2_decap_8
X_3078_ net673 _0613_ _0614_ VPWR VGND sg13g2_and2_1
XFILLER_36_871 VPWR VGND sg13g2_decap_8
X_2029_ _1452_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] VPWR VGND
+ sg13g2_inv_2
XFILLER_23_521 VPWR VGND sg13g2_decap_8
Xclkbuf_5_9__f_sap_3_inst.alu.clk_regs clknet_4_4_0_sap_3_inst.alu.clk_regs clknet_5_9__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_23_598 VPWR VGND sg13g2_decap_8
XFILLER_40_35 VPWR VGND sg13g2_fill_2
XFILLER_3_948 VPWR VGND sg13g2_decap_8
XFILLER_46_1025 VPWR VGND sg13g2_decap_4
XFILLER_2_469 VPWR VGND sg13g2_decap_8
Xfanout740 sap_3_inst.controller.opcode\[1\] net740 VPWR VGND sg13g2_buf_8
Xfanout751 net752 net751 VPWR VGND sg13g2_buf_8
Xfanout784 net785 net784 VPWR VGND sg13g2_buf_8
Xfanout773 net801 net773 VPWR VGND sg13g2_buf_8
Xfanout762 net763 net762 VPWR VGND sg13g2_buf_8
XFILLER_19_838 VPWR VGND sg13g2_decap_8
Xfanout795 net798 net795 VPWR VGND sg13g2_buf_8
XFILLER_46_668 VPWR VGND sg13g2_decap_8
XFILLER_27_893 VPWR VGND sg13g2_decap_8
XFILLER_42_874 VPWR VGND sg13g2_decap_8
XFILLER_14_565 VPWR VGND sg13g2_decap_8
XFILLER_6_764 VPWR VGND sg13g2_decap_8
X_2380_ net662 _1762_ _1791_ _1801_ VPWR VGND sg13g2_nor3_2
XFILLER_49_451 VPWR VGND sg13g2_decap_8
X_4050_ net772 VGND VPWR _0004_ sap_3_inst.controller.stage\[2\] net42 sg13g2_dfrbpq_2
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
X_3001_ _0561_ sap_3_inst.out\[1\] net673 VPWR VGND sg13g2_nand2_1
XFILLER_37_646 VPWR VGND sg13g2_decap_8
XFILLER_33_830 VPWR VGND sg13g2_decap_8
Xclkbuf_5_16__f_sap_3_inst.alu.clk_regs clknet_4_8_0_sap_3_inst.alu.clk_regs clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3903_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] _1341_
+ _1312_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] _1342_ _1306_ sg13g2_a221oi_1
XFILLER_20_513 VPWR VGND sg13g2_decap_8
X_3834_ _1281_ sap_3_inst.reg_file.array_serializer_inst.state\[0\] VPWR VGND sap_3_inst.reg_file.array_serializer_inst.state\[1\]
+ sg13g2_nand2b_2
X_3765_ net12 net599 _1231_ _1233_ _1234_ VPWR VGND sg13g2_nor4_1
X_2716_ _1538_ VPWR _0295_ VGND _1548_ _0294_ sg13g2_o21ai_1
X_3696_ _0958_ net579 _1059_ _1188_ VPWR VGND sg13g2_a21o_2
X_2647_ _0242_ net628 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] net678
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_0_918 VPWR VGND sg13g2_decap_8
X_2578_ _1989_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] net637
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_28_624 VPWR VGND sg13g2_decap_8
X_4029__7 VPWR net41 clknet_leaf_0_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_27_123 VPWR VGND sg13g2_fill_1
X_4179_ net799 VGND VPWR net81 sap_3_inst.reg_file.array_serializer_inst.bit_pos\[0\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_43_649 VPWR VGND sg13g2_decap_8
XFILLER_24_841 VPWR VGND sg13g2_decap_8
XFILLER_35_68 VPWR VGND sg13g2_fill_1
XFILLER_11_557 VPWR VGND sg13g2_decap_8
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_7_517 VPWR VGND sg13g2_decap_8
XFILLER_13_1013 VPWR VGND sg13g2_decap_8
XFILLER_3_745 VPWR VGND sg13g2_decap_8
Xfanout592 _0738_ net592 VPWR VGND sg13g2_buf_8
Xfanout570 _1077_ net570 VPWR VGND sg13g2_buf_8
Xfanout581 net582 net581 VPWR VGND sg13g2_buf_1
XFILLER_47_955 VPWR VGND sg13g2_decap_8
XFILLER_19_635 VPWR VGND sg13g2_decap_8
XFILLER_20_1017 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_465 VPWR VGND sg13g2_decap_8
XFILLER_27_690 VPWR VGND sg13g2_decap_8
XFILLER_34_627 VPWR VGND sg13g2_decap_8
XFILLER_42_671 VPWR VGND sg13g2_decap_8
XFILLER_15_885 VPWR VGND sg13g2_decap_8
XFILLER_30_822 VPWR VGND sg13g2_decap_8
XFILLER_30_899 VPWR VGND sg13g2_decap_8
X_3550_ _1002_ net557 _1068_ _1072_ VPWR VGND sg13g2_nor3_1
X_2501_ _1916_ net629 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] net631
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_561 VPWR VGND sg13g2_decap_8
X_3481_ _1011_ net547 net571 VPWR VGND sg13g2_nand2_1
X_2432_ _1853_ net633 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] net677
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2363_ _1783_ VPWR _1784_ VGND _1546_ _1549_ sg13g2_o21ai_1
X_4102_ net776 VGND VPWR _0080_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2294_ VGND VPWR _1715_ _1713_ _1540_ sg13g2_or2_1
XFILLER_38_900 VPWR VGND sg13g2_decap_8
XFILLER_49_270 VPWR VGND sg13g2_decap_4
XFILLER_38_977 VPWR VGND sg13g2_decap_8
XFILLER_21_800 VPWR VGND sg13g2_decap_8
X_3817_ net13 net603 _1269_ VPWR VGND sg13g2_nor2_1
XFILLER_21_877 VPWR VGND sg13g2_decap_8
X_3748_ _0856_ _0744_ _1219_ _1220_ VPWR VGND sg13g2_a21o_1
XFILLER_4_509 VPWR VGND sg13g2_decap_8
X_3679_ VGND VPWR _1176_ _1175_ net661 sg13g2_or2_1
XFILLER_43_1006 VPWR VGND sg13g2_decap_8
XFILLER_0_715 VPWR VGND sg13g2_decap_8
XFILLER_29_944 VPWR VGND sg13g2_decap_8
XFILLER_15_115 VPWR VGND sg13g2_fill_2
XFILLER_16_627 VPWR VGND sg13g2_decap_8
XFILLER_28_498 VPWR VGND sg13g2_decap_8
XFILLER_44_969 VPWR VGND sg13g2_decap_8
XFILLER_43_446 VPWR VGND sg13g2_decap_8
XFILLER_8_804 VPWR VGND sg13g2_decap_8
XFILLER_12_833 VPWR VGND sg13g2_decap_8
XFILLER_7_39 VPWR VGND sg13g2_fill_2
XFILLER_3_542 VPWR VGND sg13g2_decap_8
XFILLER_39_719 VPWR VGND sg13g2_decap_8
XFILLER_47_752 VPWR VGND sg13g2_decap_8
XFILLER_46_240 VPWR VGND sg13g2_fill_2
XFILLER_35_947 VPWR VGND sg13g2_decap_8
X_2981_ _0543_ _0542_ _0511_ VPWR VGND sg13g2_nand2b_1
XFILLER_15_682 VPWR VGND sg13g2_decap_8
XFILLER_30_696 VPWR VGND sg13g2_decap_8
X_3602_ _1116_ net591 _1007_ VPWR VGND sg13g2_nand2b_1
XFILLER_7_881 VPWR VGND sg13g2_decap_8
X_3533_ VPWR _0078_ _1057_ VGND sg13g2_inv_1
X_3464_ _0994_ _0989_ _0993_ net615 _1479_ VPWR VGND sg13g2_a22oi_1
X_2415_ net685 _1568_ net689 _1836_ VPWR VGND sg13g2_a21o_1
X_3395_ VGND VPWR _0787_ _0850_ _0928_ net574 sg13g2_a21oi_1
X_2346_ _1767_ _1533_ _1633_ VPWR VGND sg13g2_nand2_1
X_2277_ VGND VPWR _1584_ _1698_ _1647_ _1559_ sg13g2_a21oi_2
X_4016_ VPWR _0192_ _1427_ VGND sg13g2_inv_1
XFILLER_38_774 VPWR VGND sg13g2_decap_8
XFILLER_26_947 VPWR VGND sg13g2_decap_8
XFILLER_41_906 VPWR VGND sg13g2_decap_8
XFILLER_25_457 VPWR VGND sg13g2_decap_8
XFILLER_12_107 VPWR VGND sg13g2_fill_2
XFILLER_34_991 VPWR VGND sg13g2_decap_8
XFILLER_21_674 VPWR VGND sg13g2_decap_8
XFILLER_0_512 VPWR VGND sg13g2_decap_8
XFILLER_0_589 VPWR VGND sg13g2_decap_8
XFILLER_48_549 VPWR VGND sg13g2_decap_8
XFILLER_29_741 VPWR VGND sg13g2_decap_8
XFILLER_44_766 VPWR VGND sg13g2_decap_8
XFILLER_17_969 VPWR VGND sg13g2_decap_8
XFILLER_32_917 VPWR VGND sg13g2_decap_8
XFILLER_43_298 VPWR VGND sg13g2_fill_1
XFILLER_12_630 VPWR VGND sg13g2_decap_8
XFILLER_8_601 VPWR VGND sg13g2_decap_8
XFILLER_8_678 VPWR VGND sg13g2_decap_8
XFILLER_4_873 VPWR VGND sg13g2_decap_8
X_2200_ net732 sap_3_inst.alu.flags\[0\] net720 sap_3_inst.alu.flags\[2\] sap_3_inst.alu.flags\[3\]
+ net730 _1621_ VPWR VGND sg13g2_mux4_1
X_3180_ _0716_ net614 VPWR VGND _0635_ sg13g2_nand2b_2
XFILLER_39_516 VPWR VGND sg13g2_decap_8
X_2131_ _1552_ _1550_ _1546_ VPWR VGND sg13g2_nand2b_1
X_2062_ VPWR _1485_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_23_906 VPWR VGND sg13g2_decap_8
XFILLER_35_744 VPWR VGND sg13g2_decap_8
X_2964_ net544 _0526_ _0527_ VPWR VGND sg13g2_nor2b_1
XFILLER_16_991 VPWR VGND sg13g2_decap_8
XFILLER_33_1005 VPWR VGND sg13g2_decap_8
X_2895_ _0460_ _0458_ _0322_ net572 net749 VPWR VGND sg13g2_a22oi_1
XFILLER_30_493 VPWR VGND sg13g2_decap_8
X_3516_ net583 _0876_ _1043_ VPWR VGND sg13g2_nor2_1
X_3447_ VGND VPWR net14 _0838_ _0978_ _0632_ sg13g2_a21oi_1
X_3378_ _0911_ net656 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] net608
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2329_ _1750_ _1615_ _1641_ VPWR VGND sg13g2_nand2_1
XFILLER_38_571 VPWR VGND sg13g2_decap_8
XFILLER_26_744 VPWR VGND sg13g2_decap_8
XFILLER_41_703 VPWR VGND sg13g2_decap_8
XFILLER_40_202 VPWR VGND sg13g2_fill_2
XFILLER_4_147 VPWR VGND sg13g2_fill_2
XFILLER_1_821 VPWR VGND sg13g2_decap_8
XFILLER_49_836 VPWR VGND sg13g2_decap_8
XFILLER_1_898 VPWR VGND sg13g2_decap_8
XFILLER_48_346 VPWR VGND sg13g2_decap_8
XFILLER_1_1003 VPWR VGND sg13g2_decap_8
XFILLER_44_563 VPWR VGND sg13g2_decap_8
XFILLER_17_91 VPWR VGND sg13g2_fill_1
XFILLER_17_766 VPWR VGND sg13g2_decap_8
XFILLER_32_714 VPWR VGND sg13g2_decap_8
XFILLER_13_950 VPWR VGND sg13g2_decap_8
XFILLER_9_943 VPWR VGND sg13g2_decap_8
X_2680_ VGND VPWR _1623_ _0271_ _0272_ _0267_ sg13g2_a21oi_1
XFILLER_4_670 VPWR VGND sg13g2_decap_8
X_3301_ _0837_ net614 _0836_ VPWR VGND sg13g2_nand2b_1
X_3232_ _0768_ net643 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] net646
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3163_ _1581_ _1614_ _1575_ _0699_ VPWR VGND sg13g2_nand3_1
X_2114_ _1535_ net719 net718 VPWR VGND sg13g2_xnor2_1
XFILLER_27_508 VPWR VGND sg13g2_decap_8
X_3094_ net695 _1606_ _1622_ _0630_ VPWR VGND sg13g2_nor3_1
X_2045_ _1468_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[4\] VPWR VGND
+ sg13g2_inv_2
XFILLER_35_541 VPWR VGND sg13g2_decap_8
XFILLER_23_703 VPWR VGND sg13g2_decap_8
XFILLER_22_224 VPWR VGND sg13g2_fill_2
X_3996_ _1410_ VPWR _1413_ VGND _1434_ _1411_ sg13g2_o21ai_1
X_2947_ _0510_ _0507_ _0508_ VPWR VGND sg13g2_xnor2_1
X_2878_ VGND VPWR net754 net671 _0443_ _0413_ sg13g2_a21oi_1
XFILLER_39_880 VPWR VGND sg13g2_decap_8
XFILLER_45_349 VPWR VGND sg13g2_fill_1
XFILLER_26_541 VPWR VGND sg13g2_decap_8
XFILLER_41_500 VPWR VGND sg13g2_decap_8
XFILLER_14_747 VPWR VGND sg13g2_decap_8
XFILLER_41_577 VPWR VGND sg13g2_decap_8
XFILLER_6_946 VPWR VGND sg13g2_decap_8
XFILLER_10_986 VPWR VGND sg13g2_decap_8
XFILLER_5_467 VPWR VGND sg13g2_decap_8
XFILLER_49_633 VPWR VGND sg13g2_decap_8
XFILLER_1_695 VPWR VGND sg13g2_decap_8
XFILLER_23_1004 VPWR VGND sg13g2_decap_8
XFILLER_37_828 VPWR VGND sg13g2_decap_8
XFILLER_17_563 VPWR VGND sg13g2_decap_8
XFILLER_32_511 VPWR VGND sg13g2_decap_8
X_3850_ net769 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[1\] sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[2\]
+ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[3\] sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[4\]
+ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\] _1292_ VPWR VGND sg13g2_mux4_1
X_3781_ VPWR VGND _0633_ _1074_ _1245_ net661 _1246_ _1244_ sg13g2_a221oi_1
X_2801_ VGND VPWR _0345_ _0368_ _0369_ _0325_ sg13g2_a21oi_1
Xclkbuf_0_sap_3_inst.alu.clk sap_3_inst.alu.clk clknet_0_sap_3_inst.alu.clk VPWR VGND
+ sg13g2_buf_8
XFILLER_32_588 VPWR VGND sg13g2_decap_8
X_2732_ _0301_ _1551_ _1757_ VPWR VGND sg13g2_nand2_1
XFILLER_9_740 VPWR VGND sg13g2_decap_8
X_2663_ sap_3_inst.alu.flags\[0\] _0256_ _0248_ _0026_ VPWR VGND sg13g2_mux2_1
X_2594_ _2004_ _2002_ _2003_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_83 VPWR VGND sg13g2_decap_4
X_3215_ _0751_ _0748_ _0749_ _0750_ VPWR VGND sg13g2_and3_2
X_4195_ net793 VGND VPWR _0173_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\]
+ clknet_5_28__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_806 VPWR VGND sg13g2_decap_8
X_3146_ _0676_ VPWR _0682_ VGND _1601_ net708 sg13g2_o21ai_1
X_3077_ _0613_ _1575_ _1703_ VPWR VGND sg13g2_nand2b_1
X_2028_ VPWR _1451_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_36_850 VPWR VGND sg13g2_decap_8
XFILLER_23_500 VPWR VGND sg13g2_decap_8
XFILLER_11_739 VPWR VGND sg13g2_decap_8
XFILLER_23_577 VPWR VGND sg13g2_decap_8
X_3979_ _1401_ sap_3_inst.alu.act\[3\] net548 VPWR VGND sg13g2_nand2_1
XFILLER_40_47 VPWR VGND sg13g2_fill_2
XFILLER_3_927 VPWR VGND sg13g2_decap_8
XFILLER_46_1004 VPWR VGND sg13g2_decap_8
XFILLER_2_448 VPWR VGND sg13g2_decap_8
XFILLER_49_23 VPWR VGND sg13g2_fill_1
Xfanout741 net742 net741 VPWR VGND sg13g2_buf_8
Xfanout730 sap_3_inst.controller.opcode\[5\] net730 VPWR VGND sg13g2_buf_8
Xfanout763 _1310_ net763 VPWR VGND sg13g2_buf_8
Xfanout785 net792 net785 VPWR VGND sg13g2_buf_8
Xfanout752 sap_3_inst.alu.acc\[4\] net752 VPWR VGND sg13g2_buf_8
Xfanout774 net778 net774 VPWR VGND sg13g2_buf_8
Xfanout796 net797 net796 VPWR VGND sg13g2_buf_8
XFILLER_19_817 VPWR VGND sg13g2_decap_8
XFILLER_46_647 VPWR VGND sg13g2_decap_8
XFILLER_34_809 VPWR VGND sg13g2_decap_8
XFILLER_45_157 VPWR VGND sg13g2_fill_2
XFILLER_27_872 VPWR VGND sg13g2_decap_8
XFILLER_42_853 VPWR VGND sg13g2_decap_8
XFILLER_14_544 VPWR VGND sg13g2_decap_8
XFILLER_6_743 VPWR VGND sg13g2_decap_8
XFILLER_10_783 VPWR VGND sg13g2_decap_8
XFILLER_49_430 VPWR VGND sg13g2_decap_8
XFILLER_1_492 VPWR VGND sg13g2_decap_8
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
X_3000_ _0560_ VPWR _0042_ VGND _1456_ net673 sg13g2_o21ai_1
XFILLER_37_625 VPWR VGND sg13g2_decap_8
XFILLER_18_894 VPWR VGND sg13g2_decap_8
X_3902_ _1338_ _1339_ _1337_ _1341_ VPWR VGND _1340_ sg13g2_nand4_1
XFILLER_33_886 VPWR VGND sg13g2_decap_8
X_3833_ VPWR _0155_ net764 VGND sg13g2_inv_1
XFILLER_20_569 VPWR VGND sg13g2_decap_8
X_3764_ _0920_ _1232_ _1233_ VPWR VGND sg13g2_nor2_1
X_2715_ VGND VPWR _1569_ _0293_ _0294_ _1572_ sg13g2_a21oi_1
X_3695_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] _1130_ _1182_ _0110_
+ VPWR VGND sg13g2_mux2_1
X_2646_ _0241_ _1800_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] _1798_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2577_ VPWR VGND net3 _1987_ _1847_ net756 _1988_ _1827_ sg13g2_a221oi_1
XFILLER_28_603 VPWR VGND sg13g2_decap_8
X_4178_ net799 VGND VPWR _0156_ sap_3_inst.reg_file.array_serializer_inst.state\[1\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
X_3129_ _0663_ _0664_ _0662_ _0665_ VPWR VGND sg13g2_nand3_1
XFILLER_16_809 VPWR VGND sg13g2_decap_8
XFILLER_43_628 VPWR VGND sg13g2_decap_8
XFILLER_24_820 VPWR VGND sg13g2_decap_8
XFILLER_23_374 VPWR VGND sg13g2_decap_4
XFILLER_24_897 VPWR VGND sg13g2_decap_8
XFILLER_11_536 VPWR VGND sg13g2_decap_8
XFILLER_3_724 VPWR VGND sg13g2_decap_8
XFILLER_2_256 VPWR VGND sg13g2_fill_1
Xfanout560 net561 net560 VPWR VGND sg13g2_buf_8
XFILLER_19_614 VPWR VGND sg13g2_decap_8
Xfanout571 _0837_ net571 VPWR VGND sg13g2_buf_8
Xfanout593 _0738_ net593 VPWR VGND sg13g2_buf_1
Xfanout582 _0842_ net582 VPWR VGND sg13g2_buf_8
XFILLER_47_934 VPWR VGND sg13g2_decap_8
XFILLER_46_444 VPWR VGND sg13g2_decap_8
XFILLER_34_606 VPWR VGND sg13g2_decap_8
XFILLER_15_864 VPWR VGND sg13g2_decap_8
XFILLER_42_650 VPWR VGND sg13g2_decap_8
XFILLER_30_801 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_2_sap_3_inst.alu.clk clknet_1_1__leaf_sap_3_inst.alu.clk clknet_leaf_2_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_30_878 VPWR VGND sg13g2_decap_8
XFILLER_10_580 VPWR VGND sg13g2_decap_8
X_2500_ _1915_ net619 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] net627
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_540 VPWR VGND sg13g2_decap_8
X_3480_ _1009_ VPWR _1010_ VGND net611 _1006_ sg13g2_o21ai_1
X_2431_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] net621
+ net635 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] _1852_ net638 sg13g2_a221oi_1
XFILLER_29_1021 VPWR VGND sg13g2_decap_8
X_2362_ _1438_ _1500_ _1528_ _1781_ _1783_ VPWR VGND sg13g2_nor4_1
X_4101_ net776 VGND VPWR _0079_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\]
+ clknet_5_9__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2293_ _1540_ _1713_ _1714_ VPWR VGND sg13g2_nor2_1
XFILLER_38_956 VPWR VGND sg13g2_decap_8
XFILLER_25_639 VPWR VGND sg13g2_decap_8
XFILLER_37_499 VPWR VGND sg13g2_decap_8
XFILLER_18_691 VPWR VGND sg13g2_decap_8
XFILLER_33_683 VPWR VGND sg13g2_decap_8
XFILLER_36_1025 VPWR VGND sg13g2_decap_4
XFILLER_21_856 VPWR VGND sg13g2_decap_8
X_3816_ _1264_ VPWR _0150_ VGND _1265_ _1268_ sg13g2_o21ai_1
X_3747_ _1219_ _0844_ _0857_ VPWR VGND sg13g2_nand2b_1
X_3678_ net16 net24 net568 _1175_ VPWR VGND sg13g2_mux2_1
X_4031__9 VPWR net43 clknet_leaf_3_sap_3_inst.alu.clk VGND sg13g2_inv_1
X_2629_ VPWR _0225_ net32 VGND sg13g2_inv_1
XFILLER_29_923 VPWR VGND sg13g2_decap_8
XFILLER_16_606 VPWR VGND sg13g2_decap_8
XFILLER_44_948 VPWR VGND sg13g2_decap_8
XFILLER_43_425 VPWR VGND sg13g2_decap_8
XFILLER_28_477 VPWR VGND sg13g2_decap_8
XFILLER_12_812 VPWR VGND sg13g2_decap_8
XFILLER_23_182 VPWR VGND sg13g2_decap_4
XFILLER_24_694 VPWR VGND sg13g2_decap_8
XFILLER_7_18 VPWR VGND sg13g2_fill_1
XFILLER_12_889 VPWR VGND sg13g2_decap_8
XFILLER_3_521 VPWR VGND sg13g2_decap_8
XFILLER_11_82 VPWR VGND sg13g2_fill_1
XFILLER_3_598 VPWR VGND sg13g2_decap_8
XFILLER_47_731 VPWR VGND sg13g2_decap_8
XFILLER_19_488 VPWR VGND sg13g2_decap_8
XFILLER_35_926 VPWR VGND sg13g2_decap_8
XFILLER_15_661 VPWR VGND sg13g2_decap_8
X_2980_ _0542_ _0540_ _0541_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_992 VPWR VGND sg13g2_decap_8
X_3601_ VGND VPWR net581 _0999_ _1115_ net590 sg13g2_a21oi_1
XFILLER_30_675 VPWR VGND sg13g2_decap_8
XFILLER_7_860 VPWR VGND sg13g2_decap_8
X_3532_ _1057_ _1054_ _1056_ net557 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_6_381 VPWR VGND sg13g2_fill_2
X_3463_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] _0992_
+ net657 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] _0993_ net609 sg13g2_a221oi_1
X_2414_ VGND VPWR _1582_ _1834_ _1835_ _1616_ sg13g2_a21oi_1
X_3394_ VGND VPWR net546 _0837_ _0927_ _0926_ sg13g2_a21oi_1
XFILLER_35_0 VPWR VGND sg13g2_fill_1
X_2345_ net723 _1612_ _1727_ _1766_ VPWR VGND sg13g2_nor3_1
X_2276_ VPWR _1697_ _1696_ VGND sg13g2_inv_1
X_4015_ _1427_ _1425_ net79 _1424_ net761 VPWR VGND sg13g2_a22oi_1
XFILLER_38_753 VPWR VGND sg13g2_decap_8
XFILLER_26_926 VPWR VGND sg13g2_decap_8
XFILLER_25_436 VPWR VGND sg13g2_decap_8
XFILLER_34_970 VPWR VGND sg13g2_decap_8
XFILLER_21_653 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_568 VPWR VGND sg13g2_decap_8
XFILLER_48_528 VPWR VGND sg13g2_decap_8
XFILLER_29_720 VPWR VGND sg13g2_decap_8
XFILLER_17_948 VPWR VGND sg13g2_decap_8
XFILLER_29_797 VPWR VGND sg13g2_decap_8
XFILLER_44_745 VPWR VGND sg13g2_decap_8
XFILLER_19_1020 VPWR VGND sg13g2_decap_8
XFILLER_24_491 VPWR VGND sg13g2_decap_8
XFILLER_40_984 VPWR VGND sg13g2_decap_8
XFILLER_12_686 VPWR VGND sg13g2_decap_8
XFILLER_8_657 VPWR VGND sg13g2_decap_8
XFILLER_4_852 VPWR VGND sg13g2_decap_8
XFILLER_3_362 VPWR VGND sg13g2_fill_2
XFILLER_26_1024 VPWR VGND sg13g2_decap_4
X_2130_ _1546_ _1549_ _1551_ VPWR VGND sg13g2_nor2_2
X_2061_ VPWR _1484_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_35_723 VPWR VGND sg13g2_decap_8
XFILLER_16_970 VPWR VGND sg13g2_decap_8
XFILLER_34_244 VPWR VGND sg13g2_fill_1
X_2963_ _0513_ _0519_ _0524_ _0525_ _0526_ VPWR VGND sg13g2_nor4_1
X_2894_ _0432_ _0458_ _0459_ VPWR VGND sg13g2_nor2_1
XFILLER_30_472 VPWR VGND sg13g2_decap_8
XFILLER_31_995 VPWR VGND sg13g2_decap_8
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_94 VPWR VGND sg13g2_decap_8
X_3515_ net557 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[0\] _1042_ _0075_
+ VPWR VGND sg13g2_a21o_1
X_3446_ VGND VPWR net612 _0973_ _0977_ _0976_ sg13g2_a21oi_1
X_3377_ _0909_ VPWR _0910_ VGND _1443_ net590 sg13g2_o21ai_1
X_2328_ _1616_ _1641_ _1749_ VPWR VGND sg13g2_nor2b_1
X_2259_ _1589_ VPWR _1680_ VGND _1580_ _1646_ sg13g2_o21ai_1
XFILLER_26_723 VPWR VGND sg13g2_decap_8
XFILLER_27_48 VPWR VGND sg13g2_fill_1
XFILLER_27_59 VPWR VGND sg13g2_fill_2
XFILLER_38_550 VPWR VGND sg13g2_decap_8
XFILLER_14_929 VPWR VGND sg13g2_decap_8
XFILLER_41_759 VPWR VGND sg13g2_decap_8
XFILLER_22_995 VPWR VGND sg13g2_decap_8
XFILLER_5_649 VPWR VGND sg13g2_decap_8
XFILLER_1_800 VPWR VGND sg13g2_decap_8
XFILLER_49_815 VPWR VGND sg13g2_decap_8
XFILLER_1_877 VPWR VGND sg13g2_decap_8
XFILLER_48_325 VPWR VGND sg13g2_decap_8
XFILLER_44_542 VPWR VGND sg13g2_decap_8
XFILLER_17_745 VPWR VGND sg13g2_decap_8
XFILLER_29_594 VPWR VGND sg13g2_decap_8
XFILLER_31_258 VPWR VGND sg13g2_fill_1
XFILLER_40_781 VPWR VGND sg13g2_decap_8
XFILLER_9_922 VPWR VGND sg13g2_decap_8
XFILLER_9_999 VPWR VGND sg13g2_decap_8
X_3300_ _0692_ _0835_ _0836_ VPWR VGND sg13g2_nor2_2
X_3231_ _0759_ _0764_ _0758_ _0767_ VPWR VGND _0765_ sg13g2_nand4_1
X_3162_ _0697_ net686 _1590_ _0698_ VPWR VGND sg13g2_a21o_1
X_2113_ _1534_ _1499_ _1533_ VPWR VGND sg13g2_nand2_1
X_3093_ _0627_ VPWR _0629_ VGND net708 _0628_ sg13g2_o21ai_1
XFILLER_48_892 VPWR VGND sg13g2_decap_8
X_2044_ VPWR _1467_ sap_3_inst.alu.tmp\[6\] VGND sg13g2_inv_1
XFILLER_35_520 VPWR VGND sg13g2_decap_8
XFILLER_35_597 VPWR VGND sg13g2_decap_8
X_3995_ _1412_ _1410_ _1411_ VPWR VGND sg13g2_nand2_1
XFILLER_23_759 VPWR VGND sg13g2_decap_8
X_2946_ _0507_ _0508_ _0509_ VPWR VGND sg13g2_nor2_1
X_2877_ _0442_ net751 net671 VPWR VGND sg13g2_xnor2_1
XFILLER_30_291 VPWR VGND sg13g2_fill_1
XFILLER_31_792 VPWR VGND sg13g2_decap_8
XFILLER_1_107 VPWR VGND sg13g2_fill_2
X_3429_ _0936_ VPWR _0071_ VGND _0954_ _0960_ sg13g2_o21ai_1
XFILLER_46_829 VPWR VGND sg13g2_decap_8
XFILLER_18_509 VPWR VGND sg13g2_decap_8
XFILLER_26_520 VPWR VGND sg13g2_decap_8
XFILLER_14_726 VPWR VGND sg13g2_decap_8
XFILLER_26_597 VPWR VGND sg13g2_decap_8
XFILLER_41_556 VPWR VGND sg13g2_decap_8
XFILLER_16_1012 VPWR VGND sg13g2_decap_8
XFILLER_22_792 VPWR VGND sg13g2_decap_8
XFILLER_6_925 VPWR VGND sg13g2_decap_8
XFILLER_10_965 VPWR VGND sg13g2_decap_8
Xclkbuf_5_24__f_sap_3_inst.alu.clk_regs clknet_4_12_0_sap_3_inst.alu.clk_regs clknet_5_24__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_49_612 VPWR VGND sg13g2_decap_8
XFILLER_1_674 VPWR VGND sg13g2_decap_8
XFILLER_37_807 VPWR VGND sg13g2_decap_8
XFILLER_49_689 VPWR VGND sg13g2_decap_8
XFILLER_44_350 VPWR VGND sg13g2_fill_1
XFILLER_17_542 VPWR VGND sg13g2_decap_8
XFILLER_45_884 VPWR VGND sg13g2_decap_8
XFILLER_32_567 VPWR VGND sg13g2_decap_8
X_3780_ _1245_ net655 net16 VPWR VGND sg13g2_nand2b_1
X_2800_ _0355_ _0320_ _0368_ VPWR VGND sg13g2_xor2_1
X_2731_ _0300_ _1839_ _1716_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_262 VPWR VGND sg13g2_fill_2
XFILLER_9_796 VPWR VGND sg13g2_decap_8
X_2662_ net31 _0255_ _1858_ _0256_ VPWR VGND sg13g2_mux2_1
X_2593_ net751 net747 _2003_ VPWR VGND sg13g2_xor2_1
XFILLER_5_62 VPWR VGND sg13g2_fill_2
X_3214_ _0750_ net640 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] net612
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4194_ net773 VGND VPWR _0172_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\]
+ clknet_5_7__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3145_ _0681_ _1623_ _0680_ VPWR VGND sg13g2_nand2_1
X_3076_ _1615_ VPWR _0612_ VGND net687 _1691_ sg13g2_o21ai_1
X_2027_ VPWR _1450_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_23_556 VPWR VGND sg13g2_decap_8
X_3978_ VGND VPWR net753 net663 _1400_ _1399_ sg13g2_a21oi_1
XFILLER_11_718 VPWR VGND sg13g2_decap_8
X_2929_ _0493_ _0452_ _0491_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_906 VPWR VGND sg13g2_decap_8
Xfanout720 sap_3_inst.alu.flags\[1\] net720 VPWR VGND sg13g2_buf_8
Xfanout731 net732 net731 VPWR VGND sg13g2_buf_8
Xfanout742 sap_3_inst.controller.opcode\[0\] net742 VPWR VGND sg13g2_buf_2
Xfanout775 net777 net775 VPWR VGND sg13g2_buf_8
Xfanout753 net754 net753 VPWR VGND sg13g2_buf_8
Xfanout764 net765 net764 VPWR VGND sg13g2_buf_8
XFILLER_46_626 VPWR VGND sg13g2_decap_8
Xfanout786 net792 net786 VPWR VGND sg13g2_buf_8
Xfanout797 net798 net797 VPWR VGND sg13g2_buf_8
XFILLER_27_851 VPWR VGND sg13g2_decap_8
XFILLER_42_832 VPWR VGND sg13g2_decap_8
XFILLER_14_523 VPWR VGND sg13g2_decap_8
XFILLER_26_394 VPWR VGND sg13g2_decap_8
XFILLER_10_762 VPWR VGND sg13g2_decap_8
XFILLER_6_722 VPWR VGND sg13g2_decap_8
XFILLER_6_799 VPWR VGND sg13g2_decap_8
XFILLER_2_994 VPWR VGND sg13g2_decap_8
XFILLER_1_471 VPWR VGND sg13g2_decap_8
XFILLER_7_1021 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
XFILLER_37_604 VPWR VGND sg13g2_decap_8
XFILLER_49_486 VPWR VGND sg13g2_decap_8
XFILLER_45_681 VPWR VGND sg13g2_decap_8
XFILLER_18_873 VPWR VGND sg13g2_decap_8
X_3901_ _1340_ _1313_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] _1305_
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_865 VPWR VGND sg13g2_decap_8
X_3832_ VGND VPWR _1280_ sap_3_inst.reg_file.array_serializer_inst.state\[1\] sap_3_inst.reg_file.array_serializer_inst.state\[0\]
+ sg13g2_or2_1
XFILLER_20_548 VPWR VGND sg13g2_decap_8
X_3763_ net580 VPWR _1232_ VGND net655 _0924_ sg13g2_o21ai_1
X_2714_ _0293_ _1619_ _0292_ VPWR VGND sg13g2_nand2_1
XFILLER_9_593 VPWR VGND sg13g2_decap_8
X_3694_ _0109_ _1187_ _1049_ _1181_ _1450_ VPWR VGND sg13g2_a22oi_1
X_2645_ _0240_ _0238_ _0239_ VPWR VGND sg13g2_nand2_1
X_2576_ sap_3_inst.alu.flags\[2\] _1828_ _1987_ VPWR VGND sg13g2_and2_1
X_4177_ net799 VGND VPWR _0155_ sap_3_inst.reg_file.array_serializer_inst.state\[0\]
+ clknet_3_6__leaf_clk sg13g2_dfrbpq_2
X_3128_ _0664_ _0659_ _1575_ net706 _1577_ VPWR VGND sg13g2_a22oi_1
XFILLER_43_607 VPWR VGND sg13g2_decap_8
XFILLER_28_659 VPWR VGND sg13g2_decap_8
X_3059_ _0596_ VPWR _0065_ VGND net691 net547 sg13g2_o21ai_1
XFILLER_11_515 VPWR VGND sg13g2_decap_8
XFILLER_24_876 VPWR VGND sg13g2_decap_8
XFILLER_3_703 VPWR VGND sg13g2_decap_8
Xfanout550 _1126_ net550 VPWR VGND sg13g2_buf_8
XFILLER_47_913 VPWR VGND sg13g2_decap_8
Xfanout572 _0339_ net572 VPWR VGND sg13g2_buf_8
Xfanout583 _0830_ net583 VPWR VGND sg13g2_buf_8
Xfanout561 _0796_ net561 VPWR VGND sg13g2_buf_8
XFILLER_46_423 VPWR VGND sg13g2_decap_8
Xfanout594 _0734_ net594 VPWR VGND sg13g2_buf_8
XFILLER_15_843 VPWR VGND sg13g2_decap_8
XFILLER_30_857 VPWR VGND sg13g2_decap_8
XFILLER_41_80 VPWR VGND sg13g2_fill_1
X_2430_ _1851_ net625 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] net627
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_596 VPWR VGND sg13g2_decap_8
XFILLER_29_1000 VPWR VGND sg13g2_decap_8
X_2361_ _1438_ _1781_ _1782_ VPWR VGND sg13g2_nor2_1
XFILLER_2_791 VPWR VGND sg13g2_decap_8
X_2292_ _1511_ VPWR _1713_ VGND net722 _1564_ sg13g2_o21ai_1
X_4100_ net793 VGND VPWR _0078_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\]
+ clknet_5_27__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_2_30 VPWR VGND sg13g2_decap_8
XFILLER_38_935 VPWR VGND sg13g2_decap_8
XFILLER_2_96 VPWR VGND sg13g2_fill_2
XFILLER_46_990 VPWR VGND sg13g2_decap_8
XFILLER_18_670 VPWR VGND sg13g2_decap_8
XFILLER_25_618 VPWR VGND sg13g2_decap_8
XFILLER_33_662 VPWR VGND sg13g2_decap_8
XFILLER_36_1004 VPWR VGND sg13g2_decap_8
XFILLER_21_835 VPWR VGND sg13g2_decap_8
X_3815_ VPWR VGND _0633_ _0929_ _1267_ _0933_ _1268_ _1266_ sg13g2_a221oi_1
X_3746_ net656 VPWR _1218_ VGND net575 _0860_ sg13g2_o21ai_1
X_3677_ net578 _1173_ _1174_ VPWR VGND sg13g2_nor2_1
X_2628_ _0215_ _0224_ _0214_ net18 VPWR VGND sg13g2_nand3_1
X_2559_ _1972_ _1969_ _1970_ _1971_ VPWR VGND sg13g2_and3_1
XFILLER_29_902 VPWR VGND sg13g2_decap_8
XFILLER_28_456 VPWR VGND sg13g2_decap_8
XFILLER_29_979 VPWR VGND sg13g2_decap_8
XFILLER_46_69 VPWR VGND sg13g2_fill_1
XFILLER_44_927 VPWR VGND sg13g2_decap_8
XFILLER_43_404 VPWR VGND sg13g2_decap_8
XFILLER_15_106 VPWR VGND sg13g2_fill_2
XFILLER_24_673 VPWR VGND sg13g2_decap_8
XFILLER_12_868 VPWR VGND sg13g2_decap_8
XFILLER_8_839 VPWR VGND sg13g2_decap_8
XFILLER_3_500 VPWR VGND sg13g2_decap_8
XFILLER_3_577 VPWR VGND sg13g2_decap_8
XFILLER_47_710 VPWR VGND sg13g2_decap_8
XFILLER_4_1013 VPWR VGND sg13g2_decap_8
XFILLER_35_905 VPWR VGND sg13g2_decap_8
XFILLER_47_787 VPWR VGND sg13g2_decap_8
XFILLER_43_971 VPWR VGND sg13g2_decap_8
XFILLER_15_640 VPWR VGND sg13g2_decap_8
XFILLER_30_654 VPWR VGND sg13g2_decap_8
X_3600_ _1114_ net581 _0999_ VPWR VGND sg13g2_nand2_1
X_3531_ net557 _1055_ _1056_ VPWR VGND sg13g2_nor2b_1
X_3462_ _0990_ _0991_ net611 _0992_ VPWR VGND sg13g2_nand3_1
X_2413_ _1834_ net734 _1642_ VPWR VGND sg13g2_nand2b_1
X_3393_ net12 net571 _0926_ VPWR VGND sg13g2_nor2_1
X_2344_ _1580_ VPWR _1765_ VGND _1677_ _1764_ sg13g2_o21ai_1
XFILLER_28_0 VPWR VGND sg13g2_fill_1
X_2275_ _1696_ _1681_ _1695_ _1680_ _1679_ VPWR VGND sg13g2_a22oi_1
XFILLER_38_732 VPWR VGND sg13g2_decap_8
X_4014_ _1425_ _1426_ _0191_ VPWR VGND sg13g2_and2_1
XFILLER_26_905 VPWR VGND sg13g2_decap_8
XFILLER_25_415 VPWR VGND sg13g2_decap_8
XFILLER_37_275 VPWR VGND sg13g2_fill_2
XFILLER_37_286 VPWR VGND sg13g2_fill_1
XFILLER_12_109 VPWR VGND sg13g2_fill_1
XFILLER_21_632 VPWR VGND sg13g2_decap_8
XFILLER_32_27 VPWR VGND sg13g2_fill_1
XFILLER_10_1007 VPWR VGND sg13g2_decap_8
X_3729_ net594 _0836_ _1209_ VPWR VGND sg13g2_nor2_1
XFILLER_0_547 VPWR VGND sg13g2_decap_8
XFILLER_48_507 VPWR VGND sg13g2_decap_8
XFILLER_44_724 VPWR VGND sg13g2_decap_8
XFILLER_17_927 VPWR VGND sg13g2_decap_8
XFILLER_29_776 VPWR VGND sg13g2_decap_8
XFILLER_16_448 VPWR VGND sg13g2_fill_1
XFILLER_24_470 VPWR VGND sg13g2_decap_8
XFILLER_25_982 VPWR VGND sg13g2_decap_8
XFILLER_40_963 VPWR VGND sg13g2_decap_8
XFILLER_8_636 VPWR VGND sg13g2_decap_8
XFILLER_7_102 VPWR VGND sg13g2_decap_8
XFILLER_12_665 VPWR VGND sg13g2_decap_8
XFILLER_4_831 VPWR VGND sg13g2_decap_8
XFILLER_26_1003 VPWR VGND sg13g2_decap_8
X_2060_ VPWR _1483_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_35_702 VPWR VGND sg13g2_decap_8
XFILLER_47_584 VPWR VGND sg13g2_decap_8
XFILLER_22_407 VPWR VGND sg13g2_fill_2
XFILLER_35_779 VPWR VGND sg13g2_decap_8
X_2962_ _0523_ VPWR _0525_ VGND net745 _0327_ sg13g2_o21ai_1
X_2893_ _0456_ _0447_ _0458_ VPWR VGND sg13g2_xor2_1
XFILLER_30_451 VPWR VGND sg13g2_fill_1
XFILLER_31_974 VPWR VGND sg13g2_decap_8
X_3514_ net557 _1040_ _1041_ _1042_ VPWR VGND sg13g2_nor3_1
X_3445_ net585 VPWR _0976_ VGND net612 _0975_ sg13g2_o21ai_1
X_3376_ _0909_ net588 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] net641
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2327_ _1514_ _1747_ _1748_ VPWR VGND sg13g2_and2_1
X_2258_ net707 _1609_ net706 _1678_ _1679_ VPWR VGND sg13g2_nor4_1
XFILLER_26_702 VPWR VGND sg13g2_decap_8
X_2189_ _1610_ _1506_ _1523_ VPWR VGND sg13g2_nand2_1
XFILLER_14_908 VPWR VGND sg13g2_decap_8
XFILLER_26_779 VPWR VGND sg13g2_decap_8
XFILLER_41_738 VPWR VGND sg13g2_decap_8
XFILLER_40_226 VPWR VGND sg13g2_fill_1
XFILLER_22_974 VPWR VGND sg13g2_decap_8
XFILLER_5_628 VPWR VGND sg13g2_decap_8
XFILLER_49_1025 VPWR VGND sg13g2_decap_4
XFILLER_0_311 VPWR VGND sg13g2_fill_2
XFILLER_1_856 VPWR VGND sg13g2_decap_8
XFILLER_29_573 VPWR VGND sg13g2_decap_8
XFILLER_44_521 VPWR VGND sg13g2_decap_8
XFILLER_17_724 VPWR VGND sg13g2_decap_8
XFILLER_44_598 VPWR VGND sg13g2_decap_8
XFILLER_32_749 VPWR VGND sg13g2_decap_8
XFILLER_9_901 VPWR VGND sg13g2_decap_8
XFILLER_40_760 VPWR VGND sg13g2_decap_8
XFILLER_13_985 VPWR VGND sg13g2_decap_8
XFILLER_9_978 VPWR VGND sg13g2_decap_8
X_3230_ _0758_ _0759_ _0764_ _0765_ _0766_ VPWR VGND sg13g2_and4_1
X_3161_ _1614_ net704 net714 _0697_ VPWR VGND sg13g2_nand3_1
X_2112_ sap_3_inst.controller.stage\[0\] net718 _1533_ VPWR VGND sg13g2_nor2b_2
XFILLER_48_871 VPWR VGND sg13g2_decap_8
X_3092_ _0628_ _1583_ _1579_ VPWR VGND sg13g2_nand2b_1
XFILLER_47_381 VPWR VGND sg13g2_decap_8
X_2043_ VPWR _1466_ sap_3_inst.alu.tmp\[5\] VGND sg13g2_inv_1
XFILLER_23_738 VPWR VGND sg13g2_decap_8
XFILLER_35_576 VPWR VGND sg13g2_decap_8
X_3994_ _1411_ u_ser.bit_pos\[1\] net767 VPWR VGND sg13g2_nand2_1
Xclkbuf_4_9_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_9_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2945_ VGND VPWR net748 _1466_ _0508_ _0487_ sg13g2_a21oi_1
XFILLER_31_771 VPWR VGND sg13g2_decap_8
X_2876_ net554 net753 _0441_ _0037_ VPWR VGND sg13g2_a21o_1
XFILLER_2_609 VPWR VGND sg13g2_decap_8
X_3428_ _0717_ VPWR _0960_ VGND net576 _0957_ sg13g2_o21ai_1
X_3359_ _0890_ _0891_ _0889_ _0893_ VPWR VGND _0892_ sg13g2_nand4_1
XFILLER_46_808 VPWR VGND sg13g2_decap_8
XFILLER_38_48 VPWR VGND sg13g2_fill_1
XFILLER_14_705 VPWR VGND sg13g2_decap_8
XFILLER_26_576 VPWR VGND sg13g2_decap_8
XFILLER_41_535 VPWR VGND sg13g2_decap_8
XFILLER_13_237 VPWR VGND sg13g2_fill_2
XFILLER_22_771 VPWR VGND sg13g2_decap_8
XFILLER_10_944 VPWR VGND sg13g2_decap_8
XFILLER_6_904 VPWR VGND sg13g2_decap_8
XFILLER_1_653 VPWR VGND sg13g2_decap_8
XFILLER_0_152 VPWR VGND sg13g2_decap_8
XFILLER_49_668 VPWR VGND sg13g2_decap_8
XFILLER_17_521 VPWR VGND sg13g2_decap_8
XFILLER_45_863 VPWR VGND sg13g2_decap_8
XFILLER_17_598 VPWR VGND sg13g2_decap_8
XFILLER_44_395 VPWR VGND sg13g2_decap_8
XFILLER_32_546 VPWR VGND sg13g2_decap_8
X_2730_ _1546_ _1718_ _0299_ VPWR VGND sg13g2_nor2_1
XFILLER_13_782 VPWR VGND sg13g2_decap_8
X_2661_ _0251_ VPWR _0255_ VGND _1954_ _0254_ sg13g2_o21ai_1
XFILLER_9_775 VPWR VGND sg13g2_decap_8
X_2592_ net745 net743 _2002_ VPWR VGND sg13g2_xor2_1
XFILLER_5_992 VPWR VGND sg13g2_decap_8
X_3213_ _0749_ net587 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] net592
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4193_ net787 VGND VPWR _0171_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3144_ VGND VPWR net695 _1703_ _0680_ _1588_ sg13g2_a21oi_1
X_3075_ _0273_ VPWR _0611_ VGND net700 _1704_ sg13g2_o21ai_1
X_2026_ VPWR _1449_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_35_340 VPWR VGND sg13g2_fill_2
XFILLER_36_885 VPWR VGND sg13g2_decap_8
XFILLER_39_1013 VPWR VGND sg13g2_decap_8
XFILLER_23_535 VPWR VGND sg13g2_decap_8
X_3977_ _0431_ net664 _1399_ VPWR VGND sg13g2_nor2_1
X_2928_ _0492_ _0452_ _0491_ VPWR VGND sg13g2_nand2b_1
X_2859_ _0425_ _0422_ _0424_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
Xfanout721 _1314_ net721 VPWR VGND sg13g2_buf_8
Xfanout710 _1556_ net710 VPWR VGND sg13g2_buf_8
Xfanout732 sap_3_inst.controller.opcode\[4\] net732 VPWR VGND sg13g2_buf_8
Xfanout776 net777 net776 VPWR VGND sg13g2_buf_8
Xfanout765 _1280_ net765 VPWR VGND sg13g2_buf_8
Xfanout754 sap_3_inst.alu.acc\[3\] net754 VPWR VGND sg13g2_buf_8
Xfanout743 net744 net743 VPWR VGND sg13g2_buf_8
XFILLER_46_605 VPWR VGND sg13g2_decap_8
Xfanout787 net792 net787 VPWR VGND sg13g2_buf_2
Xfanout798 net800 net798 VPWR VGND sg13g2_buf_8
XFILLER_27_830 VPWR VGND sg13g2_decap_8
XFILLER_45_159 VPWR VGND sg13g2_fill_1
XFILLER_42_811 VPWR VGND sg13g2_decap_8
XFILLER_14_502 VPWR VGND sg13g2_decap_8
XFILLER_42_888 VPWR VGND sg13g2_decap_8
XFILLER_14_579 VPWR VGND sg13g2_decap_8
XFILLER_6_701 VPWR VGND sg13g2_decap_8
XFILLER_10_741 VPWR VGND sg13g2_decap_8
XFILLER_5_200 VPWR VGND sg13g2_fill_1
XFILLER_6_778 VPWR VGND sg13g2_decap_8
XFILLER_7_1000 VPWR VGND sg13g2_decap_8
XFILLER_2_973 VPWR VGND sg13g2_decap_8
XFILLER_1_450 VPWR VGND sg13g2_decap_8
XFILLER_49_465 VPWR VGND sg13g2_decap_8
XFILLER_18_852 VPWR VGND sg13g2_decap_8
XFILLER_45_660 VPWR VGND sg13g2_decap_8
XFILLER_17_351 VPWR VGND sg13g2_fill_2
X_3900_ _1339_ net761 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] net721
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_844 VPWR VGND sg13g2_decap_8
X_3831_ _0154_ _1125_ _1279_ net602 _1491_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_527 VPWR VGND sg13g2_decap_8
X_3762_ _1231_ _0844_ _0918_ _1230_ VPWR VGND sg13g2_and3_1
X_2713_ _0290_ _0291_ _0287_ _0292_ VPWR VGND sg13g2_nand3_1
XFILLER_9_572 VPWR VGND sg13g2_decap_8
X_3693_ _1050_ _1181_ _1187_ VPWR VGND sg13g2_nor2_1
X_2644_ _0239_ net1 _1847_ VPWR VGND sg13g2_nand2_1
X_2575_ _1986_ _1982_ _1985_ net637 _1444_ VPWR VGND sg13g2_a22oi_1
X_4176_ net777 VGND VPWR _0154_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[7\]
+ clknet_5_3__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3127_ net724 _1510_ net734 _0663_ VPWR VGND net697 sg13g2_nand4_1
XFILLER_28_638 VPWR VGND sg13g2_decap_8
X_3058_ _0596_ net727 net691 VPWR VGND sg13g2_nand2_1
XFILLER_36_682 VPWR VGND sg13g2_decap_8
XFILLER_42_129 VPWR VGND sg13g2_fill_2
X_2009_ VPWR _1432_ u_ser.state\[0\] VGND sg13g2_inv_1
XFILLER_24_855 VPWR VGND sg13g2_decap_8
XFILLER_13_1027 VPWR VGND sg13g2_fill_2
XFILLER_3_759 VPWR VGND sg13g2_decap_8
Xfanout551 _1126_ net551 VPWR VGND sg13g2_buf_2
Xfanout573 _0338_ net573 VPWR VGND sg13g2_buf_8
Xfanout562 _0716_ net562 VPWR VGND sg13g2_buf_8
Xfanout584 net586 net584 VPWR VGND sg13g2_buf_8
XFILLER_46_402 VPWR VGND sg13g2_decap_8
XFILLER_19_649 VPWR VGND sg13g2_decap_8
Xfanout595 _0734_ net595 VPWR VGND sg13g2_buf_8
XFILLER_47_969 VPWR VGND sg13g2_decap_8
XFILLER_46_479 VPWR VGND sg13g2_decap_8
XFILLER_15_822 VPWR VGND sg13g2_decap_8
XFILLER_14_354 VPWR VGND sg13g2_fill_1
XFILLER_42_685 VPWR VGND sg13g2_decap_8
XFILLER_15_899 VPWR VGND sg13g2_decap_8
XFILLER_30_836 VPWR VGND sg13g2_decap_8
XFILLER_6_575 VPWR VGND sg13g2_decap_8
X_2360_ net734 net731 _1781_ VPWR VGND sg13g2_and2_1
X_2291_ net722 _1564_ _1712_ VPWR VGND sg13g2_nor2_1
XFILLER_2_770 VPWR VGND sg13g2_decap_8
XFILLER_38_914 VPWR VGND sg13g2_decap_8
XFILLER_21_814 VPWR VGND sg13g2_decap_8
XFILLER_32_140 VPWR VGND sg13g2_fill_2
XFILLER_33_641 VPWR VGND sg13g2_decap_8
X_3814_ _1267_ net607 net12 VPWR VGND sg13g2_nand2b_1
X_3745_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] _1195_ _1211_ _0130_
+ VPWR VGND sg13g2_mux2_1
X_3676_ net574 _1172_ _1173_ VPWR VGND sg13g2_nor2_1
X_2627_ VGND VPWR _1723_ _0213_ _0224_ _0223_ sg13g2_a21oi_1
XFILLER_0_729 VPWR VGND sg13g2_decap_8
X_2558_ _1971_ net626 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] net628
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2489_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] net638
+ net621 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] _1904_ net623 sg13g2_a221oi_1
XFILLER_44_906 VPWR VGND sg13g2_decap_8
X_4159_ net781 VGND VPWR _0137_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\]
+ clknet_5_13__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_28_435 VPWR VGND sg13g2_decap_8
XFILLER_29_958 VPWR VGND sg13g2_decap_8
XFILLER_24_652 VPWR VGND sg13g2_decap_8
XFILLER_12_847 VPWR VGND sg13g2_decap_8
XFILLER_23_151 VPWR VGND sg13g2_fill_1
XFILLER_8_818 VPWR VGND sg13g2_decap_8
XFILLER_20_891 VPWR VGND sg13g2_decap_8
XFILLER_3_556 VPWR VGND sg13g2_decap_8
XFILLER_47_766 VPWR VGND sg13g2_decap_8
XFILLER_19_424 VPWR VGND sg13g2_fill_1
XFILLER_34_416 VPWR VGND sg13g2_fill_1
XFILLER_43_950 VPWR VGND sg13g2_decap_8
XFILLER_42_482 VPWR VGND sg13g2_decap_8
XFILLER_15_696 VPWR VGND sg13g2_decap_8
XFILLER_30_633 VPWR VGND sg13g2_decap_8
X_3530_ _1055_ net580 VPWR VGND _0924_ sg13g2_nand2b_2
XFILLER_7_895 VPWR VGND sg13g2_decap_8
X_3461_ _0991_ net644 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] net647
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2412_ _1833_ net686 _1832_ VPWR VGND sg13g2_nand2_1
X_3392_ _0925_ _0717_ _0921_ VPWR VGND sg13g2_nand2_1
X_2343_ _1593_ _1597_ _1590_ _1764_ VPWR VGND sg13g2_nand3_1
X_4013_ _1424_ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\] net768 _1426_
+ VPWR VGND sg13g2_a21o_1
X_2274_ _1663_ _1683_ _1684_ _1694_ _1695_ VPWR VGND sg13g2_nor4_1
XFILLER_38_711 VPWR VGND sg13g2_decap_8
XFILLER_37_210 VPWR VGND sg13g2_fill_1
XFILLER_38_788 VPWR VGND sg13g2_decap_8
XFILLER_21_611 VPWR VGND sg13g2_decap_8
XFILLER_21_688 VPWR VGND sg13g2_decap_8
X_3728_ _0122_ _1125_ _1208_ net594 _1494_ VPWR VGND sg13g2_a22oi_1
X_3659_ VGND VPWR net584 _1155_ _1159_ _1158_ sg13g2_a21oi_1
XFILLER_0_526 VPWR VGND sg13g2_decap_8
XFILLER_29_755 VPWR VGND sg13g2_decap_8
XFILLER_44_703 VPWR VGND sg13g2_decap_8
XFILLER_17_906 VPWR VGND sg13g2_decap_8
XFILLER_25_961 VPWR VGND sg13g2_decap_8
XFILLER_40_942 VPWR VGND sg13g2_decap_8
XFILLER_12_644 VPWR VGND sg13g2_decap_8
XFILLER_8_615 VPWR VGND sg13g2_decap_8
XFILLER_4_810 VPWR VGND sg13g2_decap_8
XFILLER_4_887 VPWR VGND sg13g2_decap_8
XFILLER_3_364 VPWR VGND sg13g2_fill_1
XFILLER_47_563 VPWR VGND sg13g2_decap_8
XFILLER_35_758 VPWR VGND sg13g2_decap_8
X_2961_ _0522_ VPWR _0524_ VGND _0505_ _0520_ sg13g2_o21ai_1
XFILLER_31_953 VPWR VGND sg13g2_decap_8
X_2892_ VGND VPWR _0457_ _0456_ _0447_ sg13g2_or2_1
XFILLER_33_1019 VPWR VGND sg13g2_decap_8
XFILLER_7_692 VPWR VGND sg13g2_decap_8
X_3513_ net561 net575 _1041_ VPWR VGND sg13g2_nor2_2
X_3444_ _0824_ _0974_ _0975_ VPWR VGND sg13g2_and2_1
XFILLER_40_0 VPWR VGND sg13g2_fill_1
X_3375_ _0908_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[3\] _0716_ VPWR
+ VGND sg13g2_nand2_1
X_2326_ net709 net684 net741 _1747_ VPWR VGND sg13g2_nand3_1
X_2257_ _1678_ _1593_ _1597_ VPWR VGND sg13g2_nand2_1
X_2188_ _1507_ net722 _1609_ VPWR VGND sg13g2_nor2_2
XFILLER_38_585 VPWR VGND sg13g2_decap_8
XFILLER_26_758 VPWR VGND sg13g2_decap_8
XFILLER_41_717 VPWR VGND sg13g2_decap_8
XFILLER_22_953 VPWR VGND sg13g2_decap_8
XFILLER_21_485 VPWR VGND sg13g2_decap_8
XFILLER_5_607 VPWR VGND sg13g2_decap_8
XFILLER_49_1004 VPWR VGND sg13g2_decap_8
XFILLER_1_835 VPWR VGND sg13g2_decap_8
XFILLER_17_703 VPWR VGND sg13g2_decap_8
XFILLER_29_552 VPWR VGND sg13g2_decap_8
XFILLER_44_500 VPWR VGND sg13g2_decap_8
XFILLER_1_1017 VPWR VGND sg13g2_decap_8
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_44_577 VPWR VGND sg13g2_decap_8
XFILLER_16_279 VPWR VGND sg13g2_fill_1
XFILLER_32_728 VPWR VGND sg13g2_decap_8
XFILLER_13_964 VPWR VGND sg13g2_decap_8
XFILLER_9_957 VPWR VGND sg13g2_decap_8
XFILLER_4_684 VPWR VGND sg13g2_decap_8
X_3160_ VGND VPWR _0618_ _0666_ _0696_ net686 sg13g2_a21oi_1
X_3091_ net700 _1712_ net735 _0627_ VPWR VGND sg13g2_nand3_1
XFILLER_0_890 VPWR VGND sg13g2_decap_8
X_2111_ _1532_ _1499_ _1531_ VPWR VGND sg13g2_nand2_1
Xhold1 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[0\] VPWR VGND net48 sg13g2_dlygate4sd3_1
XFILLER_48_850 VPWR VGND sg13g2_decap_8
X_2042_ VPWR _1465_ sap_3_inst.alu.tmp\[3\] VGND sg13g2_inv_1
XFILLER_47_360 VPWR VGND sg13g2_decap_8
XFILLER_35_555 VPWR VGND sg13g2_decap_8
XFILLER_23_717 VPWR VGND sg13g2_decap_8
X_3993_ u_ser.state\[0\] _1433_ _1410_ VPWR VGND sg13g2_nor2_2
X_2944_ _0505_ _0506_ _0507_ VPWR VGND sg13g2_nor2b_2
XFILLER_31_750 VPWR VGND sg13g2_decap_8
X_2875_ VPWR VGND _0440_ net554 _0439_ net546 _0441_ net616 sg13g2_a221oi_1
XFILLER_1_109 VPWR VGND sg13g2_fill_1
X_3427_ VPWR _0959_ _0958_ VGND sg13g2_inv_1
X_3358_ _0892_ net588 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] net641
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2309_ _1655_ VPWR _1730_ VGND net697 net684 sg13g2_o21ai_1
X_3289_ _0757_ _0766_ _0775_ _0823_ _0825_ VPWR VGND sg13g2_and4_1
XFILLER_39_894 VPWR VGND sg13g2_decap_8
XFILLER_26_555 VPWR VGND sg13g2_decap_8
XFILLER_41_514 VPWR VGND sg13g2_decap_8
XFILLER_22_750 VPWR VGND sg13g2_decap_8
XFILLER_10_923 VPWR VGND sg13g2_decap_8
XFILLER_1_632 VPWR VGND sg13g2_decap_8
XFILLER_49_647 VPWR VGND sg13g2_decap_8
XFILLER_23_1018 VPWR VGND sg13g2_decap_8
XFILLER_45_842 VPWR VGND sg13g2_decap_8
XFILLER_17_577 VPWR VGND sg13g2_decap_8
XFILLER_32_525 VPWR VGND sg13g2_decap_8
XFILLER_13_761 VPWR VGND sg13g2_decap_8
XFILLER_20_709 VPWR VGND sg13g2_decap_8
XFILLER_9_754 VPWR VGND sg13g2_decap_8
X_2660_ _0254_ _0252_ _0253_ VPWR VGND sg13g2_nand2_1
XFILLER_5_20 VPWR VGND sg13g2_decap_8
X_2591_ _2001_ _1999_ _2000_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_971 VPWR VGND sg13g2_decap_8
XFILLER_4_481 VPWR VGND sg13g2_decap_8
X_3212_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\] _0747_
+ net658 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] _0748_ net606 sg13g2_a221oi_1
X_4192_ net796 VGND VPWR _0170_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\]
+ clknet_5_29__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_39_102 VPWR VGND sg13g2_fill_1
X_3143_ VGND VPWR _0273_ _0678_ _0679_ _0677_ sg13g2_a21oi_1
XFILLER_39_168 VPWR VGND sg13g2_fill_2
X_3074_ _1830_ _0298_ _0610_ VPWR VGND _0609_ sg13g2_nand3b_1
X_2025_ VPWR _1448_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_36_864 VPWR VGND sg13g2_decap_8
XFILLER_23_514 VPWR VGND sg13g2_decap_8
X_3976_ _1398_ sap_3_inst.alu.act\[2\] net548 _0180_ VPWR VGND sg13g2_mux2_1
X_2927_ _0490_ _0479_ _0491_ VPWR VGND sg13g2_xor2_1
X_2858_ VGND VPWR net755 sap_3_inst.alu.tmp\[2\] _0424_ _0384_ sg13g2_a21oi_1
X_2789_ _0355_ _0356_ _0357_ VPWR VGND sg13g2_nor2b_1
XFILLER_46_1018 VPWR VGND sg13g2_decap_8
Xfanout700 net701 net700 VPWR VGND sg13g2_buf_8
Xfanout722 _1524_ net722 VPWR VGND sg13g2_buf_8
Xfanout711 _1531_ net711 VPWR VGND sg13g2_buf_8
Xfanout733 net734 net733 VPWR VGND sg13g2_buf_8
Xfanout755 net756 net755 VPWR VGND sg13g2_buf_8
Xfanout766 _0186_ net766 VPWR VGND sg13g2_buf_8
Xfanout744 sap_3_inst.alu.acc\[7\] net744 VPWR VGND sg13g2_buf_8
Xfanout777 net778 net777 VPWR VGND sg13g2_buf_8
Xfanout799 net800 net799 VPWR VGND sg13g2_buf_8
Xfanout788 net792 net788 VPWR VGND sg13g2_buf_8
XFILLER_39_691 VPWR VGND sg13g2_decap_8
XFILLER_27_886 VPWR VGND sg13g2_decap_8
Xclkbuf_5_29__f_sap_3_inst.alu.clk_regs clknet_4_14_0_sap_3_inst.alu.clk_regs clknet_5_29__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_42_867 VPWR VGND sg13g2_decap_8
XFILLER_41_355 VPWR VGND sg13g2_fill_1
XFILLER_14_558 VPWR VGND sg13g2_decap_8
XFILLER_10_720 VPWR VGND sg13g2_decap_8
XFILLER_10_797 VPWR VGND sg13g2_decap_8
XFILLER_6_757 VPWR VGND sg13g2_decap_8
XFILLER_2_952 VPWR VGND sg13g2_decap_8
XFILLER_49_444 VPWR VGND sg13g2_decap_8
XFILLER_37_639 VPWR VGND sg13g2_decap_8
XFILLER_18_831 VPWR VGND sg13g2_decap_8
XFILLER_33_823 VPWR VGND sg13g2_decap_8
X_3830_ VGND VPWR _1276_ _1278_ _1279_ net602 sg13g2_a21oi_1
XFILLER_20_506 VPWR VGND sg13g2_decap_8
X_3761_ _0916_ VPWR _1230_ VGND _0873_ _0894_ sg13g2_o21ai_1
X_2712_ _1602_ _0289_ _1580_ _0291_ VPWR VGND sg13g2_nand3_1
XFILLER_9_551 VPWR VGND sg13g2_decap_8
X_3692_ _1181_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] _1186_ _0108_
+ VPWR VGND sg13g2_a21o_1
X_2643_ _0238_ _1828_ sap_3_inst.alu.flags\[0\] _1827_ net760 VPWR VGND sg13g2_a22oi_1
X_2574_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] _1984_
+ net628 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[2\] _1985_ net630 sg13g2_a221oi_1
X_4175_ net780 VGND VPWR _0153_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\]
+ clknet_5_13__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3126_ _0662_ _1601_ _1690_ VPWR VGND sg13g2_nand2_1
XFILLER_28_617 VPWR VGND sg13g2_decap_8
X_3057_ _0595_ VPWR _0064_ VGND net691 _1899_ sg13g2_o21ai_1
XFILLER_36_661 VPWR VGND sg13g2_decap_8
XFILLER_23_311 VPWR VGND sg13g2_fill_2
XFILLER_24_834 VPWR VGND sg13g2_decap_8
X_3959_ _1387_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] net602 VPWR
+ VGND sg13g2_nand2_1
XFILLER_13_1006 VPWR VGND sg13g2_decap_8
XFILLER_3_738 VPWR VGND sg13g2_decap_8
Xfanout563 _0330_ net563 VPWR VGND sg13g2_buf_8
Xfanout574 _0845_ net574 VPWR VGND sg13g2_buf_8
Xfanout552 _0944_ net552 VPWR VGND sg13g2_buf_8
XFILLER_47_948 VPWR VGND sg13g2_decap_8
Xfanout596 net597 net596 VPWR VGND sg13g2_buf_8
Xfanout585 net586 net585 VPWR VGND sg13g2_buf_1
XFILLER_19_628 VPWR VGND sg13g2_decap_8
XFILLER_46_458 VPWR VGND sg13g2_decap_8
XFILLER_15_801 VPWR VGND sg13g2_decap_8
XFILLER_14_300 VPWR VGND sg13g2_fill_2
XFILLER_27_683 VPWR VGND sg13g2_decap_8
XFILLER_42_664 VPWR VGND sg13g2_decap_8
XFILLER_15_878 VPWR VGND sg13g2_decap_8
XFILLER_25_83 VPWR VGND sg13g2_fill_1
XFILLER_30_815 VPWR VGND sg13g2_decap_8
XFILLER_6_554 VPWR VGND sg13g2_decap_8
XFILLER_10_594 VPWR VGND sg13g2_decap_8
X_2290_ _1650_ _1702_ _1706_ _1710_ _1711_ VPWR VGND sg13g2_and4_1
XFILLER_33_620 VPWR VGND sg13g2_decap_8
X_3813_ _1266_ net604 _0935_ VPWR VGND sg13g2_nand2_1
XFILLER_33_697 VPWR VGND sg13g2_decap_8
X_3744_ VGND VPWR _1484_ _1210_ _0129_ _1217_ sg13g2_a21oi_1
X_3675_ net606 _1032_ _1172_ VPWR VGND sg13g2_nor2_1
X_2626_ VGND VPWR _0218_ _0222_ _0223_ net567 sg13g2_a21oi_1
XFILLER_0_708 VPWR VGND sg13g2_decap_8
X_2557_ _1970_ net620 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\] net630
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2488_ _1901_ _1902_ _1903_ VPWR VGND sg13g2_and2_1
X_4227_ regFile_serial_start net30 VPWR VGND sg13g2_buf_8
XFILLER_29_937 VPWR VGND sg13g2_decap_8
X_4158_ net775 VGND VPWR _0136_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\]
+ clknet_5_10__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3109_ net686 VPWR _0645_ VGND _1590_ _0638_ sg13g2_o21ai_1
X_4089_ net782 VGND VPWR _0067_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[0\]
+ clknet_5_6__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_1
XFILLER_43_439 VPWR VGND sg13g2_decap_8
XFILLER_24_631 VPWR VGND sg13g2_decap_8
XFILLER_12_826 VPWR VGND sg13g2_decap_8
XFILLER_20_870 VPWR VGND sg13g2_decap_8
XFILLER_3_535 VPWR VGND sg13g2_decap_8
XFILLER_11_63 VPWR VGND sg13g2_fill_1
XFILLER_47_745 VPWR VGND sg13g2_decap_8
XFILLER_46_277 VPWR VGND sg13g2_fill_2
XFILLER_27_480 VPWR VGND sg13g2_decap_8
XFILLER_28_981 VPWR VGND sg13g2_decap_8
XFILLER_42_461 VPWR VGND sg13g2_decap_8
XFILLER_14_141 VPWR VGND sg13g2_fill_1
XFILLER_15_675 VPWR VGND sg13g2_decap_8
XFILLER_30_612 VPWR VGND sg13g2_decap_8
XFILLER_30_689 VPWR VGND sg13g2_decap_8
XFILLER_7_874 VPWR VGND sg13g2_decap_8
XFILLER_10_391 VPWR VGND sg13g2_fill_2
X_3460_ _0990_ net649 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\] net654
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2411_ _1639_ _1661_ net733 _1832_ VPWR VGND sg13g2_nand3_1
X_3391_ _0922_ _0923_ _0924_ VPWR VGND sg13g2_and2_1
X_2342_ _1763_ _1623_ _1578_ _1598_ _1588_ VPWR VGND sg13g2_a22oi_1
X_4012_ sap_3_inst.reg_file.array_serializer_inst.word_index\[1\] _1424_ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\]
+ _1425_ VPWR VGND sg13g2_nand3_1
XFILLER_42_1021 VPWR VGND sg13g2_decap_8
X_2273_ _1686_ _1689_ _1685_ _1694_ VPWR VGND _1693_ sg13g2_nand4_1
XFILLER_38_767 VPWR VGND sg13g2_decap_8
XFILLER_19_992 VPWR VGND sg13g2_decap_8
XFILLER_37_277 VPWR VGND sg13g2_fill_1
XFILLER_34_984 VPWR VGND sg13g2_decap_8
XFILLER_21_667 VPWR VGND sg13g2_decap_8
X_3727_ net594 _1194_ _1208_ VPWR VGND sg13g2_nor2_1
X_3658_ net584 _1157_ _1158_ VPWR VGND sg13g2_nor2_1
X_3589_ _1104_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] net591 VPWR
+ VGND sg13g2_nand2_1
X_2609_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] net624 _0206_ VPWR
+ VGND sg13g2_and2_1
XFILLER_0_505 VPWR VGND sg13g2_decap_8
XFILLER_29_734 VPWR VGND sg13g2_decap_8
XFILLER_44_759 VPWR VGND sg13g2_decap_8
XFILLER_25_940 VPWR VGND sg13g2_decap_8
XFILLER_40_921 VPWR VGND sg13g2_decap_8
XFILLER_12_623 VPWR VGND sg13g2_decap_8
XFILLER_40_998 VPWR VGND sg13g2_decap_8
XFILLER_4_866 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_39_509 VPWR VGND sg13g2_decap_8
XFILLER_47_542 VPWR VGND sg13g2_decap_8
XFILLER_35_737 VPWR VGND sg13g2_decap_8
X_2960_ VGND VPWR _0523_ _0510_ _0323_ sg13g2_or2_1
XFILLER_15_461 VPWR VGND sg13g2_fill_2
XFILLER_16_984 VPWR VGND sg13g2_decap_8
XFILLER_22_409 VPWR VGND sg13g2_fill_1
X_2891_ VGND VPWR net754 _1465_ _0456_ _0430_ sg13g2_a21oi_1
XFILLER_31_932 VPWR VGND sg13g2_decap_8
XFILLER_8_42 VPWR VGND sg13g2_decap_4
Xclkbuf_5_3__f_sap_3_inst.alu.clk_regs clknet_4_1_0_sap_3_inst.alu.clk_regs clknet_5_3__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_8_64 VPWR VGND sg13g2_fill_1
XFILLER_30_486 VPWR VGND sg13g2_decap_8
XFILLER_7_671 VPWR VGND sg13g2_decap_8
X_3512_ net31 _0846_ _1039_ _1040_ VPWR VGND sg13g2_nor3_2
X_3443_ _0823_ _0775_ _0766_ _0974_ VPWR VGND sg13g2_a21o_1
X_3374_ _0905_ VPWR _0069_ VGND net562 _0901_ sg13g2_o21ai_1
X_2325_ VPWR VGND net712 _1745_ _1743_ _1741_ _1746_ _1742_ sg13g2_a221oi_1
X_2256_ _1604_ VPWR _1677_ VGND _1438_ _1610_ sg13g2_o21ai_1
XFILLER_38_564 VPWR VGND sg13g2_decap_8
X_2187_ _1608_ _1604_ _1606_ VPWR VGND sg13g2_nand2_1
XFILLER_26_737 VPWR VGND sg13g2_decap_8
XFILLER_25_258 VPWR VGND sg13g2_fill_2
XFILLER_22_932 VPWR VGND sg13g2_decap_8
XFILLER_34_781 VPWR VGND sg13g2_decap_8
XFILLER_1_814 VPWR VGND sg13g2_decap_8
XFILLER_49_829 VPWR VGND sg13g2_decap_8
XFILLER_48_339 VPWR VGND sg13g2_decap_8
XFILLER_29_531 VPWR VGND sg13g2_decap_8
XFILLER_44_556 VPWR VGND sg13g2_decap_8
XFILLER_17_759 VPWR VGND sg13g2_decap_8
XFILLER_32_707 VPWR VGND sg13g2_decap_8
XFILLER_12_420 VPWR VGND sg13g2_fill_2
XFILLER_13_943 VPWR VGND sg13g2_decap_8
Xclkbuf_5_10__f_sap_3_inst.alu.clk_regs clknet_4_5_0_sap_3_inst.alu.clk_regs clknet_5_10__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_9_936 VPWR VGND sg13g2_decap_8
XFILLER_12_453 VPWR VGND sg13g2_fill_1
XFILLER_40_795 VPWR VGND sg13g2_decap_8
XFILLER_4_663 VPWR VGND sg13g2_decap_8
X_3090_ net707 _0273_ _0626_ VPWR VGND sg13g2_nor2_1
X_2110_ net718 net719 _1531_ VPWR VGND sg13g2_nor2b_2
Xhold2 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[4\] VPWR VGND net49 sg13g2_dlygate4sd3_1
X_2041_ VPWR _1464_ sap_3_inst.alu.tmp\[2\] VGND sg13g2_inv_1
XFILLER_35_534 VPWR VGND sg13g2_decap_8
X_3992_ _1407_ VPWR _0185_ VGND net549 _1409_ sg13g2_o21ai_1
X_2943_ _0506_ net745 sap_3_inst.alu.tmp\[6\] VPWR VGND sg13g2_nand2_2
XFILLER_16_781 VPWR VGND sg13g2_decap_8
X_2874_ VGND VPWR sap_3_inst.alu.act\[3\] net669 _0440_ net616 sg13g2_a21oi_1
X_3426_ _0958_ _0922_ _0775_ _0852_ _0797_ VPWR VGND sg13g2_a22oi_1
X_3357_ _0891_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] net592 VPWR
+ VGND sg13g2_nand2_1
X_2308_ _1729_ net706 _1727_ VPWR VGND sg13g2_nand2b_1
X_3288_ _0775_ _0823_ _0766_ _0824_ VPWR VGND sg13g2_nand3_1
X_2239_ _1655_ net687 _1657_ _1660_ VPWR VGND sg13g2_a21o_1
XFILLER_39_873 VPWR VGND sg13g2_decap_8
XFILLER_26_534 VPWR VGND sg13g2_decap_8
XFILLER_13_239 VPWR VGND sg13g2_fill_1
XFILLER_10_902 VPWR VGND sg13g2_decap_8
XFILLER_16_1026 VPWR VGND sg13g2_fill_2
XFILLER_10_979 VPWR VGND sg13g2_decap_8
XFILLER_6_939 VPWR VGND sg13g2_decap_8
XFILLER_5_438 VPWR VGND sg13g2_fill_2
XFILLER_1_611 VPWR VGND sg13g2_decap_8
XFILLER_0_110 VPWR VGND sg13g2_fill_2
XFILLER_0_132 VPWR VGND sg13g2_decap_8
XFILLER_49_626 VPWR VGND sg13g2_decap_8
XFILLER_1_688 VPWR VGND sg13g2_decap_8
XFILLER_45_821 VPWR VGND sg13g2_decap_8
XFILLER_17_556 VPWR VGND sg13g2_decap_8
XFILLER_45_898 VPWR VGND sg13g2_decap_8
XFILLER_32_504 VPWR VGND sg13g2_decap_8
XFILLER_13_740 VPWR VGND sg13g2_decap_8
XFILLER_9_733 VPWR VGND sg13g2_decap_8
XFILLER_40_592 VPWR VGND sg13g2_decap_8
XFILLER_5_950 VPWR VGND sg13g2_decap_8
X_2590_ net756 net754 _2000_ VPWR VGND sg13g2_xor2_1
XFILLER_4_460 VPWR VGND sg13g2_decap_8
XFILLER_5_87 VPWR VGND sg13g2_fill_1
X_3211_ _0747_ _0745_ _0746_ VPWR VGND sg13g2_nand2_1
X_4191_ net800 VGND VPWR _0169_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[7\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
X_3142_ _1627_ _1703_ net694 _0678_ VPWR VGND _0675_ sg13g2_nand4_1
X_3073_ VGND VPWR _1515_ _0608_ _0609_ net713 sg13g2_a21oi_1
X_2024_ VPWR _1447_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_36_843 VPWR VGND sg13g2_decap_8
X_3975_ _0391_ net755 net663 _1398_ VPWR VGND sg13g2_mux2_1
X_2926_ VGND VPWR net750 sap_3_inst.alu.tmp\[4\] _0490_ _0449_ sg13g2_a21oi_1
X_2857_ VPWR _0423_ _0422_ VGND sg13g2_inv_1
X_2788_ _0356_ sap_3_inst.alu.tmp\[0\] net759 VPWR VGND sg13g2_nand2b_1
X_3409_ _0941_ net587 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] net640
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] VPWR VGND sg13g2_a22oi_1
Xfanout723 net724 net723 VPWR VGND sg13g2_buf_8
Xfanout701 _1529_ net701 VPWR VGND sg13g2_buf_2
Xfanout712 _1514_ net712 VPWR VGND sg13g2_buf_8
Xfanout767 u_ser.bit_pos\[0\] net767 VPWR VGND sg13g2_buf_8
Xfanout756 sap_3_inst.alu.acc\[2\] net756 VPWR VGND sg13g2_buf_8
Xfanout745 net746 net745 VPWR VGND sg13g2_buf_8
Xfanout734 sap_3_inst.controller.opcode\[3\] net734 VPWR VGND sg13g2_buf_8
Xfanout789 net792 net789 VPWR VGND sg13g2_buf_8
Xfanout778 net801 net778 VPWR VGND sg13g2_buf_8
Xclkbuf_4_10_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_10_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_39_670 VPWR VGND sg13g2_decap_8
XFILLER_27_865 VPWR VGND sg13g2_decap_8
XFILLER_42_846 VPWR VGND sg13g2_decap_8
XFILLER_14_537 VPWR VGND sg13g2_decap_8
XFILLER_41_367 VPWR VGND sg13g2_decap_4
XFILLER_6_736 VPWR VGND sg13g2_decap_8
XFILLER_5_213 VPWR VGND sg13g2_fill_1
XFILLER_10_776 VPWR VGND sg13g2_decap_8
XFILLER_30_40 VPWR VGND sg13g2_fill_1
XFILLER_2_931 VPWR VGND sg13g2_decap_8
XFILLER_30_95 VPWR VGND sg13g2_fill_1
XFILLER_49_423 VPWR VGND sg13g2_decap_8
XFILLER_1_485 VPWR VGND sg13g2_decap_8
XFILLER_39_71 VPWR VGND sg13g2_fill_1
XFILLER_18_810 VPWR VGND sg13g2_decap_8
XFILLER_37_618 VPWR VGND sg13g2_decap_8
XFILLER_18_887 VPWR VGND sg13g2_decap_8
XFILLER_33_802 VPWR VGND sg13g2_decap_8
XFILLER_45_695 VPWR VGND sg13g2_decap_8
XFILLER_32_312 VPWR VGND sg13g2_fill_2
XFILLER_33_879 VPWR VGND sg13g2_decap_8
X_3760_ _0133_ _0899_ _1229_ net599 _1448_ VPWR VGND sg13g2_a22oi_1
X_2711_ _0290_ _0288_ _1709_ _0286_ _1677_ VPWR VGND sg13g2_a22oi_1
XFILLER_9_530 VPWR VGND sg13g2_decap_8
X_3691_ _1181_ _1184_ _1185_ _1186_ VPWR VGND sg13g2_nor3_1
X_2642_ _1723_ _0236_ _0237_ VPWR VGND sg13g2_and2_1
X_2573_ _1984_ _1980_ _1983_ VPWR VGND sg13g2_nand2_1
X_4174_ net777 VGND VPWR _0152_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\]
+ clknet_5_8__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3125_ net733 VPWR _0661_ VGND _1749_ _1814_ sg13g2_o21ai_1
XFILLER_49_990 VPWR VGND sg13g2_decap_8
X_3056_ _0595_ net729 net691 VPWR VGND sg13g2_nand2_1
XFILLER_24_813 VPWR VGND sg13g2_decap_8
XFILLER_36_640 VPWR VGND sg13g2_decap_8
XFILLER_35_172 VPWR VGND sg13g2_fill_1
XFILLER_11_529 VPWR VGND sg13g2_decap_8
X_3958_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[4\] _1188_ net607 _0174_
+ VPWR VGND sg13g2_mux2_1
Xclkbuf_4_2_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_2_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2909_ net671 net747 _0473_ VPWR VGND sg13g2_xor2_1
X_3889_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] _1305_
+ _1329_ net762 sg13g2_a21oi_1
XFILLER_3_717 VPWR VGND sg13g2_decap_8
Xfanout542 net542 net24 VPWR VGND sg13g2_buf_8
Xfanout564 _2007_ net564 VPWR VGND sg13g2_buf_8
Xfanout575 _0843_ net575 VPWR VGND sg13g2_buf_8
Xfanout553 _0751_ net553 VPWR VGND sg13g2_buf_8
XFILLER_47_927 VPWR VGND sg13g2_decap_8
XFILLER_19_607 VPWR VGND sg13g2_decap_8
Xfanout586 _0829_ net586 VPWR VGND sg13g2_buf_8
Xfanout597 _0727_ net597 VPWR VGND sg13g2_buf_8
XFILLER_46_437 VPWR VGND sg13g2_decap_8
XFILLER_27_662 VPWR VGND sg13g2_decap_8
XFILLER_42_643 VPWR VGND sg13g2_decap_8
XFILLER_15_857 VPWR VGND sg13g2_decap_8
XFILLER_6_533 VPWR VGND sg13g2_decap_8
XFILLER_10_573 VPWR VGND sg13g2_decap_8
XFILLER_29_1014 VPWR VGND sg13g2_decap_8
XFILLER_44_8 VPWR VGND sg13g2_fill_1
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_37_437 VPWR VGND sg13g2_fill_2
XFILLER_38_949 VPWR VGND sg13g2_decap_8
XFILLER_18_684 VPWR VGND sg13g2_decap_8
XFILLER_45_492 VPWR VGND sg13g2_decap_8
XFILLER_36_1018 VPWR VGND sg13g2_decap_8
X_3812_ _1265_ net607 _0921_ VPWR VGND sg13g2_nand2_1
XFILLER_33_676 VPWR VGND sg13g2_decap_8
XFILLER_21_849 VPWR VGND sg13g2_decap_8
X_3743_ _1002_ _1068_ _1210_ _1217_ VPWR VGND sg13g2_nor3_1
X_3674_ _0105_ _1167_ _1171_ net597 _1486_ VPWR VGND sg13g2_a22oi_1
X_2625_ _0222_ _0219_ _0220_ _0221_ VPWR VGND sg13g2_and3_1
X_2556_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] net622
+ net624 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] _1969_ net678 sg13g2_a221oi_1
X_2487_ _1902_ net629 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[4\] net631
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4226_ regFile_serial net29 VPWR VGND sg13g2_buf_8
XFILLER_28_404 VPWR VGND sg13g2_decap_4
XFILLER_29_916 VPWR VGND sg13g2_decap_8
X_4157_ net774 VGND VPWR _0135_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3108_ _0644_ net686 _1703_ VPWR VGND sg13g2_nand2_1
X_4088_ net772 VGND VPWR _0066_ sap_3_inst.controller.opcode\[7\] clknet_5_5__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_43_418 VPWR VGND sg13g2_decap_8
X_3039_ _0587_ VPWR _0054_ VGND net546 net667 sg13g2_o21ai_1
XFILLER_24_610 VPWR VGND sg13g2_decap_8
XFILLER_37_982 VPWR VGND sg13g2_decap_8
XFILLER_12_805 VPWR VGND sg13g2_decap_8
XFILLER_24_687 VPWR VGND sg13g2_decap_8
XFILLER_23_186 VPWR VGND sg13g2_fill_2
XFILLER_3_514 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_47_724 VPWR VGND sg13g2_decap_8
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
XFILLER_28_960 VPWR VGND sg13g2_decap_8
XFILLER_35_919 VPWR VGND sg13g2_decap_8
XFILLER_42_440 VPWR VGND sg13g2_decap_8
XFILLER_15_654 VPWR VGND sg13g2_decap_8
XFILLER_43_985 VPWR VGND sg13g2_decap_8
XFILLER_30_668 VPWR VGND sg13g2_decap_8
XFILLER_11_893 VPWR VGND sg13g2_decap_8
XFILLER_7_853 VPWR VGND sg13g2_decap_8
XFILLER_6_396 VPWR VGND sg13g2_fill_1
X_2410_ _1675_ net713 _1526_ _1831_ VPWR VGND sg13g2_a21o_1
X_3390_ _0787_ VPWR _0923_ VGND net560 _0850_ sg13g2_o21ai_1
X_2341_ _1760_ _1515_ _1748_ _1762_ VPWR VGND sg13g2_a21o_2
XFILLER_42_1000 VPWR VGND sg13g2_decap_8
X_2272_ _1693_ _1692_ net706 _1655_ net687 VPWR VGND sg13g2_a22oi_1
X_4011_ _0190_ _1497_ _1424_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_746 VPWR VGND sg13g2_decap_8
XFILLER_26_919 VPWR VGND sg13g2_decap_8
XFILLER_19_971 VPWR VGND sg13g2_decap_8
XFILLER_25_429 VPWR VGND sg13g2_decap_8
XFILLER_34_963 VPWR VGND sg13g2_decap_8
XFILLER_21_646 VPWR VGND sg13g2_decap_8
XFILLER_20_178 VPWR VGND sg13g2_fill_1
X_3726_ _0121_ _1114_ _1207_ net595 _1485_ VPWR VGND sg13g2_a22oi_1
X_3657_ VGND VPWR _1920_ net568 _1157_ _1156_ sg13g2_a21oi_1
X_2608_ net720 VPWR _0205_ VGND _1940_ _0204_ sg13g2_o21ai_1
X_3588_ _0087_ _1101_ _1103_ net589 _1474_ VPWR VGND sg13g2_a22oi_1
X_2539_ _1952_ net618 _1950_ VPWR VGND sg13g2_nand2_1
XFILLER_29_713 VPWR VGND sg13g2_decap_8
X_4209_ net783 VGND VPWR net766 u_ser.state\[0\] clknet_3_0__leaf_clk sg13g2_dfrbpq_2
XFILLER_44_738 VPWR VGND sg13g2_decap_8
XFILLER_40_900 VPWR VGND sg13g2_decap_8
XFILLER_12_602 VPWR VGND sg13g2_decap_8
XFILLER_19_1013 VPWR VGND sg13g2_decap_8
XFILLER_25_996 VPWR VGND sg13g2_decap_8
XFILLER_24_484 VPWR VGND sg13g2_decap_8
XFILLER_40_977 VPWR VGND sg13g2_decap_8
XFILLER_12_679 VPWR VGND sg13g2_decap_8
XFILLER_11_167 VPWR VGND sg13g2_fill_2
XFILLER_4_845 VPWR VGND sg13g2_decap_8
XFILLER_26_1017 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_521 VPWR VGND sg13g2_decap_8
XFILLER_19_212 VPWR VGND sg13g2_fill_2
XFILLER_47_598 VPWR VGND sg13g2_decap_8
XFILLER_35_716 VPWR VGND sg13g2_decap_8
XFILLER_16_963 VPWR VGND sg13g2_decap_8
XFILLER_31_911 VPWR VGND sg13g2_decap_8
XFILLER_43_782 VPWR VGND sg13g2_decap_8
X_2890_ net563 VPWR _0455_ VGND net750 sap_3_inst.alu.tmp\[4\] sg13g2_o21ai_1
XFILLER_30_465 VPWR VGND sg13g2_decap_8
XFILLER_31_988 VPWR VGND sg13g2_decap_8
XFILLER_8_87 VPWR VGND sg13g2_decap_8
XFILLER_7_650 VPWR VGND sg13g2_decap_8
XFILLER_11_690 VPWR VGND sg13g2_decap_8
X_3511_ VPWR _1039_ _1038_ VGND sg13g2_inv_1
XFILLER_6_182 VPWR VGND sg13g2_fill_1
X_3442_ _0973_ _0971_ _0972_ VPWR VGND sg13g2_nand2_1
X_3373_ _0907_ _0821_ _0808_ VPWR VGND sg13g2_nand2b_1
X_2324_ net702 VPWR _1745_ VGND _1500_ _1527_ sg13g2_o21ai_1
XFILLER_26_0 VPWR VGND sg13g2_fill_1
X_2255_ VGND VPWR net709 net685 _1676_ _1538_ sg13g2_a21oi_1
X_2186_ net707 _1605_ _1607_ VPWR VGND sg13g2_nor2_2
XFILLER_38_543 VPWR VGND sg13g2_decap_8
XFILLER_26_716 VPWR VGND sg13g2_decap_8
XFILLER_22_911 VPWR VGND sg13g2_decap_8
XFILLER_34_760 VPWR VGND sg13g2_decap_8
XFILLER_21_421 VPWR VGND sg13g2_fill_2
XFILLER_22_988 VPWR VGND sg13g2_decap_8
X_3709_ net595 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] _1196_ _0115_
+ VPWR VGND sg13g2_a21o_1
XFILLER_49_808 VPWR VGND sg13g2_decap_8
XFILLER_48_318 VPWR VGND sg13g2_decap_8
XFILLER_29_510 VPWR VGND sg13g2_decap_8
XFILLER_17_738 VPWR VGND sg13g2_decap_8
XFILLER_29_587 VPWR VGND sg13g2_decap_8
XFILLER_44_535 VPWR VGND sg13g2_decap_8
XFILLER_13_922 VPWR VGND sg13g2_decap_8
XFILLER_25_793 VPWR VGND sg13g2_decap_8
XFILLER_9_915 VPWR VGND sg13g2_decap_8
XFILLER_40_774 VPWR VGND sg13g2_decap_8
XFILLER_13_999 VPWR VGND sg13g2_decap_8
XFILLER_33_62 VPWR VGND sg13g2_fill_1
XFILLER_4_642 VPWR VGND sg13g2_decap_8
XFILLER_3_152 VPWR VGND sg13g2_fill_2
Xhold3 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[6\] VPWR VGND net50 sg13g2_dlygate4sd3_1
X_2040_ _1463_ sap_3_inst.alu.tmp\[1\] VPWR VGND sg13g2_inv_2
XFILLER_48_885 VPWR VGND sg13g2_decap_8
XFILLER_35_513 VPWR VGND sg13g2_decap_8
XFILLER_47_395 VPWR VGND sg13g2_decap_8
X_3991_ VGND VPWR net744 net663 _1409_ _1408_ sg13g2_a21oi_1
XFILLER_16_760 VPWR VGND sg13g2_decap_8
X_2942_ net745 sap_3_inst.alu.tmp\[6\] _0505_ VPWR VGND sg13g2_nor2_2
X_2873_ VPWR _0439_ _0438_ VGND sg13g2_inv_1
XFILLER_31_785 VPWR VGND sg13g2_decap_8
X_3425_ _0957_ _0919_ net552 VPWR VGND sg13g2_xnor2_1
X_3356_ _0890_ net656 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] net608
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2307_ _1612_ _1727_ _1728_ VPWR VGND sg13g2_nor2_1
X_3287_ _0787_ net560 _0808_ _0820_ _0823_ VPWR VGND sg13g2_and4_1
X_2238_ VGND VPWR _1659_ _1658_ _1612_ sg13g2_or2_1
XFILLER_39_852 VPWR VGND sg13g2_decap_8
XFILLER_26_513 VPWR VGND sg13g2_decap_8
X_2169_ _1522_ _1573_ _1520_ _1590_ VPWR VGND sg13g2_nand3_1
XFILLER_14_719 VPWR VGND sg13g2_decap_8
XFILLER_41_549 VPWR VGND sg13g2_decap_8
XFILLER_16_1005 VPWR VGND sg13g2_decap_8
XFILLER_22_785 VPWR VGND sg13g2_decap_8
XFILLER_6_918 VPWR VGND sg13g2_decap_8
XFILLER_10_958 VPWR VGND sg13g2_decap_8
XFILLER_49_605 VPWR VGND sg13g2_decap_8
XFILLER_1_667 VPWR VGND sg13g2_decap_8
XFILLER_45_800 VPWR VGND sg13g2_decap_8
XFILLER_17_535 VPWR VGND sg13g2_decap_8
XFILLER_29_395 VPWR VGND sg13g2_decap_4
XFILLER_45_877 VPWR VGND sg13g2_decap_8
XFILLER_44_376 VPWR VGND sg13g2_decap_4
XFILLER_25_590 VPWR VGND sg13g2_decap_8
XFILLER_40_571 VPWR VGND sg13g2_decap_8
XFILLER_9_712 VPWR VGND sg13g2_decap_8
XFILLER_12_240 VPWR VGND sg13g2_fill_1
XFILLER_13_796 VPWR VGND sg13g2_decap_8
XFILLER_8_233 VPWR VGND sg13g2_fill_2
XFILLER_9_789 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_4
X_3210_ _0746_ net643 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\] net652
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4190_ net797 VGND VPWR _0168_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[6\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
X_3141_ _1604_ _0675_ _0677_ VPWR VGND sg13g2_nor2_1
X_3072_ _0598_ VPWR _0608_ VGND _0313_ _0607_ sg13g2_o21ai_1
XFILLER_36_822 VPWR VGND sg13g2_decap_8
XFILLER_48_682 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk_div_out clk_div_out clknet_0_clk_div_out VPWR VGND sg13g2_buf_8
X_2023_ VPWR _1446_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_35_321 VPWR VGND sg13g2_fill_1
XFILLER_39_1027 VPWR VGND sg13g2_fill_2
XFILLER_36_899 VPWR VGND sg13g2_decap_8
X_3974_ _1397_ sap_3_inst.alu.act\[1\] net549 _0179_ VPWR VGND sg13g2_mux2_1
XFILLER_23_549 VPWR VGND sg13g2_decap_8
X_2925_ _0323_ VPWR _0489_ VGND net564 _0459_ sg13g2_o21ai_1
X_2856_ VGND VPWR _0422_ _0417_ _0415_ sg13g2_or2_1
XFILLER_31_582 VPWR VGND sg13g2_decap_8
X_2787_ sap_3_inst.alu.tmp\[1\] net758 _0355_ VPWR VGND sg13g2_xor2_1
Xfanout713 _1512_ net713 VPWR VGND sg13g2_buf_8
Xfanout724 _1505_ net724 VPWR VGND sg13g2_buf_8
Xfanout702 _1513_ net702 VPWR VGND sg13g2_buf_8
X_3408_ _0937_ _0938_ net610 _0940_ VPWR VGND _0939_ sg13g2_nand4_1
Xfanout735 net736 net735 VPWR VGND sg13g2_buf_8
Xfanout757 sap_3_inst.alu.acc\[1\] net757 VPWR VGND sg13g2_buf_8
Xfanout746 sap_3_inst.alu.acc\[6\] net746 VPWR VGND sg13g2_buf_8
Xfanout779 net781 net779 VPWR VGND sg13g2_buf_8
Xfanout768 sap_3_inst.reg_file.array_serializer_inst.word_index\[1\] net768 VPWR VGND
+ sg13g2_buf_8
X_3339_ _0874_ _0859_ _0871_ VPWR VGND sg13g2_xnor2_1
XFILLER_46_619 VPWR VGND sg13g2_decap_8
XFILLER_27_844 VPWR VGND sg13g2_decap_8
XFILLER_42_825 VPWR VGND sg13g2_decap_8
XFILLER_14_516 VPWR VGND sg13g2_decap_8
XFILLER_26_387 VPWR VGND sg13g2_decap_8
XFILLER_22_582 VPWR VGND sg13g2_decap_8
XFILLER_6_715 VPWR VGND sg13g2_decap_8
XFILLER_10_755 VPWR VGND sg13g2_decap_8
XFILLER_2_910 VPWR VGND sg13g2_decap_8
XFILLER_49_402 VPWR VGND sg13g2_decap_8
XFILLER_7_1014 VPWR VGND sg13g2_decap_8
XFILLER_2_987 VPWR VGND sg13g2_decap_8
XFILLER_1_464 VPWR VGND sg13g2_decap_8
XFILLER_49_479 VPWR VGND sg13g2_decap_8
XFILLER_18_866 VPWR VGND sg13g2_decap_8
XFILLER_45_674 VPWR VGND sg13g2_decap_8
XFILLER_32_357 VPWR VGND sg13g2_fill_2
XFILLER_33_858 VPWR VGND sg13g2_decap_8
X_2710_ _1593_ _1597_ _1590_ _0289_ VPWR VGND _1708_ sg13g2_nand4_1
XFILLER_13_593 VPWR VGND sg13g2_decap_8
XFILLER_9_586 VPWR VGND sg13g2_decap_8
X_3690_ net575 _0876_ _1185_ VPWR VGND sg13g2_nor2_2
X_2641_ _0236_ _0231_ _0235_ net639 _1460_ VPWR VGND sg13g2_a22oi_1
X_2572_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] net637
+ net622 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] _1983_ net624 sg13g2_a221oi_1
X_4173_ net774 VGND VPWR _0151_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\]
+ clknet_5_2__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3124_ _1439_ _1508_ net733 _0660_ VPWR VGND _0659_ sg13g2_nand4_1
X_3055_ _0594_ VPWR _0063_ VGND net691 _1920_ sg13g2_o21ai_1
XFILLER_36_696 VPWR VGND sg13g2_decap_8
XFILLER_24_869 VPWR VGND sg13g2_decap_8
XFILLER_11_508 VPWR VGND sg13g2_decap_8
X_3957_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] _1130_ net608 _0173_
+ VPWR VGND sg13g2_mux2_1
X_2908_ _0472_ net747 net671 VPWR VGND sg13g2_nand2_1
X_3888_ _1328_ _1313_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] _1308_
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2839_ _0396_ _0398_ _0332_ _0406_ VPWR VGND _0405_ sg13g2_nand4_1
XFILLER_47_906 VPWR VGND sg13g2_decap_8
Xfanout543 net544 net543 VPWR VGND sg13g2_buf_8
Xfanout554 net555 net554 VPWR VGND sg13g2_buf_8
Xfanout565 net567 net565 VPWR VGND sg13g2_buf_8
Xfanout598 net599 net598 VPWR VGND sg13g2_buf_8
XFILLER_46_416 VPWR VGND sg13g2_decap_8
Xfanout587 _0740_ net587 VPWR VGND sg13g2_buf_8
Xfanout576 _0843_ net576 VPWR VGND sg13g2_buf_8
XFILLER_27_641 VPWR VGND sg13g2_decap_8
XFILLER_42_622 VPWR VGND sg13g2_decap_8
XFILLER_15_836 VPWR VGND sg13g2_decap_8
XFILLER_42_699 VPWR VGND sg13g2_decap_8
XFILLER_10_552 VPWR VGND sg13g2_decap_8
XFILLER_6_512 VPWR VGND sg13g2_decap_8
XFILLER_6_589 VPWR VGND sg13g2_decap_8
XFILLER_2_784 VPWR VGND sg13g2_decap_8
XFILLER_38_928 VPWR VGND sg13g2_decap_8
XFILLER_18_663 VPWR VGND sg13g2_decap_8
XFILLER_46_983 VPWR VGND sg13g2_decap_8
XFILLER_45_471 VPWR VGND sg13g2_decap_8
XFILLER_32_132 VPWR VGND sg13g2_fill_2
XFILLER_33_655 VPWR VGND sg13g2_decap_8
XFILLER_21_828 VPWR VGND sg13g2_decap_8
X_3811_ _1264_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] net604 VPWR
+ VGND sg13g2_nand2_1
XFILLER_14_880 VPWR VGND sg13g2_decap_8
X_3742_ _1210_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] _1216_ _0128_
+ VPWR VGND sg13g2_a21o_1
X_3673_ VPWR VGND _1170_ _1070_ _1169_ _1117_ _1171_ _1168_ sg13g2_a221oi_1
X_2624_ _0221_ net626 sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] net628
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2555_ _1966_ _1967_ _1968_ VPWR VGND sg13g2_and2_1
X_2486_ _1901_ net619 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\] net633
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4225_ sap_3_outputReg_start_sync net28 VPWR VGND sg13g2_buf_1
X_4156_ net782 VGND VPWR _0134_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\]
+ clknet_5_26__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3107_ _1658_ net686 _1616_ _0643_ VPWR VGND sg13g2_a21o_1
XFILLER_28_449 VPWR VGND sg13g2_decap_8
X_4087_ net770 VGND VPWR _0065_ sap_3_inst.controller.opcode\[6\] clknet_5_5__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_37_961 VPWR VGND sg13g2_decap_8
X_3038_ _0587_ sap_3_inst.alu.tmp\[3\] net667 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_1_sap_3_inst.alu.clk clknet_1_1__leaf_sap_3_inst.alu.clk clknet_leaf_1_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_36_493 VPWR VGND sg13g2_decap_8
XFILLER_24_666 VPWR VGND sg13g2_decap_8
XFILLER_47_703 VPWR VGND sg13g2_decap_8
XFILLER_4_1006 VPWR VGND sg13g2_decap_8
XFILLER_14_110 VPWR VGND sg13g2_fill_1
XFILLER_15_633 VPWR VGND sg13g2_decap_8
XFILLER_43_964 VPWR VGND sg13g2_decap_8
XFILLER_42_496 VPWR VGND sg13g2_decap_8
XFILLER_30_647 VPWR VGND sg13g2_decap_8
XFILLER_7_832 VPWR VGND sg13g2_decap_8
XFILLER_11_872 VPWR VGND sg13g2_decap_8
X_2340_ VGND VPWR _1748_ _1761_ _1760_ _1515_ sg13g2_a21oi_2
X_2271_ VGND VPWR _1692_ _1691_ _1690_ sg13g2_or2_1
XFILLER_2_581 VPWR VGND sg13g2_decap_8
X_4010_ _1435_ _1288_ _1424_ VPWR VGND sg13g2_nor2_2
XFILLER_38_725 VPWR VGND sg13g2_decap_8
XFILLER_19_950 VPWR VGND sg13g2_decap_8
XFILLER_46_780 VPWR VGND sg13g2_decap_8
XFILLER_25_408 VPWR VGND sg13g2_decap_8
XFILLER_34_942 VPWR VGND sg13g2_decap_8
XFILLER_21_625 VPWR VGND sg13g2_decap_8
X_3725_ net595 _1068_ _1207_ VPWR VGND sg13g2_nor2_1
X_3656_ net13 net568 _1156_ VPWR VGND sg13g2_nor2_1
X_2607_ _0199_ _0200_ _0201_ _0203_ _0204_ VPWR VGND sg13g2_nor4_1
X_3587_ _1103_ _0957_ net577 _0946_ net584 VPWR VGND sg13g2_a22oi_1
X_2538_ _1951_ net732 _1928_ VPWR VGND sg13g2_nand2_2
X_2469_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] _1885_
+ net619 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] _1886_ net623 sg13g2_a221oi_1
X_4208_ net790 VGND VPWR _0185_ sap_3_inst.alu.act\[7\] clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_4139_ net773 VGND VPWR _0117_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\]
+ clknet_5_7__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_769 VPWR VGND sg13g2_decap_8
XFILLER_44_717 VPWR VGND sg13g2_decap_8
XFILLER_24_463 VPWR VGND sg13g2_decap_8
XFILLER_25_975 VPWR VGND sg13g2_decap_8
XFILLER_40_956 VPWR VGND sg13g2_decap_8
XFILLER_8_629 VPWR VGND sg13g2_decap_8
XFILLER_12_658 VPWR VGND sg13g2_decap_8
XFILLER_7_139 VPWR VGND sg13g2_fill_1
XFILLER_4_824 VPWR VGND sg13g2_decap_8
XFILLER_47_500 VPWR VGND sg13g2_decap_8
XFILLER_19_202 VPWR VGND sg13g2_fill_2
XFILLER_47_577 VPWR VGND sg13g2_decap_8
XFILLER_19_268 VPWR VGND sg13g2_fill_2
XFILLER_16_942 VPWR VGND sg13g2_decap_8
XFILLER_43_761 VPWR VGND sg13g2_decap_8
XFILLER_15_463 VPWR VGND sg13g2_fill_1
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_30_444 VPWR VGND sg13g2_decap_8
XFILLER_31_967 VPWR VGND sg13g2_decap_8
X_3510_ _1038_ net561 net586 VPWR VGND sg13g2_nand2_1
XFILLER_10_190 VPWR VGND sg13g2_fill_1
X_3441_ _0969_ VPWR _0972_ VGND _0931_ _0945_ sg13g2_o21ai_1
X_3372_ _0906_ _0808_ _0875_ VPWR VGND sg13g2_xnor2_1
X_2323_ sap_3_inst.controller.stage\[2\] _1527_ _1744_ VPWR VGND sg13g2_nor2_1
X_2254_ _1675_ net715 net710 VPWR VGND sg13g2_nand2_2
XFILLER_38_522 VPWR VGND sg13g2_decap_8
X_2185_ VGND VPWR _1606_ _1567_ _1517_ sg13g2_or2_1
XFILLER_25_205 VPWR VGND sg13g2_fill_2
XFILLER_38_599 VPWR VGND sg13g2_decap_8
XFILLER_33_271 VPWR VGND sg13g2_fill_1
XFILLER_22_967 VPWR VGND sg13g2_decap_8
XFILLER_21_499 VPWR VGND sg13g2_decap_8
XFILLER_4_109 VPWR VGND sg13g2_decap_4
X_3708_ net594 _0861_ _1040_ _1196_ VPWR VGND sg13g2_nor3_1
XFILLER_49_1018 VPWR VGND sg13g2_decap_8
X_3639_ net597 _0861_ _1142_ _1143_ VPWR VGND sg13g2_nor3_1
XFILLER_1_849 VPWR VGND sg13g2_decap_8
XFILLER_44_514 VPWR VGND sg13g2_decap_8
XFILLER_17_717 VPWR VGND sg13g2_decap_8
XFILLER_29_566 VPWR VGND sg13g2_decap_8
XFILLER_17_53 VPWR VGND sg13g2_fill_2
XFILLER_13_901 VPWR VGND sg13g2_decap_8
XFILLER_17_75 VPWR VGND sg13g2_fill_1
XFILLER_25_772 VPWR VGND sg13g2_decap_8
XFILLER_40_753 VPWR VGND sg13g2_decap_8
XFILLER_13_978 VPWR VGND sg13g2_decap_8
XFILLER_12_477 VPWR VGND sg13g2_fill_1
XFILLER_32_1022 VPWR VGND sg13g2_decap_8
XFILLER_4_621 VPWR VGND sg13g2_decap_8
XFILLER_4_698 VPWR VGND sg13g2_decap_8
Xclkbuf_5_8__f_sap_3_inst.alu.clk_regs clknet_4_4_0_sap_3_inst.alu.clk_regs clknet_5_8__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
Xhold4 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[3\] VPWR VGND net51 sg13g2_dlygate4sd3_1
XFILLER_48_864 VPWR VGND sg13g2_decap_8
XFILLER_47_374 VPWR VGND sg13g2_decap_8
X_3990_ _0542_ net663 _1408_ VPWR VGND sg13g2_nor2_1
XFILLER_35_569 VPWR VGND sg13g2_decap_8
X_2941_ _0503_ _1936_ _0504_ VPWR VGND _0502_ sg13g2_nand3b_1
X_2872_ VPWR VGND _0421_ net669 _0437_ net543 _0438_ _0425_ sg13g2_a221oi_1
XFILLER_31_764 VPWR VGND sg13g2_decap_8
XFILLER_8_993 VPWR VGND sg13g2_decap_8
X_3424_ net559 _0918_ net552 _0956_ VPWR VGND sg13g2_nor3_1
X_3355_ _0889_ net611 _0887_ _0888_ VPWR VGND sg13g2_and3_1
X_2306_ net714 VPWR _1727_ VGND net710 net705 sg13g2_o21ai_1
X_3286_ _0808_ _0820_ net561 _0822_ VPWR VGND sg13g2_nand3_1
X_2237_ _1658_ _1527_ net705 VPWR VGND sg13g2_nand2_2
XFILLER_39_831 VPWR VGND sg13g2_decap_8
X_2168_ net735 net737 _1521_ _1589_ VGND VPWR _1574_ sg13g2_nor4_2
X_2099_ net726 net727 _1520_ VPWR VGND sg13g2_nor2_2
XFILLER_26_569 VPWR VGND sg13g2_decap_8
XFILLER_41_528 VPWR VGND sg13g2_decap_8
XFILLER_10_937 VPWR VGND sg13g2_decap_8
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
XFILLER_22_764 VPWR VGND sg13g2_decap_8
XFILLER_21_285 VPWR VGND sg13g2_fill_1
XFILLER_0_112 VPWR VGND sg13g2_fill_1
Xclkbuf_5_15__f_sap_3_inst.alu.clk_regs clknet_4_7_0_sap_3_inst.alu.clk_regs clknet_5_15__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_0_145 VPWR VGND sg13g2_decap_8
XFILLER_0_123 VPWR VGND sg13g2_decap_4
XFILLER_1_646 VPWR VGND sg13g2_decap_8
XFILLER_45_856 VPWR VGND sg13g2_decap_8
XFILLER_17_514 VPWR VGND sg13g2_decap_8
XFILLER_44_388 VPWR VGND sg13g2_decap_8
XFILLER_32_539 VPWR VGND sg13g2_decap_8
XFILLER_40_550 VPWR VGND sg13g2_decap_8
XFILLER_13_775 VPWR VGND sg13g2_decap_8
XFILLER_9_768 VPWR VGND sg13g2_decap_8
XFILLER_5_985 VPWR VGND sg13g2_decap_8
XFILLER_5_34 VPWR VGND sg13g2_fill_2
XFILLER_4_495 VPWR VGND sg13g2_decap_8
X_3140_ _0676_ _1627_ _1703_ VPWR VGND sg13g2_nand2_1
XFILLER_48_661 VPWR VGND sg13g2_decap_8
X_3071_ _1835_ _0603_ _0605_ _0606_ _0607_ VPWR VGND sg13g2_nor4_1
XFILLER_36_801 VPWR VGND sg13g2_decap_8
X_2022_ VPWR _1445_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_36_878 VPWR VGND sg13g2_decap_8
XFILLER_39_1006 VPWR VGND sg13g2_decap_8
XFILLER_23_528 VPWR VGND sg13g2_decap_8
X_3973_ _0358_ net758 net664 _1397_ VPWR VGND sg13g2_mux2_1
X_2924_ _0486_ _0487_ _0488_ VPWR VGND sg13g2_nor2_1
XFILLER_31_561 VPWR VGND sg13g2_decap_8
X_2855_ VPWR VGND _1936_ _0420_ _0414_ net752 _0421_ net572 sg13g2_a221oi_1
XFILLER_8_790 VPWR VGND sg13g2_decap_8
X_2786_ _0354_ _1455_ _1463_ VPWR VGND sg13g2_nand2_1
Xfanout703 _1513_ net703 VPWR VGND sg13g2_buf_1
Xfanout714 _1501_ net714 VPWR VGND sg13g2_buf_8
X_3407_ _0939_ net649 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] net651
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] VPWR VGND sg13g2_a22oi_1
Xfanout758 sap_3_inst.alu.acc\[1\] net758 VPWR VGND sg13g2_buf_1
Xfanout725 sap_3_inst.controller.opcode\[7\] net725 VPWR VGND sg13g2_buf_8
Xfanout736 sap_3_inst.controller.opcode\[3\] net736 VPWR VGND sg13g2_buf_8
Xfanout747 net749 net747 VPWR VGND sg13g2_buf_8
X_3338_ _0873_ _0857_ _0872_ VPWR VGND sg13g2_nand2_2
Xfanout769 net80 net769 VPWR VGND sg13g2_buf_8
X_3269_ _1453_ _0713_ _0731_ _0805_ VPWR VGND sg13g2_nor3_1
XFILLER_27_823 VPWR VGND sg13g2_decap_8
XFILLER_42_804 VPWR VGND sg13g2_decap_8
XFILLER_22_561 VPWR VGND sg13g2_decap_8
XFILLER_10_734 VPWR VGND sg13g2_decap_8
XFILLER_2_966 VPWR VGND sg13g2_decap_8
XFILLER_1_443 VPWR VGND sg13g2_decap_8
XFILLER_49_458 VPWR VGND sg13g2_decap_8
XFILLER_18_845 VPWR VGND sg13g2_decap_8
XFILLER_45_653 VPWR VGND sg13g2_decap_8
XFILLER_32_314 VPWR VGND sg13g2_fill_1
XFILLER_33_837 VPWR VGND sg13g2_decap_8
XFILLER_41_892 VPWR VGND sg13g2_decap_8
XFILLER_13_572 VPWR VGND sg13g2_decap_8
XFILLER_9_565 VPWR VGND sg13g2_decap_8
X_2640_ _0235_ _0232_ _0233_ _0234_ VPWR VGND sg13g2_and3_1
X_2571_ _1979_ _1981_ _1982_ VPWR VGND sg13g2_and2_1
XFILLER_5_782 VPWR VGND sg13g2_decap_8
XFILLER_45_1010 VPWR VGND sg13g2_decap_8
X_4172_ net782 VGND VPWR _0150_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\]
+ clknet_5_7__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3123_ _1504_ _1675_ _0659_ VPWR VGND sg13g2_nor2_1
X_3054_ _0594_ net731 net691 VPWR VGND sg13g2_nand2_1
XFILLER_36_675 VPWR VGND sg13g2_decap_8
XFILLER_24_848 VPWR VGND sg13g2_decap_8
X_3956_ _1386_ VPWR _0172_ VGND _1445_ net608 sg13g2_o21ai_1
X_2907_ net671 net751 _0444_ _0471_ VPWR VGND sg13g2_a21o_1
X_3887_ _1327_ VPWR _0162_ VGND _1325_ _1326_ sg13g2_o21ai_1
X_2838_ VPWR VGND _0322_ _0404_ _0391_ net758 _0405_ net573 sg13g2_a221oi_1
X_2769_ _1949_ _0198_ _0338_ VPWR VGND sg13g2_nor2_1
Xfanout555 _0319_ net555 VPWR VGND sg13g2_buf_8
Xfanout544 _0331_ net544 VPWR VGND sg13g2_buf_8
Xfanout566 net567 net566 VPWR VGND sg13g2_buf_1
Xfanout588 _0740_ net588 VPWR VGND sg13g2_buf_8
Xfanout599 _0724_ net599 VPWR VGND sg13g2_buf_8
Xfanout577 net582 net577 VPWR VGND sg13g2_buf_8
XFILLER_27_620 VPWR VGND sg13g2_decap_8
XFILLER_42_601 VPWR VGND sg13g2_decap_8
XFILLER_15_815 VPWR VGND sg13g2_decap_8
XFILLER_27_697 VPWR VGND sg13g2_decap_8
XFILLER_26_174 VPWR VGND sg13g2_fill_1
XFILLER_42_678 VPWR VGND sg13g2_decap_8
XFILLER_41_144 VPWR VGND sg13g2_fill_2
XFILLER_14_369 VPWR VGND sg13g2_fill_2
XFILLER_30_829 VPWR VGND sg13g2_decap_8
XFILLER_23_892 VPWR VGND sg13g2_decap_8
XFILLER_10_531 VPWR VGND sg13g2_decap_8
XFILLER_6_568 VPWR VGND sg13g2_decap_8
XFILLER_2_763 VPWR VGND sg13g2_decap_8
XFILLER_49_244 VPWR VGND sg13g2_fill_1
XFILLER_38_907 VPWR VGND sg13g2_decap_8
XFILLER_46_962 VPWR VGND sg13g2_decap_8
XFILLER_18_642 VPWR VGND sg13g2_decap_8
XFILLER_45_450 VPWR VGND sg13g2_decap_8
XFILLER_33_634 VPWR VGND sg13g2_decap_8
XFILLER_21_807 VPWR VGND sg13g2_decap_8
X_3810_ _0149_ _0901_ _1263_ net603 _1446_ VPWR VGND sg13g2_a22oi_1
XFILLER_32_155 VPWR VGND sg13g2_fill_1
X_3741_ _1133_ _1134_ net556 _1216_ VPWR VGND sg13g2_nor3_1
XFILLER_32_166 VPWR VGND sg13g2_fill_2
XFILLER_9_384 VPWR VGND sg13g2_fill_2
X_3672_ VGND VPWR _1170_ net569 net15 sg13g2_or2_1
X_2623_ _0220_ net630 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] net636
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2554_ _1967_ net634 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] net636
+ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
X_2485_ VGND VPWR net676 _1899_ _0031_ _1900_ sg13g2_a21oi_1
X_4224_ sap_3_outputReg_serial net27 VPWR VGND sg13g2_buf_1
X_4155_ net774 VGND VPWR _0133_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\]
+ clknet_5_1__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3106_ _1651_ net686 _1607_ _0642_ VPWR VGND sg13g2_a21o_1
X_4086_ net771 VGND VPWR _0064_ sap_3_inst.controller.opcode\[5\] clknet_5_5__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_37_940 VPWR VGND sg13g2_decap_8
X_3037_ net19 sap_3_inst.alu.tmp\[2\] net667 _0053_ VPWR VGND sg13g2_mux2_1
XFILLER_24_645 VPWR VGND sg13g2_decap_8
X_3939_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\] _1373_
+ _1314_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] _1374_ _1312_ sg13g2_a221oi_1
XFILLER_20_884 VPWR VGND sg13g2_decap_8
XFILLER_3_549 VPWR VGND sg13g2_decap_8
XFILLER_11_88 VPWR VGND sg13g2_fill_1
XFILLER_47_759 VPWR VGND sg13g2_decap_8
XFILLER_15_612 VPWR VGND sg13g2_decap_8
XFILLER_28_995 VPWR VGND sg13g2_decap_8
XFILLER_36_41 VPWR VGND sg13g2_fill_2
XFILLER_43_943 VPWR VGND sg13g2_decap_8
XFILLER_27_494 VPWR VGND sg13g2_decap_8
XFILLER_36_85 VPWR VGND sg13g2_fill_2
XFILLER_42_475 VPWR VGND sg13g2_decap_8
XFILLER_15_689 VPWR VGND sg13g2_decap_8
XFILLER_30_626 VPWR VGND sg13g2_decap_8
XFILLER_11_851 VPWR VGND sg13g2_decap_8
XFILLER_7_811 VPWR VGND sg13g2_decap_8
XFILLER_7_888 VPWR VGND sg13g2_decap_8
XFILLER_2_560 VPWR VGND sg13g2_decap_8
X_2270_ _1536_ _1625_ _1691_ VPWR VGND sg13g2_nor2_1
XFILLER_38_704 VPWR VGND sg13g2_decap_8
XFILLER_34_921 VPWR VGND sg13g2_decap_8
XFILLER_21_604 VPWR VGND sg13g2_decap_8
XFILLER_34_998 VPWR VGND sg13g2_decap_8
X_3724_ _1206_ VPWR _0120_ VGND _1477_ net643 sg13g2_o21ai_1
X_3655_ _0946_ VPWR _1155_ VGND net652 _0947_ sg13g2_o21ai_1
X_2606_ _1952_ _0202_ _0203_ VPWR VGND sg13g2_nor2b_1
X_3586_ _1102_ net577 _0957_ VPWR VGND sg13g2_nand2_1
XFILLER_0_519 VPWR VGND sg13g2_decap_8
X_2537_ net732 _1928_ _1950_ VPWR VGND sg13g2_and2_1
X_2468_ _1883_ _1884_ _1882_ _1885_ VPWR VGND sg13g2_nand3_1
X_4207_ net790 VGND VPWR _0184_ sap_3_inst.alu.act\[6\] clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_2399_ _1819_ VPWR _1820_ VGND _1551_ _1814_ sg13g2_o21ai_1
X_4138_ net773 VGND VPWR _0116_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_748 VPWR VGND sg13g2_decap_8
X_4069_ net789 VGND VPWR _0047_ sap_3_inst.out\[5\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_24_442 VPWR VGND sg13g2_decap_8
XFILLER_25_954 VPWR VGND sg13g2_decap_8
XFILLER_36_291 VPWR VGND sg13g2_fill_1
XFILLER_40_935 VPWR VGND sg13g2_decap_8
XFILLER_12_637 VPWR VGND sg13g2_decap_8
XFILLER_8_608 VPWR VGND sg13g2_decap_8
XFILLER_11_169 VPWR VGND sg13g2_fill_1
XFILLER_20_681 VPWR VGND sg13g2_decap_8
XFILLER_4_803 VPWR VGND sg13g2_decap_8
XFILLER_47_556 VPWR VGND sg13g2_decap_8
XFILLER_16_921 VPWR VGND sg13g2_decap_8
XFILLER_28_792 VPWR VGND sg13g2_decap_8
XFILLER_43_740 VPWR VGND sg13g2_decap_8
XFILLER_42_250 VPWR VGND sg13g2_fill_2
XFILLER_16_998 VPWR VGND sg13g2_decap_8
XFILLER_31_946 VPWR VGND sg13g2_decap_8
XFILLER_8_23 VPWR VGND sg13g2_fill_2
XFILLER_7_685 VPWR VGND sg13g2_decap_8
X_3440_ _0930_ net552 _0882_ _0971_ VPWR VGND _0970_ sg13g2_nand4_1
X_3371_ _0905_ _0904_ net614 net562 sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[2\]
+ VPWR VGND sg13g2_a22oi_1
X_2322_ net709 net684 net740 _1743_ VPWR VGND sg13g2_nand3_1
X_2253_ net715 _1556_ _1674_ VPWR VGND sg13g2_and2_1
XFILLER_38_501 VPWR VGND sg13g2_decap_8
X_2184_ _1517_ _1567_ _1605_ VPWR VGND sg13g2_nor2_2
XFILLER_38_578 VPWR VGND sg13g2_decap_8
XFILLER_34_795 VPWR VGND sg13g2_decap_8
XFILLER_22_946 VPWR VGND sg13g2_decap_8
XFILLER_21_478 VPWR VGND sg13g2_decap_8
XFILLER_30_990 VPWR VGND sg13g2_decap_8
X_3707_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\] _1195_ _1182_ _0114_
+ VPWR VGND sg13g2_mux2_1
X_3638_ VPWR VGND _1141_ _1138_ _1140_ _0727_ _1142_ _1039_ sg13g2_a221oi_1
X_3569_ VPWR VGND _1087_ net589 _0884_ net577 _1088_ _0874_ sg13g2_a221oi_1
XFILLER_1_828 VPWR VGND sg13g2_decap_8
XFILLER_0_338 VPWR VGND sg13g2_fill_1
XFILLER_29_545 VPWR VGND sg13g2_decap_8
XFILLER_25_751 VPWR VGND sg13g2_decap_8
XFILLER_40_732 VPWR VGND sg13g2_decap_8
XFILLER_13_957 VPWR VGND sg13g2_decap_8
XFILLER_32_1001 VPWR VGND sg13g2_decap_8
XFILLER_4_600 VPWR VGND sg13g2_decap_8
XFILLER_4_677 VPWR VGND sg13g2_decap_8
XFILLER_3_154 VPWR VGND sg13g2_fill_1
XFILLER_3_143 VPWR VGND sg13g2_decap_4
XFILLER_0_883 VPWR VGND sg13g2_decap_8
XFILLER_48_843 VPWR VGND sg13g2_decap_8
Xhold5 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[7\] VPWR VGND net52 sg13g2_dlygate4sd3_1
XFILLER_47_353 VPWR VGND sg13g2_decap_8
XFILLER_35_548 VPWR VGND sg13g2_decap_8
XFILLER_16_795 VPWR VGND sg13g2_decap_8
X_2940_ _0500_ _0501_ _0472_ _0503_ VPWR VGND sg13g2_nand3_1
X_2871_ net543 _0434_ _0435_ _0436_ _0437_ VPWR VGND sg13g2_nor4_1
XFILLER_31_743 VPWR VGND sg13g2_decap_8
XFILLER_8_972 VPWR VGND sg13g2_decap_8
X_3423_ _0918_ net552 _0955_ VPWR VGND sg13g2_nor2_1
X_3354_ _0888_ net645 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] net653
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_31_0 VPWR VGND sg13g2_fill_1
X_2305_ VPWR VGND _1594_ _1725_ _1646_ _1608_ _1726_ _1637_ sg13g2_a221oi_1
X_3285_ _0821_ net561 _0820_ VPWR VGND sg13g2_nand2_1
XFILLER_39_810 VPWR VGND sg13g2_decap_8
X_2236_ net722 _1528_ _1595_ _1625_ _1657_ VPWR VGND sg13g2_nor4_1
XFILLER_38_320 VPWR VGND sg13g2_fill_1
XFILLER_39_887 VPWR VGND sg13g2_decap_8
X_2167_ _1506_ _1561_ _1436_ _1588_ VPWR VGND sg13g2_nand3_1
XFILLER_41_507 VPWR VGND sg13g2_decap_8
X_2098_ VGND VPWR _1519_ net729 net732 sg13g2_or2_1
XFILLER_26_548 VPWR VGND sg13g2_decap_8
XFILLER_22_743 VPWR VGND sg13g2_decap_8
XFILLER_34_592 VPWR VGND sg13g2_decap_8
XFILLER_10_916 VPWR VGND sg13g2_decap_8
Xclkbuf_regs_0_clk_div_two sap_3_inst.alu.clk sap_3_inst.alu.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_1_625 VPWR VGND sg13g2_decap_8
XFILLER_45_835 VPWR VGND sg13g2_decap_8
XFILLER_32_518 VPWR VGND sg13g2_decap_8
XFILLER_13_754 VPWR VGND sg13g2_decap_8
XFILLER_8_235 VPWR VGND sg13g2_fill_1
XFILLER_9_747 VPWR VGND sg13g2_decap_8
XFILLER_5_964 VPWR VGND sg13g2_decap_8
XFILLER_4_474 VPWR VGND sg13g2_decap_8
XFILLER_0_680 VPWR VGND sg13g2_decap_8
X_3070_ _0599_ _0601_ _1730_ _0606_ VPWR VGND _0602_ sg13g2_nand4_1
XFILLER_48_640 VPWR VGND sg13g2_decap_8
X_2021_ VPWR _1444_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[2\] VGND
+ sg13g2_inv_1
XFILLER_47_150 VPWR VGND sg13g2_fill_1
XFILLER_36_857 VPWR VGND sg13g2_decap_8
XFILLER_23_507 VPWR VGND sg13g2_decap_8
X_3972_ VGND VPWR _1462_ net549 _0178_ _1396_ sg13g2_a21oi_1
XFILLER_16_592 VPWR VGND sg13g2_decap_8
X_2923_ VGND VPWR _0457_ _0485_ _0487_ _0479_ sg13g2_a21oi_1
XFILLER_31_540 VPWR VGND sg13g2_decap_8
X_2854_ _0419_ VPWR _0420_ VGND _0417_ _0418_ sg13g2_o21ai_1
X_2785_ _0353_ net757 sap_3_inst.alu.tmp\[1\] VPWR VGND sg13g2_nand2_1
Xfanout704 net705 net704 VPWR VGND sg13g2_buf_8
Xfanout715 _1501_ net715 VPWR VGND sg13g2_buf_1
X_3406_ _0938_ net643 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] net646
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] VPWR VGND sg13g2_a22oi_1
Xfanout737 net738 net737 VPWR VGND sg13g2_buf_8
Xfanout748 net749 net748 VPWR VGND sg13g2_buf_1
Xfanout726 sap_3_inst.controller.opcode\[7\] net726 VPWR VGND sg13g2_buf_2
X_3337_ _0872_ _0871_ VPWR VGND sg13g2_inv_2
Xfanout759 net760 net759 VPWR VGND sg13g2_buf_8
X_3268_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[2\] net640 _0804_ VPWR
+ VGND sg13g2_and2_1
XFILLER_27_802 VPWR VGND sg13g2_decap_8
X_2219_ _1640_ _1533_ net705 VPWR VGND sg13g2_nand2_1
X_3199_ _0735_ net644 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\] net646
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_684 VPWR VGND sg13g2_decap_8
XFILLER_27_879 VPWR VGND sg13g2_decap_8
XFILLER_41_326 VPWR VGND sg13g2_fill_1
XFILLER_22_540 VPWR VGND sg13g2_decap_8
XFILLER_10_713 VPWR VGND sg13g2_decap_8
XFILLER_2_945 VPWR VGND sg13g2_decap_8
XFILLER_49_437 VPWR VGND sg13g2_decap_8
XFILLER_1_499 VPWR VGND sg13g2_decap_8
XFILLER_18_824 VPWR VGND sg13g2_decap_8
XFILLER_45_632 VPWR VGND sg13g2_decap_8
XFILLER_17_323 VPWR VGND sg13g2_fill_1
XFILLER_33_816 VPWR VGND sg13g2_decap_8
XFILLER_41_871 VPWR VGND sg13g2_decap_8
XFILLER_13_551 VPWR VGND sg13g2_decap_8
XFILLER_32_359 VPWR VGND sg13g2_fill_1
XFILLER_9_544 VPWR VGND sg13g2_decap_8
X_2570_ _1981_ net636 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[2\] net679
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_761 VPWR VGND sg13g2_decap_8
X_4171_ net771 VGND VPWR _0149_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[2\]
+ clknet_5_0__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3122_ _0652_ net702 _0655_ _0658_ VPWR VGND sg13g2_a21o_2
X_3053_ _0593_ VPWR _0062_ VGND net691 net546 sg13g2_o21ai_1
XFILLER_36_654 VPWR VGND sg13g2_decap_8
XFILLER_24_827 VPWR VGND sg13g2_decap_8
X_3955_ _1386_ _1385_ _1201_ VPWR VGND sg13g2_nand2b_1
X_4032__10 VPWR net44 clknet_leaf_1_sap_3_inst.alu.clk VGND sg13g2_inv_1
X_2906_ net554 net751 _0470_ _0038_ VPWR VGND sg13g2_a21o_1
XFILLER_32_882 VPWR VGND sg13g2_decap_8
X_3886_ _1327_ net48 net764 VPWR VGND sg13g2_nand2_1
X_2837_ _0404_ _1936_ _0402_ _0403_ VPWR VGND sg13g2_and3_1
X_2768_ net720 _1950_ _0337_ VPWR VGND sg13g2_and2_1
XFILLER_2_208 VPWR VGND sg13g2_fill_1
X_2699_ net566 _1963_ net12 VPWR VGND sg13g2_nor2b_2
Xfanout556 _1210_ net556 VPWR VGND sg13g2_buf_8
Xfanout545 net545 net19 VPWR VGND sg13g2_buf_8
Xfanout578 net579 net578 VPWR VGND sg13g2_buf_8
Xfanout567 _1673_ net567 VPWR VGND sg13g2_buf_8
Xfanout589 net591 net589 VPWR VGND sg13g2_buf_8
XFILLER_39_481 VPWR VGND sg13g2_decap_8
XFILLER_27_676 VPWR VGND sg13g2_decap_8
XFILLER_41_101 VPWR VGND sg13g2_fill_1
XFILLER_14_337 VPWR VGND sg13g2_fill_1
XFILLER_42_657 VPWR VGND sg13g2_decap_8
XFILLER_14_348 VPWR VGND sg13g2_fill_1
XFILLER_30_808 VPWR VGND sg13g2_decap_8
XFILLER_10_510 VPWR VGND sg13g2_decap_8
XFILLER_23_871 VPWR VGND sg13g2_decap_8
XFILLER_10_587 VPWR VGND sg13g2_decap_8
XFILLER_6_547 VPWR VGND sg13g2_decap_8
XFILLER_2_742 VPWR VGND sg13g2_decap_8
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_25 VPWR VGND sg13g2_fill_1
XFILLER_46_941 VPWR VGND sg13g2_decap_8
XFILLER_18_621 VPWR VGND sg13g2_decap_8
XFILLER_33_613 VPWR VGND sg13g2_decap_8
XFILLER_18_698 VPWR VGND sg13g2_decap_8
XFILLER_32_134 VPWR VGND sg13g2_fill_1
X_3740_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] _1188_ _1211_ _0127_
+ VPWR VGND sg13g2_mux2_1
X_3671_ _1169_ net547 net569 VPWR VGND sg13g2_nand2_1
X_2622_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] net622
+ net634 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\] _0219_ net679 sg13g2_a221oi_1
X_2553_ _1966_ net632 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] _1794_
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2484_ sap_3_inst.alu.flags\[5\] net676 _1900_ VPWR VGND sg13g2_nor2_1
X_4223_ mem_mar_we net26 VPWR VGND sg13g2_buf_1
X_4154_ net770 VGND VPWR _0132_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[1\]
+ clknet_5_4__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3105_ _0641_ net680 _0640_ VPWR VGND sg13g2_nand2b_1
X_4085_ net770 VGND VPWR _0063_ sap_3_inst.controller.opcode\[4\] clknet_5_0__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3036_ VGND VPWR _1463_ net668 _0052_ _0586_ sg13g2_a21oi_1
XFILLER_37_996 VPWR VGND sg13g2_decap_8
XFILLER_24_624 VPWR VGND sg13g2_decap_8
XFILLER_12_819 VPWR VGND sg13g2_decap_8
X_3938_ _1370_ _1371_ _1368_ _1373_ VPWR VGND _1372_ sg13g2_nand4_1
X_3869_ sap_3_inst.reg_file.array_serializer_inst.word_index\[2\] sap_3_inst.reg_file.array_serializer_inst.word_index\[3\]
+ _1309_ _1310_ VPWR VGND sg13g2_a21o_2
XFILLER_20_863 VPWR VGND sg13g2_decap_8
XFILLER_3_528 VPWR VGND sg13g2_decap_8
XFILLER_47_738 VPWR VGND sg13g2_decap_8
XFILLER_28_974 VPWR VGND sg13g2_decap_8
XFILLER_43_922 VPWR VGND sg13g2_decap_8
XFILLER_27_473 VPWR VGND sg13g2_decap_8
XFILLER_42_454 VPWR VGND sg13g2_decap_8
XFILLER_15_668 VPWR VGND sg13g2_decap_8
XFILLER_30_605 VPWR VGND sg13g2_decap_8
XFILLER_43_999 VPWR VGND sg13g2_decap_8
XFILLER_35_1010 VPWR VGND sg13g2_decap_8
XFILLER_11_830 VPWR VGND sg13g2_decap_8
XFILLER_7_867 VPWR VGND sg13g2_decap_8
XFILLER_42_1014 VPWR VGND sg13g2_decap_8
XFILLER_19_985 VPWR VGND sg13g2_decap_8
XFILLER_34_900 VPWR VGND sg13g2_decap_8
XFILLER_18_473 VPWR VGND sg13g2_fill_2
XFILLER_34_977 VPWR VGND sg13g2_decap_8
X_3723_ net643 _1112_ _1206_ VPWR VGND _1133_ sg13g2_nand3b_1
X_3654_ _1149_ VPWR _0102_ VGND _1153_ _1154_ sg13g2_o21ai_1
X_2605_ _1943_ _1944_ _0202_ VPWR VGND sg13g2_nor2b_2
X_3585_ net589 _1100_ _1101_ VPWR VGND sg13g2_nor2_1
X_2536_ _1948_ VPWR _1949_ VGND _1612_ _1627_ sg13g2_o21ai_1
X_2467_ _1884_ net631 sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[5\] net677
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4206_ net790 VGND VPWR _0183_ sap_3_inst.alu.act\[5\] clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_2398_ net689 _1816_ _1817_ _1818_ _1819_ VPWR VGND sg13g2_or4_1
XFILLER_29_727 VPWR VGND sg13g2_decap_8
X_4137_ net796 VGND VPWR _0115_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[0\]
+ clknet_5_30__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4068_ net789 VGND VPWR _0046_ sap_3_inst.out\[4\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3019_ sap_3_inst.alu.tmp\[6\] net746 _0539_ _0572_ VPWR VGND sg13g2_a21o_1
XFILLER_24_421 VPWR VGND sg13g2_decap_8
XFILLER_25_933 VPWR VGND sg13g2_decap_8
XFILLER_37_793 VPWR VGND sg13g2_decap_8
XFILLER_19_1027 VPWR VGND sg13g2_fill_2
XFILLER_40_914 VPWR VGND sg13g2_decap_8
XFILLER_12_616 VPWR VGND sg13g2_decap_8
XFILLER_24_498 VPWR VGND sg13g2_decap_8
XFILLER_20_660 VPWR VGND sg13g2_decap_8
XFILLER_4_859 VPWR VGND sg13g2_decap_8
XFILLER_47_535 VPWR VGND sg13g2_decap_8
XFILLER_16_900 VPWR VGND sg13g2_decap_8
XFILLER_28_771 VPWR VGND sg13g2_decap_8
XFILLER_16_977 VPWR VGND sg13g2_decap_8
XFILLER_43_796 VPWR VGND sg13g2_decap_8
XFILLER_30_413 VPWR VGND sg13g2_fill_1
XFILLER_31_925 VPWR VGND sg13g2_decap_8
XFILLER_8_46 VPWR VGND sg13g2_fill_1
XFILLER_30_479 VPWR VGND sg13g2_decap_8
XFILLER_8_79 VPWR VGND sg13g2_fill_2
XFILLER_7_664 VPWR VGND sg13g2_decap_8
X_3370_ _0610_ _0902_ _0903_ _0904_ VPWR VGND sg13g2_nor3_1
XFILLER_3_892 VPWR VGND sg13g2_decap_8
X_2321_ VGND VPWR net739 _1720_ _1742_ net712 sg13g2_a21oi_1
X_2252_ _1673_ _1537_ _1672_ net715 _1499_ VPWR VGND sg13g2_a22oi_1
X_2183_ _1519_ _1567_ _1595_ _1604_ VPWR VGND sg13g2_or3_1
XFILLER_38_557 VPWR VGND sg13g2_decap_8
XFILLER_19_782 VPWR VGND sg13g2_decap_8
Xclkbuf_5_23__f_sap_3_inst.alu.clk_regs clknet_4_11_0_sap_3_inst.alu.clk_regs clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_22_925 VPWR VGND sg13g2_decap_8
XFILLER_34_774 VPWR VGND sg13g2_decap_8
X_3706_ _1024_ net578 _1194_ _1195_ VPWR VGND sg13g2_a21o_2
X_3637_ VGND VPWR _1141_ net569 net9 sg13g2_or2_1
XFILLER_1_807 VPWR VGND sg13g2_decap_8
X_3568_ _1085_ _1086_ _1087_ VPWR VGND sg13g2_nor2_1
X_2519_ _1932_ _1559_ _1627_ VPWR VGND sg13g2_nand2_1
X_3499_ _1028_ net553 _0825_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_524 VPWR VGND sg13g2_decap_8
XFILLER_44_549 VPWR VGND sg13g2_decap_8
XFILLER_25_730 VPWR VGND sg13g2_decap_8
XFILLER_37_590 VPWR VGND sg13g2_decap_8
XFILLER_40_711 VPWR VGND sg13g2_decap_8
XFILLER_13_936 VPWR VGND sg13g2_decap_8
XFILLER_40_788 VPWR VGND sg13g2_decap_8
XFILLER_9_929 VPWR VGND sg13g2_decap_8
XFILLER_12_468 VPWR VGND sg13g2_fill_1
XFILLER_4_656 VPWR VGND sg13g2_decap_8
XFILLER_3_122 VPWR VGND sg13g2_decap_8
XFILLER_0_862 VPWR VGND sg13g2_decap_8
XFILLER_48_822 VPWR VGND sg13g2_decap_8
Xhold6 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[1\] VPWR VGND net53 sg13g2_dlygate4sd3_1
XFILLER_47_332 VPWR VGND sg13g2_decap_8
XFILLER_48_899 VPWR VGND sg13g2_decap_8
XFILLER_35_527 VPWR VGND sg13g2_decap_8
XFILLER_16_774 VPWR VGND sg13g2_decap_8
XFILLER_43_593 VPWR VGND sg13g2_decap_8
X_2870_ net753 _0327_ _0436_ VPWR VGND sg13g2_nor2_1
XFILLER_31_722 VPWR VGND sg13g2_decap_8
XFILLER_12_980 VPWR VGND sg13g2_decap_8
XFILLER_30_265 VPWR VGND sg13g2_fill_1
XFILLER_31_799 VPWR VGND sg13g2_decap_8
XFILLER_8_951 VPWR VGND sg13g2_decap_8
X_3422_ VPWR VGND _0950_ _0953_ _0949_ net584 _0954_ _0948_ sg13g2_a221oi_1
X_3353_ _0887_ net648 sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] net650
+ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2304_ _1627_ _1662_ _1725_ VPWR VGND sg13g2_nor2_1
X_3284_ _0814_ _0819_ _0820_ VPWR VGND sg13g2_and2_1
X_2235_ net722 _1528_ _1595_ _1656_ VPWR VGND sg13g2_nor3_1
X_2166_ net738 _1507_ _1562_ _1587_ VPWR VGND sg13g2_nor3_2
XFILLER_39_866 VPWR VGND sg13g2_decap_8
XFILLER_26_527 VPWR VGND sg13g2_decap_8
X_2097_ sap_3_inst.controller.opcode\[4\] net730 _1518_ VPWR VGND sg13g2_nor2_2
XFILLER_34_571 VPWR VGND sg13g2_decap_8
XFILLER_22_722 VPWR VGND sg13g2_decap_8
XFILLER_16_1019 VPWR VGND sg13g2_decap_8
X_2999_ _0560_ sap_3_inst.out\[0\] net673 VPWR VGND sg13g2_nand2_1
XFILLER_22_799 VPWR VGND sg13g2_decap_8
XFILLER_0_103 VPWR VGND sg13g2_decap_8
XFILLER_1_604 VPWR VGND sg13g2_decap_8
XFILLER_49_619 VPWR VGND sg13g2_decap_8
XFILLER_45_814 VPWR VGND sg13g2_decap_8
XFILLER_44_313 VPWR VGND sg13g2_decap_4
XFILLER_17_549 VPWR VGND sg13g2_decap_8
XFILLER_13_733 VPWR VGND sg13g2_decap_8
XFILLER_9_726 VPWR VGND sg13g2_decap_8
XFILLER_40_585 VPWR VGND sg13g2_decap_8
XFILLER_5_943 VPWR VGND sg13g2_decap_8
XFILLER_5_36 VPWR VGND sg13g2_fill_1
XFILLER_5_69 VPWR VGND sg13g2_fill_1
XFILLER_4_453 VPWR VGND sg13g2_decap_8
X_2020_ VPWR _1443_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] VGND
+ sg13g2_inv_1
XFILLER_48_696 VPWR VGND sg13g2_decap_8
XFILLER_36_836 VPWR VGND sg13g2_decap_8
X_3971_ net549 _1395_ _1396_ VPWR VGND sg13g2_nor2_1
X_2922_ _0486_ _0457_ _0479_ _0485_ VPWR VGND sg13g2_and3_1
XFILLER_16_571 VPWR VGND sg13g2_decap_8
X_2853_ _0419_ _0340_ _0415_ net573 net755 VPWR VGND sg13g2_a22oi_1
XFILLER_31_596 VPWR VGND sg13g2_decap_8
X_2784_ VGND VPWR _1456_ net555 _0034_ _0352_ sg13g2_a21oi_1
X_3405_ _0937_ net655 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\] net606
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] VPWR VGND sg13g2_a22oi_1
Xfanout705 _1624_ net705 VPWR VGND sg13g2_buf_8
Xfanout716 sap_3_inst.controller.stage\[3\] net716 VPWR VGND sg13g2_buf_8
Xfanout727 sap_3_inst.controller.opcode\[6\] net727 VPWR VGND sg13g2_buf_8
Xfanout749 sap_3_inst.alu.acc\[5\] net749 VPWR VGND sg13g2_buf_8
Xfanout738 sap_3_inst.controller.opcode\[2\] net738 VPWR VGND sg13g2_buf_8
X_3336_ _0870_ VPWR _0871_ VGND sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[1\]
+ net610 sg13g2_o21ai_1
XFILLER_22_1023 VPWR VGND sg13g2_decap_4
X_3267_ _1454_ _0673_ _0713_ _0803_ VPWR VGND sg13g2_nor3_1
XFILLER_39_663 VPWR VGND sg13g2_decap_8
X_2218_ _1533_ net705 _1639_ VPWR VGND sg13g2_and2_1
X_3198_ _0734_ _0710_ _0719_ VPWR VGND sg13g2_nand2_2
X_2149_ _1570_ net699 _1568_ VPWR VGND sg13g2_nand2_1
XFILLER_27_858 VPWR VGND sg13g2_decap_8
XFILLER_42_839 VPWR VGND sg13g2_decap_8
XFILLER_35_891 VPWR VGND sg13g2_decap_8
XFILLER_22_596 VPWR VGND sg13g2_decap_8
XFILLER_10_769 VPWR VGND sg13g2_decap_8
XFILLER_6_729 VPWR VGND sg13g2_decap_8
XFILLER_2_924 VPWR VGND sg13g2_decap_8
XFILLER_49_416 VPWR VGND sg13g2_decap_8
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_478 VPWR VGND sg13g2_decap_8
XFILLER_18_803 VPWR VGND sg13g2_decap_8
XFILLER_45_611 VPWR VGND sg13g2_decap_8
XFILLER_44_121 VPWR VGND sg13g2_fill_1
XFILLER_45_688 VPWR VGND sg13g2_decap_8
XFILLER_26_891 VPWR VGND sg13g2_decap_8
XFILLER_41_850 VPWR VGND sg13g2_decap_8
XFILLER_13_530 VPWR VGND sg13g2_decap_8
XFILLER_9_523 VPWR VGND sg13g2_decap_8
XFILLER_5_740 VPWR VGND sg13g2_decap_8
X_4170_ net773 VGND VPWR _0148_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[1\]
+ clknet_5_1__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3121_ VGND VPWR _0655_ _0657_ _0652_ net702 sg13g2_a21oi_2
XFILLER_49_983 VPWR VGND sg13g2_decap_8
X_3052_ _0593_ net734 net691 VPWR VGND sg13g2_nand2_1
XFILLER_48_493 VPWR VGND sg13g2_decap_8
XFILLER_36_633 VPWR VGND sg13g2_decap_8
XFILLER_23_305 VPWR VGND sg13g2_fill_1
XFILLER_24_806 VPWR VGND sg13g2_decap_8
Xclkbuf_4_13_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_13_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3954_ VGND VPWR net580 _0906_ _1385_ net604 sg13g2_a21oi_1
XFILLER_32_861 VPWR VGND sg13g2_decap_8
X_2905_ VPWR VGND _0469_ net554 _0468_ _1920_ _0470_ net616 sg13g2_a221oi_1
X_3885_ net762 _1460_ net765 _1326_ VPWR VGND sg13g2_a21o_1
X_2836_ VGND VPWR _0403_ _0401_ _0400_ sg13g2_or2_1
X_2767_ net563 VPWR _0336_ VGND net759 sap_3_inst.alu.tmp\[0\] sg13g2_o21ai_1
X_2698_ net567 _1986_ net11 VPWR VGND sg13g2_nor2b_2
XFILLER_6_90 VPWR VGND sg13g2_fill_2
Xfanout557 net558 net557 VPWR VGND sg13g2_buf_8
Xfanout546 _1975_ net546 VPWR VGND sg13g2_buf_8
Xfanout579 net582 net579 VPWR VGND sg13g2_buf_8
Xfanout568 _1139_ net568 VPWR VGND sg13g2_buf_8
X_3319_ VGND VPWR _0855_ _0854_ _0757_ sg13g2_or2_1
XFILLER_27_655 VPWR VGND sg13g2_decap_8
XFILLER_42_636 VPWR VGND sg13g2_decap_8
XFILLER_41_146 VPWR VGND sg13g2_fill_1
XFILLER_23_850 VPWR VGND sg13g2_decap_8
XFILLER_25_88 VPWR VGND sg13g2_fill_2
XFILLER_6_526 VPWR VGND sg13g2_decap_8
XFILLER_10_566 VPWR VGND sg13g2_decap_8
XFILLER_2_721 VPWR VGND sg13g2_decap_8
XFILLER_29_1007 VPWR VGND sg13g2_decap_8
XFILLER_2_798 VPWR VGND sg13g2_decap_8
XFILLER_2_37 VPWR VGND sg13g2_fill_1
XFILLER_49_279 VPWR VGND sg13g2_fill_2
XFILLER_46_920 VPWR VGND sg13g2_decap_8
XFILLER_18_600 VPWR VGND sg13g2_decap_8
XFILLER_18_677 VPWR VGND sg13g2_decap_8
XFILLER_46_997 VPWR VGND sg13g2_decap_8
XFILLER_45_485 VPWR VGND sg13g2_decap_8
XFILLER_33_669 VPWR VGND sg13g2_decap_8
XFILLER_14_894 VPWR VGND sg13g2_decap_8
XFILLER_32_168 VPWR VGND sg13g2_fill_1
Xclkbuf_4_5_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_5_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3670_ _1168_ net597 _1007_ VPWR VGND sg13g2_nand2b_1
XFILLER_12_1022 VPWR VGND sg13g2_decap_8
X_2621_ _0216_ _0217_ _0218_ VPWR VGND sg13g2_and2_1
X_2552_ _1965_ net4 _1847_ VPWR VGND sg13g2_nand2_1
X_2483_ _1899_ net22 VPWR VGND sg13g2_inv_4
X_4222_ mem_ram_we net25 VPWR VGND sg13g2_buf_1
XFILLER_29_909 VPWR VGND sg13g2_decap_8
X_4153_ net795 VGND VPWR _0131_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\]
+ clknet_5_28__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3104_ _0640_ _0613_ _0628_ _0639_ VPWR VGND sg13g2_and3_1
X_4084_ net770 VGND VPWR _0062_ sap_3_inst.controller.opcode\[3\] clknet_5_0__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_49_780 VPWR VGND sg13g2_decap_8
X_3035_ net18 net668 _0586_ VPWR VGND sg13g2_nor2_1
XFILLER_24_603 VPWR VGND sg13g2_decap_8
XFILLER_37_975 VPWR VGND sg13g2_decap_8
X_3937_ _1372_ _1305_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] _1302_
+ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_842 VPWR VGND sg13g2_decap_8
X_3868_ sap_3_inst.reg_file.array_serializer_inst.word_index\[0\] sap_3_inst.reg_file.array_serializer_inst.word_index\[1\]
+ sap_3_inst.reg_file.array_serializer_inst.word_index\[3\] sap_3_inst.reg_file.array_serializer_inst.word_index\[2\]
+ _1309_ VPWR VGND sg13g2_nor4_1
X_2819_ _0384_ _0385_ _0386_ VPWR VGND sg13g2_nor2b_1
X_3799_ VGND VPWR _1482_ net601 _0145_ _1256_ sg13g2_a21oi_1
XFILLER_3_507 VPWR VGND sg13g2_decap_8
XFILLER_11_68 VPWR VGND sg13g2_fill_2
XFILLER_47_717 VPWR VGND sg13g2_decap_8
XFILLER_28_953 VPWR VGND sg13g2_decap_8
XFILLER_43_901 VPWR VGND sg13g2_decap_8
XFILLER_27_452 VPWR VGND sg13g2_decap_8
XFILLER_36_87 VPWR VGND sg13g2_fill_1
XFILLER_43_978 VPWR VGND sg13g2_decap_8
XFILLER_42_433 VPWR VGND sg13g2_decap_8
XFILLER_15_647 VPWR VGND sg13g2_decap_8
XFILLER_6_301 VPWR VGND sg13g2_fill_2
XFILLER_11_886 VPWR VGND sg13g2_decap_8
XFILLER_7_846 VPWR VGND sg13g2_decap_8
XFILLER_2_595 VPWR VGND sg13g2_decap_8
XFILLER_38_739 VPWR VGND sg13g2_decap_8
XFILLER_18_430 VPWR VGND sg13g2_fill_2
XFILLER_19_964 VPWR VGND sg13g2_decap_8
XFILLER_46_794 VPWR VGND sg13g2_decap_8
XFILLER_45_271 VPWR VGND sg13g2_fill_2
XFILLER_34_956 VPWR VGND sg13g2_decap_8
XFILLER_14_691 VPWR VGND sg13g2_decap_8
XFILLER_21_639 VPWR VGND sg13g2_decap_8
X_3722_ _0119_ _1102_ _1205_ net594 _1472_ VPWR VGND sg13g2_a22oi_1
X_3653_ _1154_ net653 _0921_ VPWR VGND sg13g2_nand2_1
X_2604_ net618 _1951_ _0201_ VPWR VGND sg13g2_nor2_2
XFILLER_6_890 VPWR VGND sg13g2_decap_8
X_3584_ VGND VPWR _1920_ net570 _1100_ _1099_ sg13g2_a21oi_1
X_2535_ VGND VPWR net735 _1928_ _1948_ _1947_ sg13g2_a21oi_1
X_2466_ _1883_ net621 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[5\] net633
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4205_ net790 VGND VPWR _0182_ sap_3_inst.alu.act\[4\] clknet_5_23__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_4136_ net779 VGND VPWR _0114_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[7\]
+ clknet_5_15__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_2397_ VGND VPWR _1578_ _1640_ _1818_ _1612_ sg13g2_a21oi_1
XFILLER_29_706 VPWR VGND sg13g2_decap_8
X_4067_ net784 VGND VPWR _0045_ sap_3_inst.out\[3\] clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3018_ _0478_ _0507_ _0514_ _0540_ _0571_ VPWR VGND sg13g2_and4_1
XFILLER_24_400 VPWR VGND sg13g2_decap_8
XFILLER_25_912 VPWR VGND sg13g2_decap_8
XFILLER_37_772 VPWR VGND sg13g2_decap_8
XFILLER_19_1006 VPWR VGND sg13g2_decap_8
XFILLER_24_477 VPWR VGND sg13g2_decap_8
XFILLER_25_989 VPWR VGND sg13g2_decap_8
XFILLER_11_138 VPWR VGND sg13g2_fill_1
XFILLER_7_109 VPWR VGND sg13g2_decap_4
XFILLER_4_838 VPWR VGND sg13g2_decap_8
XFILLER_47_514 VPWR VGND sg13g2_decap_8
XFILLER_28_750 VPWR VGND sg13g2_decap_8
XFILLER_35_709 VPWR VGND sg13g2_decap_8
XFILLER_15_433 VPWR VGND sg13g2_fill_2
XFILLER_16_956 VPWR VGND sg13g2_decap_8
XFILLER_43_775 VPWR VGND sg13g2_decap_8
XFILLER_42_252 VPWR VGND sg13g2_fill_1
XFILLER_31_904 VPWR VGND sg13g2_decap_8
XFILLER_7_643 VPWR VGND sg13g2_decap_8
XFILLER_11_683 VPWR VGND sg13g2_decap_8
XFILLER_6_142 VPWR VGND sg13g2_fill_1
XFILLER_3_871 VPWR VGND sg13g2_decap_8
X_2320_ _1740_ VPWR _1741_ VGND _1735_ _1738_ sg13g2_o21ai_1
X_2251_ _1672_ net703 _1671_ VPWR VGND sg13g2_nand2_1
X_2182_ _1519_ _1567_ _1595_ _1603_ VPWR VGND sg13g2_nor3_1
XFILLER_38_536 VPWR VGND sg13g2_decap_8
XFILLER_26_709 VPWR VGND sg13g2_decap_8
XFILLER_19_761 VPWR VGND sg13g2_decap_8
XFILLER_46_591 VPWR VGND sg13g2_decap_8
XFILLER_33_230 VPWR VGND sg13g2_fill_1
XFILLER_34_753 VPWR VGND sg13g2_decap_8
XFILLER_22_904 VPWR VGND sg13g2_decap_8
XFILLER_33_241 VPWR VGND sg13g2_fill_2
X_3705_ _1194_ _1073_ net24 VPWR VGND sg13g2_nand2b_1
X_3636_ _1140_ net568 net31 VPWR VGND sg13g2_nand2b_1
X_3567_ _1086_ net576 _0880_ VPWR VGND sg13g2_nand2_2
X_2518_ net685 _1549_ _1930_ _1931_ VPWR VGND sg13g2_a21o_1
XFILLER_25_1010 VPWR VGND sg13g2_decap_8
X_3498_ _1027_ _1005_ _1020_ VPWR VGND sg13g2_xnor2_1
X_2449_ VPWR VGND net7 _1867_ _1847_ net745 _1868_ _1827_ sg13g2_a221oi_1
XFILLER_29_503 VPWR VGND sg13g2_decap_8
X_4119_ net796 VGND VPWR _0097_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\]
+ clknet_5_31__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_44_528 VPWR VGND sg13g2_decap_8
XFILLER_17_89 VPWR VGND sg13g2_fill_2
X_4027__5 VPWR net39 clknet_leaf_2_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_13_915 VPWR VGND sg13g2_decap_8
XFILLER_25_786 VPWR VGND sg13g2_decap_8
XFILLER_9_908 VPWR VGND sg13g2_decap_8
XFILLER_40_767 VPWR VGND sg13g2_decap_8
XFILLER_12_447 VPWR VGND sg13g2_fill_1
XFILLER_4_635 VPWR VGND sg13g2_decap_8
XFILLER_0_841 VPWR VGND sg13g2_decap_8
XFILLER_48_801 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_decap_4
Xhold7 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[2\] VPWR VGND net54 sg13g2_dlygate4sd3_1
XFILLER_48_878 VPWR VGND sg13g2_decap_8
XFILLER_47_388 VPWR VGND sg13g2_decap_8
XFILLER_35_506 VPWR VGND sg13g2_decap_8
XFILLER_16_753 VPWR VGND sg13g2_decap_8
XFILLER_31_701 VPWR VGND sg13g2_decap_8
XFILLER_43_572 VPWR VGND sg13g2_decap_8
XFILLER_31_778 VPWR VGND sg13g2_decap_8
XFILLER_8_930 VPWR VGND sg13g2_decap_8
XFILLER_7_473 VPWR VGND sg13g2_fill_2
X_3421_ VGND VPWR _0953_ _0952_ net579 sg13g2_or2_1
X_3352_ _0886_ _0877_ _0863_ _0068_ VPWR VGND sg13g2_a21o_1
X_2303_ _1724_ _1620_ _1698_ VPWR VGND sg13g2_nand2_1
X_3283_ _0815_ _0816_ _0817_ _0818_ _0819_ VPWR VGND sg13g2_and4_1
X_2234_ net729 _1507_ net722 _1655_ VPWR VGND sg13g2_nor3_2
XFILLER_39_845 VPWR VGND sg13g2_decap_8
X_2165_ _1585_ VPWR _1586_ VGND _1576_ _1579_ sg13g2_o21ai_1
XFILLER_26_506 VPWR VGND sg13g2_decap_8
X_2096_ VGND VPWR _1517_ net741 net739 sg13g2_or2_1
XFILLER_0_1023 VPWR VGND sg13g2_decap_4
XFILLER_38_399 VPWR VGND sg13g2_fill_2
XFILLER_22_701 VPWR VGND sg13g2_decap_8
XFILLER_34_550 VPWR VGND sg13g2_decap_8
XFILLER_22_778 VPWR VGND sg13g2_decap_8
X_2998_ net555 net743 _0559_ _0041_ VPWR VGND sg13g2_a21o_1
X_3619_ _0093_ _1128_ _1049_ net551 _1452_ VPWR VGND sg13g2_a22oi_1
XFILLER_29_355 VPWR VGND sg13g2_fill_2
XFILLER_17_528 VPWR VGND sg13g2_decap_8
XFILLER_13_712 VPWR VGND sg13g2_decap_8
XFILLER_25_583 VPWR VGND sg13g2_decap_8
XFILLER_44_98 VPWR VGND sg13g2_fill_2
XFILLER_9_705 VPWR VGND sg13g2_decap_8
XFILLER_40_564 VPWR VGND sg13g2_decap_8
XFILLER_13_789 VPWR VGND sg13g2_decap_8
XFILLER_5_922 VPWR VGND sg13g2_decap_8
XFILLER_5_999 VPWR VGND sg13g2_decap_8
XFILLER_48_675 VPWR VGND sg13g2_decap_8
XFILLER_36_815 VPWR VGND sg13g2_decap_8
X_3970_ _0321_ net759 net664 _1395_ VPWR VGND sg13g2_mux2_1
XFILLER_16_550 VPWR VGND sg13g2_decap_8
XFILLER_44_892 VPWR VGND sg13g2_decap_8
X_2921_ _0485_ net750 sap_3_inst.alu.tmp\[4\] VPWR VGND sg13g2_nand2b_1
X_2852_ VGND VPWR _0333_ _0416_ _0418_ net563 sg13g2_a21oi_1
XFILLER_31_575 VPWR VGND sg13g2_decap_8
X_2783_ VPWR VGND _0351_ net555 _0350_ net31 _0352_ net617 sg13g2_a221oi_1
X_3404_ _0936_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[4\] net562 VPWR
+ VGND sg13g2_nand2_1
Xfanout706 _1611_ net706 VPWR VGND sg13g2_buf_8
Xfanout739 sap_3_inst.controller.opcode\[1\] net739 VPWR VGND sg13g2_buf_8
Xfanout717 sap_3_inst.controller.stage\[2\] net717 VPWR VGND sg13g2_buf_8
Xfanout728 sap_3_inst.controller.opcode\[6\] net728 VPWR VGND sg13g2_buf_2
X_3335_ _0867_ _0868_ _0864_ _0870_ VPWR VGND _0869_ sg13g2_nand4_1
X_3266_ _0798_ _0799_ _0800_ _0801_ _0802_ VPWR VGND sg13g2_and4_1
X_2217_ net718 net705 _1638_ VPWR VGND sg13g2_and2_1
XFILLER_22_1002 VPWR VGND sg13g2_decap_8
XFILLER_39_642 VPWR VGND sg13g2_decap_8
X_3197_ _0658_ net665 _0711_ _0733_ VPWR VGND sg13g2_nor3_1
XFILLER_27_837 VPWR VGND sg13g2_decap_8
XFILLER_38_152 VPWR VGND sg13g2_fill_2
X_2148_ _1542_ _1555_ _1566_ _1569_ VGND VPWR _1568_ sg13g2_nor4_2
XFILLER_26_325 VPWR VGND sg13g2_fill_1
XFILLER_42_818 VPWR VGND sg13g2_decap_8
X_2079_ VGND VPWR _1500_ net716 net717 sg13g2_or2_1
XFILLER_14_509 VPWR VGND sg13g2_decap_8
XFILLER_35_870 VPWR VGND sg13g2_decap_8
XFILLER_22_575 VPWR VGND sg13g2_decap_8
XFILLER_6_708 VPWR VGND sg13g2_decap_8
XFILLER_10_748 VPWR VGND sg13g2_decap_8
XFILLER_2_903 VPWR VGND sg13g2_decap_8
XFILLER_7_1007 VPWR VGND sg13g2_decap_8
XFILLER_1_457 VPWR VGND sg13g2_decap_8
XFILLER_29_130 VPWR VGND sg13g2_fill_1
XFILLER_44_111 VPWR VGND sg13g2_fill_2
XFILLER_18_859 VPWR VGND sg13g2_decap_8
XFILLER_45_667 VPWR VGND sg13g2_decap_8
XFILLER_26_870 VPWR VGND sg13g2_decap_8
XFILLER_32_328 VPWR VGND sg13g2_fill_1
XFILLER_9_502 VPWR VGND sg13g2_decap_8
XFILLER_13_586 VPWR VGND sg13g2_decap_8
XFILLER_9_579 VPWR VGND sg13g2_decap_8
XFILLER_5_796 VPWR VGND sg13g2_decap_8
XFILLER_45_1024 VPWR VGND sg13g2_decap_4
X_3120_ VPWR _0656_ _0655_ VGND sg13g2_inv_1
XFILLER_49_962 VPWR VGND sg13g2_decap_8
XFILLER_48_472 VPWR VGND sg13g2_decap_8
X_3051_ VGND VPWR _1436_ net692 _0061_ _0592_ sg13g2_a21oi_1
XFILLER_36_612 VPWR VGND sg13g2_decap_8
XFILLER_17_892 VPWR VGND sg13g2_decap_8
XFILLER_36_689 VPWR VGND sg13g2_decap_8
X_3953_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] _1047_ net609 _0171_
+ VPWR VGND sg13g2_mux2_1
XFILLER_32_840 VPWR VGND sg13g2_decap_8
X_2904_ VGND VPWR sap_3_inst.alu.act\[4\] net669 _0469_ net616 sg13g2_a21oi_1
X_3884_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] _1324_
+ net721 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] _1325_ _1313_ sg13g2_a221oi_1
X_2835_ _0402_ _0400_ _0401_ VPWR VGND sg13g2_nand2_1
X_2766_ _0321_ VPWR _0335_ VGND net544 _0334_ sg13g2_o21ai_1
X_2697_ net567 _0213_ net10 VPWR VGND sg13g2_nor2b_2
Xfanout547 _1878_ net547 VPWR VGND sg13g2_buf_8
X_3318_ _0776_ _0788_ _0767_ _0854_ VPWR VGND _0849_ sg13g2_nand4_1
Xfanout558 _1037_ net558 VPWR VGND sg13g2_buf_8
Xfanout569 _1139_ net569 VPWR VGND sg13g2_buf_2
XFILLER_46_409 VPWR VGND sg13g2_decap_8
X_3249_ _0658_ net665 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[3\] _0785_
+ VPWR VGND net659 sg13g2_nand4_1
XFILLER_27_634 VPWR VGND sg13g2_decap_8
XFILLER_42_615 VPWR VGND sg13g2_decap_8
XFILLER_15_829 VPWR VGND sg13g2_decap_8
XFILLER_25_23 VPWR VGND sg13g2_fill_1
XFILLER_6_505 VPWR VGND sg13g2_decap_8
XFILLER_10_545 VPWR VGND sg13g2_decap_8
XFILLER_2_700 VPWR VGND sg13g2_decap_8
XFILLER_2_777 VPWR VGND sg13g2_decap_8
XFILLER_46_976 VPWR VGND sg13g2_decap_8
XFILLER_45_464 VPWR VGND sg13g2_decap_8
XFILLER_18_656 VPWR VGND sg13g2_decap_8
XFILLER_33_648 VPWR VGND sg13g2_decap_8
XFILLER_14_873 VPWR VGND sg13g2_decap_8
XFILLER_12_1001 VPWR VGND sg13g2_decap_8
X_2620_ _0217_ net624 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] net632
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2551_ _1964_ _1828_ sap_3_inst.alu.flags\[3\] _1827_ net754 VPWR VGND sg13g2_a22oi_1
X_2482_ _1899_ _1888_ _1889_ _1898_ VPWR VGND sg13g2_and3_2
XFILLER_5_593 VPWR VGND sg13g2_decap_8
X_4152_ net779 VGND VPWR _0130_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[7\]
+ clknet_5_15__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3103_ _1581_ _1620_ _1575_ _0639_ VPWR VGND sg13g2_nand3_1
X_4083_ net770 VGND VPWR _0061_ sap_3_inst.controller.opcode\[2\] clknet_5_5__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3034_ net17 sap_3_inst.alu.tmp\[0\] net668 _0051_ VPWR VGND sg13g2_mux2_1
XFILLER_37_954 VPWR VGND sg13g2_decap_8
XFILLER_24_659 VPWR VGND sg13g2_decap_8
X_3936_ _1371_ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[6\] _1308_
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_821 VPWR VGND sg13g2_decap_8
X_3867_ _1300_ _1307_ _1308_ VPWR VGND sg13g2_nor2_2
XFILLER_31_191 VPWR VGND sg13g2_fill_1
X_2818_ _0367_ _0382_ _0353_ _0385_ VPWR VGND sg13g2_nand3_1
XFILLER_20_898 VPWR VGND sg13g2_decap_8
X_3798_ net601 _1002_ _1071_ _1256_ VPWR VGND sg13g2_nor3_1
X_2749_ _0315_ VPWR _0318_ VGND _0311_ net670 sg13g2_o21ai_1
XFILLER_46_228 VPWR VGND sg13g2_fill_2
XFILLER_28_932 VPWR VGND sg13g2_decap_8
XFILLER_27_431 VPWR VGND sg13g2_decap_8
XFILLER_15_626 VPWR VGND sg13g2_decap_8
XFILLER_43_957 VPWR VGND sg13g2_decap_8
XFILLER_42_489 VPWR VGND sg13g2_decap_8
XFILLER_10_353 VPWR VGND sg13g2_fill_1
XFILLER_7_825 VPWR VGND sg13g2_decap_8
XFILLER_11_865 VPWR VGND sg13g2_decap_8
Xclkbuf_5_31__f_sap_3_inst.alu.clk_regs clknet_4_15_0_sap_3_inst.alu.clk_regs clknet_5_31__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_2_574 VPWR VGND sg13g2_decap_8
XFILLER_38_718 VPWR VGND sg13g2_decap_8
XFILLER_19_943 VPWR VGND sg13g2_decap_8
XFILLER_46_773 VPWR VGND sg13g2_decap_8
XFILLER_34_935 VPWR VGND sg13g2_decap_8
XFILLER_21_618 VPWR VGND sg13g2_decap_8
XFILLER_14_670 VPWR VGND sg13g2_decap_8
X_3721_ net594 _1059_ _1205_ VPWR VGND sg13g2_nor2_1
X_3652_ VPWR VGND _0933_ _0929_ _1152_ _1150_ _1153_ _1151_ sg13g2_a221oi_1
X_2603_ _1936_ _1945_ _0200_ VPWR VGND sg13g2_nor2_2
X_3583_ net13 net570 _1099_ VPWR VGND sg13g2_nor2_1
X_2534_ _1550_ _1747_ _1947_ VPWR VGND sg13g2_nor2_2
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_2465_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] net635
+ _1882_ net638 sg13g2_a21oi_1
X_4204_ net789 VGND VPWR _0181_ sap_3_inst.alu.act\[3\] clknet_5_21__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_2396_ net724 _1559_ _1584_ _1817_ VPWR VGND sg13g2_nor3_1
XFILLER_3_92 VPWR VGND sg13g2_decap_8
X_4135_ net796 VGND VPWR _0113_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\]
+ clknet_5_30__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4066_ net784 VGND VPWR _0044_ sap_3_inst.out\[2\] clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_37_751 VPWR VGND sg13g2_decap_8
X_3017_ _0570_ _0447_ _0569_ VPWR VGND sg13g2_nand2_1
XFILLER_25_968 VPWR VGND sg13g2_decap_8
XFILLER_24_456 VPWR VGND sg13g2_decap_8
XFILLER_40_949 VPWR VGND sg13g2_decap_8
X_3919_ _1356_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[4\] _1311_
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_4_817 VPWR VGND sg13g2_decap_8
XFILLER_20_695 VPWR VGND sg13g2_decap_8
XFILLER_16_935 VPWR VGND sg13g2_decap_8
XFILLER_43_754 VPWR VGND sg13g2_decap_8
XFILLER_7_622 VPWR VGND sg13g2_decap_8
XFILLER_11_662 VPWR VGND sg13g2_decap_8
XFILLER_6_132 VPWR VGND sg13g2_fill_2
XFILLER_7_699 VPWR VGND sg13g2_decap_8
XFILLER_6_198 VPWR VGND sg13g2_fill_2
XFILLER_3_850 VPWR VGND sg13g2_decap_8
XFILLER_2_360 VPWR VGND sg13g2_fill_1
X_2250_ _1538_ VPWR _1671_ VGND _1548_ _1670_ sg13g2_o21ai_1
X_2181_ VGND VPWR _1602_ _1601_ _1594_ sg13g2_or2_1
XFILLER_38_515 VPWR VGND sg13g2_decap_8
XFILLER_19_740 VPWR VGND sg13g2_decap_8
XFILLER_46_570 VPWR VGND sg13g2_decap_8
XFILLER_34_732 VPWR VGND sg13g2_decap_8
XFILLER_15_990 VPWR VGND sg13g2_decap_8
X_3704_ _1191_ VPWR _0113_ VGND _1181_ _1193_ sg13g2_o21ai_1
X_3635_ _1139_ net652 _0836_ VPWR VGND sg13g2_nand2b_1
X_3566_ net32 net10 _1078_ _1085_ VPWR VGND sg13g2_mux2_1
X_3497_ VGND VPWR net610 _1024_ _1026_ net576 sg13g2_a21oi_1
X_2517_ _1930_ net682 _1929_ VPWR VGND sg13g2_nand2b_1
X_2448_ sap_3_inst.alu.flags\[6\] _1828_ _1867_ VPWR VGND sg13g2_and2_1
X_2379_ _1800_ net662 _1761_ _1792_ VPWR VGND sg13g2_and3_2
X_4118_ net776 VGND VPWR _0096_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\]
+ clknet_5_14__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_559 VPWR VGND sg13g2_decap_8
XFILLER_44_507 VPWR VGND sg13g2_decap_8
X_4049_ net772 VGND VPWR _0003_ sap_3_inst.controller.stage\[1\] net41 sg13g2_dfrbpq_2
XFILLER_24_220 VPWR VGND sg13g2_fill_1
XFILLER_25_765 VPWR VGND sg13g2_decap_8
XFILLER_40_746 VPWR VGND sg13g2_decap_8
XFILLER_21_982 VPWR VGND sg13g2_decap_8
XFILLER_32_1015 VPWR VGND sg13g2_decap_8
XFILLER_20_492 VPWR VGND sg13g2_decap_8
XFILLER_4_614 VPWR VGND sg13g2_decap_8
XFILLER_0_820 VPWR VGND sg13g2_decap_8
XFILLER_0_897 VPWR VGND sg13g2_decap_8
Xhold8 sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[5\] VPWR VGND net55 sg13g2_dlygate4sd3_1
XFILLER_48_857 VPWR VGND sg13g2_decap_8
XFILLER_47_367 VPWR VGND sg13g2_decap_8
XFILLER_16_732 VPWR VGND sg13g2_decap_8
XFILLER_43_551 VPWR VGND sg13g2_decap_8
XFILLER_30_201 VPWR VGND sg13g2_fill_2
XFILLER_31_757 VPWR VGND sg13g2_decap_8
XFILLER_8_986 VPWR VGND sg13g2_decap_8
XFILLER_48_1011 VPWR VGND sg13g2_decap_8
X_3420_ net574 _0852_ _0951_ _0952_ VPWR VGND sg13g2_nor3_1
X_3351_ _0879_ _0880_ net576 _0886_ VPWR VGND _0884_ sg13g2_nand4_1
Xclkbuf_5_28__f_sap_3_inst.alu.clk_regs clknet_4_14_0_sap_3_inst.alu.clk_regs clknet_5_28__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2302_ _1723_ _1537_ net567 _1722_ VPWR VGND sg13g2_and3_2
X_3282_ _0672_ _0712_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] _0818_
+ VPWR VGND sg13g2_nand3_1
X_2233_ _1654_ _1647_ _1579_ _1593_ _1590_ VPWR VGND sg13g2_a22oi_1
XFILLER_39_824 VPWR VGND sg13g2_decap_8
X_2164_ _1585_ _1581_ _1583_ VPWR VGND sg13g2_nand2_1
XFILLER_0_1002 VPWR VGND sg13g2_decap_8
X_2095_ net740 net741 _1516_ VPWR VGND sg13g2_nor2_1
XFILLER_0_71 VPWR VGND sg13g2_fill_2
XFILLER_21_223 VPWR VGND sg13g2_fill_2
XFILLER_22_757 VPWR VGND sg13g2_decap_8
XFILLER_9_80 VPWR VGND sg13g2_decap_4
X_2997_ net555 _0533_ _0558_ _0559_ VPWR VGND sg13g2_nor3_1
XFILLER_21_267 VPWR VGND sg13g2_fill_1
X_3618_ _1050_ net551 _1128_ VPWR VGND sg13g2_nor2_1
XFILLER_1_639 VPWR VGND sg13g2_decap_8
X_3549_ VGND VPWR _1071_ _1070_ _1068_ sg13g2_or2_1
XFILLER_17_507 VPWR VGND sg13g2_decap_8
XFILLER_45_849 VPWR VGND sg13g2_decap_8
XFILLER_44_348 VPWR VGND sg13g2_fill_2
XFILLER_44_359 VPWR VGND sg13g2_decap_4
XFILLER_25_562 VPWR VGND sg13g2_decap_8
XFILLER_40_543 VPWR VGND sg13g2_decap_8
XFILLER_13_768 VPWR VGND sg13g2_decap_8
XFILLER_5_901 VPWR VGND sg13g2_decap_8
XFILLER_5_27 VPWR VGND sg13g2_decap_8
XFILLER_5_978 VPWR VGND sg13g2_decap_8
XFILLER_4_488 VPWR VGND sg13g2_decap_8
XFILLER_48_654 VPWR VGND sg13g2_decap_8
XFILLER_0_694 VPWR VGND sg13g2_decap_8
XFILLER_44_871 VPWR VGND sg13g2_decap_8
X_2920_ _0483_ VPWR _0484_ VGND net748 _0327_ sg13g2_o21ai_1
XFILLER_31_554 VPWR VGND sg13g2_decap_8
X_2851_ net753 sap_3_inst.alu.tmp\[3\] _0417_ VPWR VGND sg13g2_nor2_1
X_2782_ VGND VPWR _1462_ net670 _0351_ net617 sg13g2_a21oi_1
XFILLER_8_783 VPWR VGND sg13g2_decap_8
X_3403_ _0908_ VPWR _0070_ VGND _0925_ _0934_ sg13g2_o21ai_1
Xfanout707 net708 net707 VPWR VGND sg13g2_buf_8
Xfanout718 sap_3_inst.controller.stage\[1\] net718 VPWR VGND sg13g2_buf_8
Xfanout729 sap_3_inst.controller.opcode\[5\] net729 VPWR VGND sg13g2_buf_8
X_3334_ _0869_ net588 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[1\] net592
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[1\] VPWR VGND sg13g2_a22oi_1
X_3265_ _0695_ _0719_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[2\] _0801_
+ VPWR VGND sg13g2_nand3_1
X_2216_ _1637_ _1636_ VPWR VGND sg13g2_inv_2
XFILLER_39_621 VPWR VGND sg13g2_decap_8
X_3196_ _0657_ _0670_ _0711_ _0732_ VPWR VGND sg13g2_nor3_1
XFILLER_27_816 VPWR VGND sg13g2_decap_8
X_2147_ _1509_ _1562_ _1568_ VPWR VGND sg13g2_nor2_2
XFILLER_39_698 VPWR VGND sg13g2_decap_8
X_2078_ net717 net716 _1499_ VPWR VGND sg13g2_nor2_2
XFILLER_10_727 VPWR VGND sg13g2_decap_8
XFILLER_22_554 VPWR VGND sg13g2_decap_8
XFILLER_2_959 VPWR VGND sg13g2_decap_8
XFILLER_45_646 VPWR VGND sg13g2_decap_8
XFILLER_17_337 VPWR VGND sg13g2_fill_1
XFILLER_18_838 VPWR VGND sg13g2_decap_8
XFILLER_41_885 VPWR VGND sg13g2_decap_8
XFILLER_13_565 VPWR VGND sg13g2_decap_8
XFILLER_9_558 VPWR VGND sg13g2_decap_8
XFILLER_5_775 VPWR VGND sg13g2_decap_8
XFILLER_45_1003 VPWR VGND sg13g2_decap_8
XFILLER_49_941 VPWR VGND sg13g2_decap_8
XFILLER_0_491 VPWR VGND sg13g2_decap_8
X_3050_ net692 net19 _0592_ VPWR VGND sg13g2_nor2_1
XFILLER_48_451 VPWR VGND sg13g2_decap_8
XFILLER_36_668 VPWR VGND sg13g2_decap_8
XFILLER_17_871 VPWR VGND sg13g2_decap_8
X_3952_ net604 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[0\] _1384_ _0170_
+ VPWR VGND sg13g2_a21o_1
X_2903_ _0468_ _0466_ _0467_ VPWR VGND sg13g2_nand2_1
X_3883_ _1324_ _1323_ _1322_ VPWR VGND sg13g2_nand2b_1
X_2834_ VGND VPWR net760 _0371_ _0401_ _0370_ sg13g2_a21oi_1
XFILLER_32_896 VPWR VGND sg13g2_decap_8
XFILLER_8_580 VPWR VGND sg13g2_decap_8
X_2765_ VGND VPWR _0334_ _0333_ _0322_ sg13g2_or2_1
X_2696_ net566 _0236_ net9 VPWR VGND sg13g2_nor2b_2
XFILLER_6_92 VPWR VGND sg13g2_fill_1
Xfanout548 net549 net548 VPWR VGND sg13g2_buf_8
X_3317_ _0788_ _0849_ _0776_ _0853_ VPWR VGND sg13g2_nand3_1
Xfanout559 net560 net559 VPWR VGND sg13g2_buf_8
X_3248_ _0672_ net659 sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[3\] _0784_
+ VPWR VGND sg13g2_nand3_1
XFILLER_27_613 VPWR VGND sg13g2_decap_8
X_3179_ _0715_ _0672_ net659 VPWR VGND sg13g2_nand2_2
XFILLER_39_495 VPWR VGND sg13g2_decap_8
XFILLER_15_808 VPWR VGND sg13g2_decap_8
XFILLER_26_167 VPWR VGND sg13g2_decap_8
XFILLER_41_126 VPWR VGND sg13g2_fill_2
XFILLER_25_57 VPWR VGND sg13g2_fill_1
XFILLER_23_885 VPWR VGND sg13g2_decap_8
XFILLER_10_524 VPWR VGND sg13g2_decap_8
XFILLER_2_756 VPWR VGND sg13g2_decap_8
XFILLER_18_635 VPWR VGND sg13g2_decap_8
XFILLER_46_955 VPWR VGND sg13g2_decap_8
XFILLER_45_443 VPWR VGND sg13g2_decap_8
XFILLER_33_627 VPWR VGND sg13g2_decap_8
XFILLER_14_852 VPWR VGND sg13g2_decap_8
XFILLER_41_682 VPWR VGND sg13g2_decap_8
X_2550_ _1963_ _1958_ _1962_ net637 _1440_ VPWR VGND sg13g2_a22oi_1
X_2481_ VGND VPWR _1723_ _1887_ _1898_ _1897_ sg13g2_a21oi_1
XFILLER_5_572 VPWR VGND sg13g2_decap_8
X_4151_ net780 VGND VPWR _0129_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[6\]
+ clknet_5_30__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4082_ net785 VGND VPWR _0060_ sap_3_inst.controller.opcode\[1\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_3102_ net714 net704 net731 _0638_ VPWR VGND sg13g2_nand3_1
X_3033_ _1843_ VPWR _0585_ VGND _1836_ _0584_ sg13g2_o21ai_1
XFILLER_37_933 VPWR VGND sg13g2_decap_8
XFILLER_24_638 VPWR VGND sg13g2_decap_8
XFILLER_20_800 VPWR VGND sg13g2_decap_8
X_3935_ _1370_ _1316_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] _1313_
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_32_693 VPWR VGND sg13g2_decap_8
X_3866_ _1307_ _1497_ net768 VPWR VGND sg13g2_nand2_2
XFILLER_20_877 VPWR VGND sg13g2_decap_8
X_3797_ net599 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[5\] _1255_ _0144_
+ VPWR VGND sg13g2_a21o_1
X_2817_ VGND VPWR _0353_ _0367_ _0384_ _0382_ sg13g2_a21oi_1
X_2748_ _0317_ _0202_ _0316_ VPWR VGND sg13g2_nand2b_1
X_2679_ _0269_ _0270_ _0268_ _0271_ VPWR VGND sg13g2_nand3_1
Xclkbuf_5_2__f_sap_3_inst.alu.clk_regs clknet_4_1_0_sap_3_inst.alu.clk_regs clknet_5_2__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_28_911 VPWR VGND sg13g2_decap_8
XFILLER_27_421 VPWR VGND sg13g2_fill_1
XFILLER_43_936 VPWR VGND sg13g2_decap_8
XFILLER_15_605 VPWR VGND sg13g2_decap_8
XFILLER_27_487 VPWR VGND sg13g2_decap_8
XFILLER_28_988 VPWR VGND sg13g2_decap_8
XFILLER_42_468 VPWR VGND sg13g2_decap_8
XFILLER_30_619 VPWR VGND sg13g2_decap_8
XFILLER_23_682 VPWR VGND sg13g2_decap_8
XFILLER_35_1024 VPWR VGND sg13g2_decap_4
XFILLER_7_804 VPWR VGND sg13g2_decap_8
XFILLER_11_844 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_4
XFILLER_2_553 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_19_922 VPWR VGND sg13g2_decap_8
XFILLER_46_752 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_sap_3_inst.alu.clk clknet_1_0__leaf_sap_3_inst.alu.clk clknet_leaf_0_sap_3_inst.alu.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_19_999 VPWR VGND sg13g2_decap_8
XFILLER_34_914 VPWR VGND sg13g2_decap_8
XFILLER_45_273 VPWR VGND sg13g2_fill_1
XFILLER_33_435 VPWR VGND sg13g2_fill_2
X_3720_ VPWR _0118_ _1204_ VGND sg13g2_inv_1
XFILLER_13_181 VPWR VGND sg13g2_fill_1
XFILLER_9_163 VPWR VGND sg13g2_fill_2
X_3651_ _1152_ _0727_ _0935_ VPWR VGND sg13g2_nand2_1
X_2602_ _0197_ _0198_ net564 _0199_ VPWR VGND sg13g2_nand3_1
X_3582_ _1098_ VPWR _0086_ VGND _1443_ net593 sg13g2_o21ai_1
X_2533_ _1943_ _1944_ _1946_ VPWR VGND sg13g2_nor2_2
X_2464_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] _1880_
+ net625 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] _1881_ net627 sg13g2_a221oi_1
X_4203_ net789 VGND VPWR _0180_ sap_3_inst.alu.act\[2\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_2395_ net736 _1815_ _1816_ VPWR VGND sg13g2_nor2_1
X_4134_ net779 VGND VPWR _0112_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_3_71 VPWR VGND sg13g2_decap_4
XFILLER_3_1011 VPWR VGND sg13g2_decap_8
XFILLER_28_229 VPWR VGND sg13g2_fill_1
X_4065_ net783 VGND VPWR _0043_ sap_3_inst.out\[1\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_37_730 VPWR VGND sg13g2_decap_8
X_3016_ _0569_ _0479_ _0507_ _0540_ VPWR VGND sg13g2_and3_1
XFILLER_24_435 VPWR VGND sg13g2_decap_8
XFILLER_25_947 VPWR VGND sg13g2_decap_8
XFILLER_40_928 VPWR VGND sg13g2_decap_8
XFILLER_11_118 VPWR VGND sg13g2_fill_1
XFILLER_33_991 VPWR VGND sg13g2_decap_8
XFILLER_32_490 VPWR VGND sg13g2_decap_8
X_3918_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[4\] _1302_
+ _1355_ net763 sg13g2_a21oi_1
XFILLER_20_674 VPWR VGND sg13g2_decap_8
X_3849_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[0\] sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\]
+ _1291_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_47_549 VPWR VGND sg13g2_decap_8
XFILLER_16_914 VPWR VGND sg13g2_decap_8
XFILLER_28_785 VPWR VGND sg13g2_decap_8
XFILLER_43_733 VPWR VGND sg13g2_decap_8
XFILLER_15_435 VPWR VGND sg13g2_fill_1
XFILLER_27_273 VPWR VGND sg13g2_fill_1
XFILLER_31_939 VPWR VGND sg13g2_decap_8
XFILLER_11_641 VPWR VGND sg13g2_decap_8
XFILLER_7_601 VPWR VGND sg13g2_decap_8
XFILLER_7_678 VPWR VGND sg13g2_decap_8
XFILLER_12_91 VPWR VGND sg13g2_fill_1
X_2180_ VGND VPWR _1601_ _1599_ _1596_ sg13g2_or2_1
XFILLER_34_711 VPWR VGND sg13g2_decap_8
XFILLER_19_796 VPWR VGND sg13g2_decap_8
XFILLER_22_939 VPWR VGND sg13g2_decap_8
XFILLER_34_788 VPWR VGND sg13g2_decap_8
XFILLER_30_983 VPWR VGND sg13g2_decap_8
X_3703_ _1192_ VPWR _1193_ VGND net581 _1071_ sg13g2_o21ai_1
X_3634_ _0847_ VPWR _1138_ VGND _0828_ _0830_ sg13g2_o21ai_1
X_3565_ net590 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] _1084_ _0083_
+ VPWR VGND sg13g2_a21o_1
X_3496_ net576 _1024_ _1025_ VPWR VGND sg13g2_nor2_1
X_2516_ net694 _1550_ _1716_ _1929_ VPWR VGND sg13g2_nor3_1
X_2447_ _1866_ _1861_ _1865_ net639 _1479_ VPWR VGND sg13g2_a22oi_1
X_2378_ _1799_ net662 _1762_ _1790_ VPWR VGND sg13g2_and3_2
X_4117_ net776 VGND VPWR _0095_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\]
+ clknet_5_9__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_538 VPWR VGND sg13g2_decap_8
X_4048_ net770 VGND VPWR _0002_ sap_3_inst.controller.stage\[0\] net40 sg13g2_dfrbpq_2
XFILLER_25_744 VPWR VGND sg13g2_decap_8
XFILLER_40_725 VPWR VGND sg13g2_decap_8
XFILLER_21_961 VPWR VGND sg13g2_decap_8
XFILLER_3_103 VPWR VGND sg13g2_fill_1
XFILLER_3_136 VPWR VGND sg13g2_decap_8
XFILLER_48_836 VPWR VGND sg13g2_decap_8
Xhold9 u_ser.shadow_reg\[6\] VPWR VGND net56 sg13g2_dlygate4sd3_1
XFILLER_0_876 VPWR VGND sg13g2_decap_8
XFILLER_47_346 VPWR VGND sg13g2_decap_8
XFILLER_16_711 VPWR VGND sg13g2_decap_8
XFILLER_28_582 VPWR VGND sg13g2_decap_8
XFILLER_43_530 VPWR VGND sg13g2_decap_8
XFILLER_16_788 VPWR VGND sg13g2_decap_8
XFILLER_31_736 VPWR VGND sg13g2_decap_8
XFILLER_8_965 VPWR VGND sg13g2_decap_8
XFILLER_12_994 VPWR VGND sg13g2_decap_8
XFILLER_7_475 VPWR VGND sg13g2_fill_1
X_3350_ VPWR _0885_ _0884_ VGND sg13g2_inv_1
X_2301_ net703 VPWR _1722_ VGND _1676_ _1721_ sg13g2_o21ai_1
X_3281_ net659 _0719_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] _0817_
+ VPWR VGND sg13g2_nand3_1
XFILLER_39_803 VPWR VGND sg13g2_decap_8
X_2232_ _1653_ _1652_ _1615_ _1643_ net707 VPWR VGND sg13g2_a22oi_1
X_2163_ _1584_ _1573_ VPWR VGND _1567_ sg13g2_nand2b_2
XFILLER_0_50 VPWR VGND sg13g2_decap_8
X_2094_ _1504_ _1510_ _1515_ VPWR VGND net733 sg13g2_nand3b_1
XFILLER_19_593 VPWR VGND sg13g2_decap_8
XFILLER_22_736 VPWR VGND sg13g2_decap_8
XFILLER_34_585 VPWR VGND sg13g2_decap_8
XFILLER_10_909 VPWR VGND sg13g2_decap_8
X_2996_ VPWR VGND _0557_ _0310_ _0556_ sap_3_inst.alu.act\[7\] _0558_ net669 sg13g2_a221oi_1
XFILLER_9_92 VPWR VGND sg13g2_decap_4
XFILLER_30_780 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_clk_div_out clknet_0_clk_div_out clknet_1_1__leaf_clk_div_out VPWR
+ VGND sg13g2_buf_8
X_3617_ _1047_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] net550 _0092_
+ VPWR VGND sg13g2_mux2_1
X_3548_ VGND VPWR _0757_ _0854_ _1070_ _1069_ sg13g2_a21oi_1
XFILLER_0_117 VPWR VGND sg13g2_fill_1
XFILLER_1_618 VPWR VGND sg13g2_decap_8
XFILLER_0_139 VPWR VGND sg13g2_fill_1
X_3479_ VPWR _1009_ _1008_ VGND sg13g2_inv_1
XFILLER_28_46 VPWR VGND sg13g2_fill_1
XFILLER_45_828 VPWR VGND sg13g2_decap_8
XFILLER_44_305 VPWR VGND sg13g2_fill_2
XFILLER_25_541 VPWR VGND sg13g2_decap_8
XFILLER_40_522 VPWR VGND sg13g2_decap_8
XFILLER_13_747 VPWR VGND sg13g2_decap_8
XFILLER_40_599 VPWR VGND sg13g2_decap_8
XFILLER_5_957 VPWR VGND sg13g2_decap_8
XFILLER_4_467 VPWR VGND sg13g2_decap_8
XFILLER_0_673 VPWR VGND sg13g2_decap_8
XFILLER_48_633 VPWR VGND sg13g2_decap_8
XFILLER_44_850 VPWR VGND sg13g2_decap_8
XFILLER_16_585 VPWR VGND sg13g2_decap_8
X_2850_ _0416_ net753 sap_3_inst.alu.tmp\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_31_533 VPWR VGND sg13g2_decap_8
XFILLER_15_1011 VPWR VGND sg13g2_decap_8
X_2781_ _0347_ _0349_ _0335_ _0350_ VPWR VGND sg13g2_nand3_1
XFILLER_12_791 VPWR VGND sg13g2_decap_8
XFILLER_8_762 VPWR VGND sg13g2_decap_8
X_3402_ _0935_ _0787_ _0822_ VPWR VGND sg13g2_xnor2_1
Xfanout708 _1603_ net708 VPWR VGND sg13g2_buf_8
Xfanout719 sap_3_inst.controller.stage\[0\] net719 VPWR VGND sg13g2_buf_8
X_3333_ _0868_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\] net641 VPWR
+ VGND sg13g2_nand2_1
XFILLER_22_0 VPWR VGND sg13g2_fill_2
X_3264_ _0800_ net650 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[2\] net653
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_600 VPWR VGND sg13g2_decap_8
X_2215_ _1636_ net716 _1635_ VPWR VGND sg13g2_nand2_2
X_3195_ _0731_ _0658_ net665 VPWR VGND sg13g2_nand2_1
XFILLER_39_677 VPWR VGND sg13g2_decap_8
X_2146_ net726 net728 net738 _1567_ VPWR VGND sg13g2_nand3_1
XFILLER_22_533 VPWR VGND sg13g2_decap_8
XFILLER_10_706 VPWR VGND sg13g2_decap_8
X_2979_ VGND VPWR net746 _1467_ _0541_ _0509_ sg13g2_a21oi_1
XFILLER_2_938 VPWR VGND sg13g2_decap_8
XFILLER_18_817 VPWR VGND sg13g2_decap_8
XFILLER_45_625 VPWR VGND sg13g2_decap_8
XFILLER_44_113 VPWR VGND sg13g2_fill_1
XFILLER_17_305 VPWR VGND sg13g2_fill_1
XFILLER_29_176 VPWR VGND sg13g2_fill_1
XFILLER_29_198 VPWR VGND sg13g2_fill_2
XFILLER_33_809 VPWR VGND sg13g2_decap_8
XFILLER_44_157 VPWR VGND sg13g2_fill_2
XFILLER_13_544 VPWR VGND sg13g2_decap_8
XFILLER_25_382 VPWR VGND sg13g2_decap_8
XFILLER_41_864 VPWR VGND sg13g2_decap_8
XFILLER_9_537 VPWR VGND sg13g2_decap_8
XFILLER_5_754 VPWR VGND sg13g2_decap_8
XFILLER_49_920 VPWR VGND sg13g2_decap_8
XFILLER_0_470 VPWR VGND sg13g2_decap_8
XFILLER_1_982 VPWR VGND sg13g2_decap_8
XFILLER_48_430 VPWR VGND sg13g2_decap_8
XFILLER_49_997 VPWR VGND sg13g2_decap_8
XFILLER_17_850 VPWR VGND sg13g2_decap_8
XFILLER_36_647 VPWR VGND sg13g2_decap_8
X_3951_ net604 _1040_ _1041_ _1384_ VPWR VGND sg13g2_nor3_1
X_2902_ VGND VPWR net544 _0450_ _0467_ _0314_ sg13g2_a21oi_1
XFILLER_32_875 VPWR VGND sg13g2_decap_8
X_3882_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] _1317_
+ _1323_ net762 sg13g2_a21oi_1
X_2833_ _0400_ net756 _1947_ VPWR VGND sg13g2_xnor2_1
X_2764_ _0197_ net618 _0333_ VPWR VGND sg13g2_nor2b_2
X_2695_ _1637_ _0282_ _0283_ _0005_ VPWR VGND sg13g2_nor3_1
X_3316_ _0775_ _0851_ _0852_ VPWR VGND sg13g2_nor2_1
Xfanout549 _1394_ net549 VPWR VGND sg13g2_buf_8
X_3247_ net659 _0719_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\] _0783_
+ VPWR VGND sg13g2_nand3_1
X_3178_ _0673_ _0713_ _0714_ VPWR VGND sg13g2_nor2_1
XFILLER_39_474 VPWR VGND sg13g2_decap_8
X_2129_ net737 _1520_ _1550_ VPWR VGND net739 sg13g2_nand3b_1
XFILLER_27_669 VPWR VGND sg13g2_decap_8
XFILLER_23_864 VPWR VGND sg13g2_decap_8
XFILLER_10_503 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_fill_2
XFILLER_2_735 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_46_934 VPWR VGND sg13g2_decap_8
XFILLER_18_614 VPWR VGND sg13g2_decap_8
XFILLER_45_422 VPWR VGND sg13g2_decap_8
XFILLER_33_606 VPWR VGND sg13g2_decap_8
XFILLER_45_499 VPWR VGND sg13g2_decap_8
XFILLER_14_831 VPWR VGND sg13g2_decap_8
XFILLER_41_661 VPWR VGND sg13g2_decap_8
XFILLER_13_330 VPWR VGND sg13g2_fill_1
X_2480_ VGND VPWR _1892_ _1896_ _1897_ net565 sg13g2_a21oi_1
XFILLER_5_551 VPWR VGND sg13g2_decap_8
X_4150_ net779 VGND VPWR _0128_ sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\]
+ clknet_5_12__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_3101_ _1549_ net687 net731 _0637_ VPWR VGND sg13g2_nand3_1
X_4081_ net770 VGND VPWR _0059_ sap_3_inst.controller.opcode\[0\] clknet_5_4__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_49_794 VPWR VGND sg13g2_decap_8
X_3032_ _0584_ _1545_ _1729_ VPWR VGND sg13g2_nand2_1
XFILLER_37_912 VPWR VGND sg13g2_decap_8
XFILLER_24_617 VPWR VGND sg13g2_decap_8
XFILLER_37_989 VPWR VGND sg13g2_decap_8
XFILLER_23_127 VPWR VGND sg13g2_fill_2
X_3934_ _1369_ _1315_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] _1306_
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] VPWR VGND sg13g2_a22oi_1
X_3865_ _1497_ net768 sap_3_inst.reg_file.array_serializer_inst.word_index\[3\] _1306_
+ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.word_index\[2\] sg13g2_nor4_2
XFILLER_32_672 VPWR VGND sg13g2_decap_8
X_2816_ VPWR _0383_ _0382_ VGND sg13g2_inv_1
XFILLER_20_856 VPWR VGND sg13g2_decap_8
X_3796_ net598 _1133_ _1134_ _1255_ VPWR VGND sg13g2_nor3_1
X_2747_ net618 _1951_ _0316_ VPWR VGND sg13g2_and2_1
X_2678_ _1605_ VPWR _0270_ VGND net696 _1637_ sg13g2_o21ai_1
XFILLER_28_967 VPWR VGND sg13g2_decap_8
XFILLER_43_915 VPWR VGND sg13g2_decap_8
XFILLER_27_466 VPWR VGND sg13g2_decap_8
XFILLER_42_447 VPWR VGND sg13g2_decap_8
XFILLER_35_1003 VPWR VGND sg13g2_decap_8
XFILLER_11_823 VPWR VGND sg13g2_decap_8
XFILLER_23_661 VPWR VGND sg13g2_decap_8
XFILLER_2_532 VPWR VGND sg13g2_decap_8
XFILLER_42_1007 VPWR VGND sg13g2_decap_8
XFILLER_19_901 VPWR VGND sg13g2_decap_8
XFILLER_46_731 VPWR VGND sg13g2_decap_8
XFILLER_19_978 VPWR VGND sg13g2_decap_8
XFILLER_9_153 VPWR VGND sg13g2_fill_1
X_3650_ VGND VPWR _1151_ net569 net12 sg13g2_or2_1
X_2601_ _0198_ _1943_ _1944_ VPWR VGND sg13g2_nand2_2
X_3581_ net593 _0921_ _1098_ VPWR VGND _1097_ sg13g2_nand3b_1
X_2532_ _1945_ _1943_ VPWR VGND _1944_ sg13g2_nand2b_2
X_2463_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] net629 _1880_ VPWR
+ VGND sg13g2_and2_1
X_4202_ net788 VGND VPWR _0179_ sap_3_inst.alu.act\[1\] clknet_5_20__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
X_2394_ _1815_ _1690_ _1655_ _1661_ _1639_ VPWR VGND sg13g2_a22oi_1
X_4133_ net779 VGND VPWR _0111_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\]
+ clknet_5_14__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4064_ net783 VGND VPWR _0042_ sap_3_inst.out\[0\] clknet_5_16__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_49_591 VPWR VGND sg13g2_decap_8
X_3015_ net564 _0326_ _1953_ _0568_ VPWR VGND _0567_ sg13g2_nand4_1
XFILLER_25_926 VPWR VGND sg13g2_decap_8
XFILLER_37_786 VPWR VGND sg13g2_decap_8
XFILLER_24_414 VPWR VGND sg13g2_decap_8
XFILLER_40_907 VPWR VGND sg13g2_decap_8
XFILLER_12_609 VPWR VGND sg13g2_decap_8
XFILLER_33_970 VPWR VGND sg13g2_decap_8
X_3917_ _1354_ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[4\] _1312_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_653 VPWR VGND sg13g2_decap_8
X_3848_ net66 _0156_ _1290_ VPWR VGND sg13g2_nor2_1
X_3779_ _1020_ _0997_ _1244_ VPWR VGND sg13g2_xor2_1
XFILLER_47_528 VPWR VGND sg13g2_decap_8
XFILLER_28_764 VPWR VGND sg13g2_decap_8
XFILLER_43_712 VPWR VGND sg13g2_decap_8
XFILLER_15_414 VPWR VGND sg13g2_fill_2
XFILLER_31_918 VPWR VGND sg13g2_decap_8
XFILLER_43_789 VPWR VGND sg13g2_decap_8
XFILLER_24_981 VPWR VGND sg13g2_decap_8
XFILLER_11_620 VPWR VGND sg13g2_decap_8
XFILLER_10_174 VPWR VGND sg13g2_fill_1
XFILLER_7_657 VPWR VGND sg13g2_decap_8
XFILLER_11_697 VPWR VGND sg13g2_decap_8
XFILLER_3_885 VPWR VGND sg13g2_decap_8
XFILLER_33_8 VPWR VGND sg13g2_fill_1
XFILLER_19_775 VPWR VGND sg13g2_decap_8
XFILLER_22_918 VPWR VGND sg13g2_decap_8
XFILLER_34_767 VPWR VGND sg13g2_decap_8
XFILLER_18_1020 VPWR VGND sg13g2_decap_8
XFILLER_30_962 VPWR VGND sg13g2_decap_8
X_3702_ net580 VPWR _1192_ VGND net647 _1001_ sg13g2_o21ai_1
X_3633_ net550 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[7\] _1137_ _0098_
+ VPWR VGND sg13g2_a21o_1
X_3564_ net590 _0861_ _1083_ _1084_ VPWR VGND sg13g2_nor3_1
X_2515_ _1923_ VPWR _1928_ VGND net690 _1927_ sg13g2_o21ai_1
X_3495_ _0858_ _1023_ _1024_ VPWR VGND sg13g2_nor2b_2
X_2446_ _1865_ _1862_ _1863_ _1864_ VPWR VGND sg13g2_and3_1
XFILLER_25_1024 VPWR VGND sg13g2_decap_4
X_2377_ net662 _1762_ _1793_ _1798_ VPWR VGND sg13g2_nor3_2
X_4116_ net793 VGND VPWR _0094_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[3\]
+ clknet_5_27__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_29_517 VPWR VGND sg13g2_decap_8
X_4047_ net786 VGND VPWR _0029_ sap_3_inst.alu.flags\[3\] net39 sg13g2_dfrbpq_1
XFILLER_25_723 VPWR VGND sg13g2_decap_8
XFILLER_37_583 VPWR VGND sg13g2_decap_8
XFILLER_40_704 VPWR VGND sg13g2_decap_8
XFILLER_13_929 VPWR VGND sg13g2_decap_8
XFILLER_21_940 VPWR VGND sg13g2_decap_8
XFILLER_4_649 VPWR VGND sg13g2_decap_8
XFILLER_3_115 VPWR VGND sg13g2_decap_8
XFILLER_0_855 VPWR VGND sg13g2_decap_8
XFILLER_48_815 VPWR VGND sg13g2_decap_8
XFILLER_28_561 VPWR VGND sg13g2_decap_8
XFILLER_16_767 VPWR VGND sg13g2_decap_8
XFILLER_43_586 VPWR VGND sg13g2_decap_8
XFILLER_31_715 VPWR VGND sg13g2_decap_8
XFILLER_11_450 VPWR VGND sg13g2_fill_2
XFILLER_12_973 VPWR VGND sg13g2_decap_8
XFILLER_8_944 VPWR VGND sg13g2_decap_8
XFILLER_3_682 VPWR VGND sg13g2_decap_8
X_2300_ _1541_ _1719_ _1720_ _1721_ VPWR VGND sg13g2_nor3_1
X_3280_ _0816_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] net641 VPWR
+ VGND sg13g2_nand2_1
X_2231_ _1652_ _1579_ _1651_ VPWR VGND sg13g2_nand2_1
X_2162_ _1567_ _1574_ _1583_ VPWR VGND sg13g2_nor2_2
XFILLER_39_859 VPWR VGND sg13g2_decap_8
X_2093_ net736 net724 _1511_ _1514_ VPWR VGND sg13g2_nor3_2
XFILLER_47_892 VPWR VGND sg13g2_decap_8
X_2076__1 VPWR net35 clknet_1_0__leaf_clk_div_out VGND sg13g2_inv_1
XFILLER_19_572 VPWR VGND sg13g2_decap_8
XFILLER_0_73 VPWR VGND sg13g2_fill_1
XFILLER_22_715 VPWR VGND sg13g2_decap_8
XFILLER_34_564 VPWR VGND sg13g2_decap_8
X_2995_ VGND VPWR net543 _0552_ _0557_ net670 sg13g2_a21oi_1
X_3616_ net551 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] _1127_ _0091_
+ VPWR VGND sg13g2_a21o_1
X_3547_ _1069_ _0844_ _0855_ VPWR VGND sg13g2_nand2_1
X_3478_ net586 VPWR _1008_ VGND net615 _1007_ sg13g2_o21ai_1
X_2429_ _1850_ net619 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[7\] net631
+ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_45_807 VPWR VGND sg13g2_decap_8
XFILLER_44_317 VPWR VGND sg13g2_fill_2
XFILLER_25_520 VPWR VGND sg13g2_decap_8
XFILLER_44_68 VPWR VGND sg13g2_fill_2
XFILLER_40_501 VPWR VGND sg13g2_decap_8
XFILLER_13_726 VPWR VGND sg13g2_decap_8
XFILLER_25_597 VPWR VGND sg13g2_decap_8
XFILLER_40_578 VPWR VGND sg13g2_decap_8
XFILLER_9_719 VPWR VGND sg13g2_decap_8
XFILLER_5_936 VPWR VGND sg13g2_decap_8
XFILLER_4_402 VPWR VGND sg13g2_fill_1
XFILLER_48_612 VPWR VGND sg13g2_decap_8
XFILLER_0_652 VPWR VGND sg13g2_decap_8
XFILLER_48_689 VPWR VGND sg13g2_decap_8
XFILLER_29_881 VPWR VGND sg13g2_decap_8
XFILLER_36_829 VPWR VGND sg13g2_decap_8
XFILLER_16_564 VPWR VGND sg13g2_decap_8
XFILLER_31_512 VPWR VGND sg13g2_decap_8
XFILLER_8_741 VPWR VGND sg13g2_decap_8
X_2780_ _0342_ _0346_ _0348_ _0349_ VPWR VGND sg13g2_nor3_1
XFILLER_12_770 VPWR VGND sg13g2_decap_8
XFILLER_31_589 VPWR VGND sg13g2_decap_8
X_3401_ _0927_ _0929_ _0933_ _0934_ VPWR VGND sg13g2_nor3_1
X_3332_ _0867_ net611 _0865_ _0866_ VPWR VGND sg13g2_and3_1
Xfanout709 _1565_ net709 VPWR VGND sg13g2_buf_8
X_3263_ _0799_ net645 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[2\] net648
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2214_ _1635_ sap_3_inst.controller.stage\[2\] net719 net718 VPWR VGND sg13g2_and3_2
XFILLER_22_1016 VPWR VGND sg13g2_decap_8
X_3194_ _0730_ net649 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[0\] net653
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_15_0 VPWR VGND sg13g2_fill_2
X_2145_ _1521_ net709 _1566_ VPWR VGND sg13g2_nor2_1
XFILLER_22_1027 VPWR VGND sg13g2_fill_2
XFILLER_39_656 VPWR VGND sg13g2_decap_8
XFILLER_35_884 VPWR VGND sg13g2_decap_8
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_22_512 VPWR VGND sg13g2_decap_8
X_2978_ sap_3_inst.alu.tmp\[7\] net743 _0540_ VPWR VGND sg13g2_xor2_1
XFILLER_22_589 VPWR VGND sg13g2_decap_8
XFILLER_2_917 VPWR VGND sg13g2_decap_8
XFILLER_49_409 VPWR VGND sg13g2_decap_8
XFILLER_29_100 VPWR VGND sg13g2_fill_1
XFILLER_45_604 VPWR VGND sg13g2_decap_8
XFILLER_26_884 VPWR VGND sg13g2_decap_8
XFILLER_38_1012 VPWR VGND sg13g2_decap_8
XFILLER_41_843 VPWR VGND sg13g2_decap_8
XFILLER_13_523 VPWR VGND sg13g2_decap_8
XFILLER_25_394 VPWR VGND sg13g2_decap_8
XFILLER_9_516 VPWR VGND sg13g2_decap_8
XFILLER_5_733 VPWR VGND sg13g2_decap_8
XFILLER_4_210 VPWR VGND sg13g2_fill_1
XFILLER_1_961 VPWR VGND sg13g2_decap_8
XFILLER_49_976 VPWR VGND sg13g2_decap_8
XFILLER_48_486 VPWR VGND sg13g2_decap_8
XFILLER_36_626 VPWR VGND sg13g2_decap_8
X_3950_ _1280_ net52 _1383_ _0169_ VPWR VGND sg13g2_a21o_1
X_2901_ _0465_ VPWR _0466_ VGND _0444_ _0445_ sg13g2_o21ai_1
XFILLER_32_854 VPWR VGND sg13g2_decap_8
X_3881_ _1319_ _1320_ _1318_ _1322_ VPWR VGND _1321_ sg13g2_nand4_1
X_2832_ _0399_ net756 net672 VPWR VGND sg13g2_nand2_1
XFILLER_31_386 VPWR VGND sg13g2_fill_1
X_2763_ VPWR _0332_ net543 VGND sg13g2_inv_1
X_2694_ net716 _1635_ _0283_ VPWR VGND sg13g2_nor2_1
XFILLER_6_83 VPWR VGND sg13g2_decap_8
X_3315_ _0851_ _0788_ _0849_ VPWR VGND sg13g2_nand2_1
X_3246_ _0782_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[3\] net641 VPWR
+ VGND sg13g2_nand2_1
X_3177_ _0694_ _0711_ _0691_ _0713_ VPWR VGND sg13g2_nand3_1
X_2128_ net739 _1436_ _1521_ _1549_ VPWR VGND sg13g2_nor3_2
XFILLER_27_648 VPWR VGND sg13g2_decap_8
XFILLER_42_629 VPWR VGND sg13g2_decap_8
X_2059_ VPWR _1482_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_26_147 VPWR VGND sg13g2_fill_2
XFILLER_23_843 VPWR VGND sg13g2_decap_8
XFILLER_35_681 VPWR VGND sg13g2_decap_8
XFILLER_22_375 VPWR VGND sg13g2_decap_4
XFILLER_10_559 VPWR VGND sg13g2_decap_8
XFILLER_6_519 VPWR VGND sg13g2_decap_8
XFILLER_2_714 VPWR VGND sg13g2_decap_8
XFILLER_46_913 VPWR VGND sg13g2_decap_8
XFILLER_45_401 VPWR VGND sg13g2_decap_8
XFILLER_45_478 VPWR VGND sg13g2_decap_8
XFILLER_14_810 VPWR VGND sg13g2_decap_8
XFILLER_26_681 VPWR VGND sg13g2_decap_8
XFILLER_41_640 VPWR VGND sg13g2_decap_8
XFILLER_14_887 VPWR VGND sg13g2_decap_8
XFILLER_12_1015 VPWR VGND sg13g2_decap_8
XFILLER_5_530 VPWR VGND sg13g2_decap_8
XFILLER_31_91 VPWR VGND sg13g2_fill_1
X_3100_ _1553_ net684 net731 _0636_ VPWR VGND _1716_ sg13g2_nand4_1
X_4080_ net791 VGND VPWR _0058_ sap_3_inst.alu.tmp\[7\] clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_49_773 VPWR VGND sg13g2_decap_8
X_3031_ _0562_ sap_3_inst.alu.carry _0583_ _0050_ VPWR VGND sg13g2_a21o_1
XFILLER_37_968 VPWR VGND sg13g2_decap_8
XFILLER_32_651 VPWR VGND sg13g2_decap_8
X_3933_ VGND VPWR sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[6\] _1311_
+ _1368_ net763 sg13g2_a21oi_1
X_3864_ net768 _1304_ _1305_ VPWR VGND sg13g2_nor2_2
X_2815_ _0382_ net755 sap_3_inst.alu.tmp\[2\] VPWR VGND sg13g2_xnor2_1
XFILLER_20_835 VPWR VGND sg13g2_decap_8
X_3795_ VGND VPWR _1470_ net599 _0143_ _1254_ sg13g2_a21oi_1
XFILLER_9_880 VPWR VGND sg13g2_decap_8
X_2746_ net618 _1950_ _1946_ _0315_ VPWR VGND sg13g2_nand3_1
X_2677_ _1599_ VPWR _0269_ VGND net696 _1626_ sg13g2_o21ai_1
X_3229_ _0760_ _0761_ _0762_ _0763_ _0765_ VPWR VGND sg13g2_and4_1
XFILLER_27_401 VPWR VGND sg13g2_decap_4
XFILLER_28_946 VPWR VGND sg13g2_decap_8
XFILLER_27_445 VPWR VGND sg13g2_decap_8
XFILLER_42_426 VPWR VGND sg13g2_fill_2
XFILLER_14_117 VPWR VGND sg13g2_fill_2
XFILLER_36_990 VPWR VGND sg13g2_decap_8
XFILLER_14_139 VPWR VGND sg13g2_fill_2
XFILLER_23_640 VPWR VGND sg13g2_decap_8
XFILLER_11_802 VPWR VGND sg13g2_decap_8
XFILLER_10_312 VPWR VGND sg13g2_fill_2
XFILLER_7_839 VPWR VGND sg13g2_decap_8
XFILLER_11_879 VPWR VGND sg13g2_decap_8
XFILLER_6_349 VPWR VGND sg13g2_fill_1
Xclkbuf_4_8_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_8_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_2_511 VPWR VGND sg13g2_decap_8
XFILLER_2_588 VPWR VGND sg13g2_decap_8
XFILLER_46_710 VPWR VGND sg13g2_decap_8
XFILLER_19_957 VPWR VGND sg13g2_decap_8
XFILLER_46_787 VPWR VGND sg13g2_decap_8
XFILLER_34_949 VPWR VGND sg13g2_decap_8
XFILLER_33_459 VPWR VGND sg13g2_fill_2
XFILLER_42_993 VPWR VGND sg13g2_decap_8
XFILLER_14_684 VPWR VGND sg13g2_decap_8
XFILLER_9_110 VPWR VGND sg13g2_fill_2
XFILLER_9_165 VPWR VGND sg13g2_fill_1
X_2600_ _0197_ _1946_ _1951_ VPWR VGND sg13g2_nand2_2
X_3580_ VPWR VGND _1096_ _0929_ _1095_ _0933_ _1097_ _1094_ sg13g2_a221oi_1
X_2531_ _1521_ net695 net709 _1944_ VPWR VGND sg13g2_nor3_2
XFILLER_6_883 VPWR VGND sg13g2_decap_8
X_4201_ net788 VGND VPWR _0178_ sap_3_inst.alu.act\[0\] clknet_5_17__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_2462_ VGND VPWR net675 _1878_ _0032_ _1879_ sg13g2_a21oi_1
X_2393_ _1550_ _1559_ _1814_ VPWR VGND sg13g2_nor2_2
X_4132_ net795 VGND VPWR _0110_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\]
+ clknet_5_28__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_49_570 VPWR VGND sg13g2_decap_8
X_4063_ net791 VGND VPWR _0041_ sap_3_inst.alu.acc\[7\] clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
X_3014_ _1944_ VPWR _0567_ VGND net732 _1943_ sg13g2_o21ai_1
XFILLER_25_905 VPWR VGND sg13g2_decap_8
XFILLER_37_765 VPWR VGND sg13g2_decap_8
X_3916_ _1353_ net721 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[4\] _1308_
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[4\] VPWR VGND sg13g2_a22oi_1
Xclkbuf_5_7__f_sap_3_inst.alu.clk_regs clknet_4_3_0_sap_3_inst.alu.clk_regs clknet_5_7__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_20_632 VPWR VGND sg13g2_decap_8
X_3847_ regFile_serial_start net75 _0155_ _0160_ VPWR VGND sg13g2_a21o_1
X_3778_ _0137_ _1114_ _1243_ net601 _1483_ VPWR VGND sg13g2_a22oi_1
X_2729_ _1504_ net713 net733 _0298_ VPWR VGND sg13g2_nand3_1
XFILLER_47_507 VPWR VGND sg13g2_decap_8
XFILLER_47_46 VPWR VGND sg13g2_fill_1
XFILLER_28_743 VPWR VGND sg13g2_decap_8
XFILLER_16_949 VPWR VGND sg13g2_decap_8
XFILLER_43_768 VPWR VGND sg13g2_decap_8
XFILLER_24_960 VPWR VGND sg13g2_decap_8
XFILLER_10_120 VPWR VGND sg13g2_fill_2
XFILLER_11_676 VPWR VGND sg13g2_decap_8
XFILLER_7_636 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_fill_2
XFILLER_3_864 VPWR VGND sg13g2_decap_8
XFILLER_38_529 VPWR VGND sg13g2_decap_8
XFILLER_18_220 VPWR VGND sg13g2_fill_2
XFILLER_19_754 VPWR VGND sg13g2_decap_8
XFILLER_46_584 VPWR VGND sg13g2_decap_8
XFILLER_18_264 VPWR VGND sg13g2_fill_1
XFILLER_34_746 VPWR VGND sg13g2_decap_8
Xclkbuf_5_14__f_sap_3_inst.alu.clk_regs clknet_4_7_0_sap_3_inst.alu.clk_regs clknet_5_14__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_42_790 VPWR VGND sg13g2_decap_8
XFILLER_30_941 VPWR VGND sg13g2_decap_8
X_3701_ _1191_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] _1181_ VPWR
+ VGND sg13g2_nand2_1
X_3632_ _1025_ _1075_ net550 _1137_ VPWR VGND sg13g2_nor3_1
XFILLER_6_680 VPWR VGND sg13g2_decap_8
X_3563_ _0846_ _1082_ _1083_ VPWR VGND sg13g2_nor2_1
XFILLER_45_0 VPWR VGND sg13g2_fill_1
X_2514_ VGND VPWR net688 _1568_ _1927_ _1925_ sg13g2_a21oi_1
X_3494_ net553 VPWR _1023_ VGND net559 _0855_ sg13g2_o21ai_1
X_2445_ _1864_ net621 sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] net627
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_25_1003 VPWR VGND sg13g2_decap_8
X_2376_ _1797_ net662 _1762_ _1772_ VPWR VGND sg13g2_and3_2
X_4115_ net795 VGND VPWR _0093_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[2\]
+ clknet_5_27__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4046_ net786 VGND VPWR _0028_ sap_3_inst.alu.flags\[2\] net38 sg13g2_dfrbpq_1
XFILLER_25_702 VPWR VGND sg13g2_decap_8
XFILLER_37_562 VPWR VGND sg13g2_decap_8
XFILLER_13_908 VPWR VGND sg13g2_decap_8
XFILLER_24_234 VPWR VGND sg13g2_fill_1
XFILLER_25_779 VPWR VGND sg13g2_decap_8
XFILLER_21_996 VPWR VGND sg13g2_decap_8
XFILLER_4_628 VPWR VGND sg13g2_decap_8
XFILLER_0_834 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_28_540 VPWR VGND sg13g2_decap_8
XFILLER_16_746 VPWR VGND sg13g2_decap_8
XFILLER_43_565 VPWR VGND sg13g2_decap_8
XFILLER_8_923 VPWR VGND sg13g2_decap_8
XFILLER_12_952 VPWR VGND sg13g2_decap_8
XFILLER_48_1025 VPWR VGND sg13g2_decap_4
XFILLER_3_661 VPWR VGND sg13g2_decap_8
X_2230_ _1651_ _1633_ net714 net704 net711 VPWR VGND sg13g2_a22oi_1
X_2161_ _1582_ _1535_ net710 VPWR VGND sg13g2_nand2_2
XFILLER_39_838 VPWR VGND sg13g2_decap_8
X_2092_ _1513_ _1508_ _1510_ VPWR VGND sg13g2_nand2_1
XFILLER_19_551 VPWR VGND sg13g2_decap_8
XFILLER_38_359 VPWR VGND sg13g2_fill_1
XFILLER_47_871 VPWR VGND sg13g2_decap_8
XFILLER_0_1016 VPWR VGND sg13g2_decap_8
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_381 VPWR VGND sg13g2_decap_8
XFILLER_0_96 VPWR VGND sg13g2_decap_8
XFILLER_34_543 VPWR VGND sg13g2_decap_8
X_2994_ net544 _0537_ _0550_ _0555_ _0556_ VPWR VGND sg13g2_or4_1
X_3615_ _1040_ _1041_ net550 _1127_ VPWR VGND sg13g2_nor3_1
X_3546_ _1068_ net547 _1067_ VPWR VGND sg13g2_nand2_2
X_3477_ _0824_ _0757_ _1007_ VPWR VGND sg13g2_xor2_1
X_2428_ _1849_ _1829_ _1848_ VPWR VGND sg13g2_nand2_1
X_2359_ _1626_ VPWR _1780_ VGND _1596_ _1599_ sg13g2_o21ai_1
XFILLER_38_893 VPWR VGND sg13g2_decap_8
XFILLER_13_705 VPWR VGND sg13g2_decap_8
XFILLER_25_576 VPWR VGND sg13g2_decap_8
XFILLER_40_557 VPWR VGND sg13g2_decap_8
XFILLER_5_915 VPWR VGND sg13g2_decap_8
XFILLER_21_793 VPWR VGND sg13g2_decap_8
XFILLER_4_447 VPWR VGND sg13g2_fill_2
XFILLER_0_631 VPWR VGND sg13g2_decap_8
XFILLER_48_668 VPWR VGND sg13g2_decap_8
XFILLER_36_808 VPWR VGND sg13g2_decap_8
XFILLER_29_860 VPWR VGND sg13g2_decap_8
XFILLER_16_543 VPWR VGND sg13g2_decap_8
XFILLER_44_885 VPWR VGND sg13g2_decap_8
XFILLER_31_568 VPWR VGND sg13g2_decap_8
XFILLER_8_720 VPWR VGND sg13g2_decap_8
XFILLER_8_797 VPWR VGND sg13g2_decap_8
X_3400_ VGND VPWR net583 _0933_ _0932_ _0931_ sg13g2_a21oi_2
X_3331_ _0866_ net650 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[1\] net653
+ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_4_992 VPWR VGND sg13g2_decap_8
X_3262_ _0798_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[2\] net656 VPWR
+ VGND sg13g2_nand2_1
X_2213_ _1634_ net717 net716 VPWR VGND sg13g2_nand2_1
X_3193_ _0710_ _0728_ _0729_ VPWR VGND sg13g2_and2_1
XFILLER_39_635 VPWR VGND sg13g2_decap_8
X_2144_ _1565_ net737 _1563_ VPWR VGND sg13g2_nand2_2
X_2075_ VPWR _1498_ net768 VGND sg13g2_inv_1
XFILLER_19_392 VPWR VGND sg13g2_fill_1
XFILLER_35_863 VPWR VGND sg13g2_decap_8
X_4035__13 VPWR net47 clknet_leaf_1_sap_3_inst.alu.clk VGND sg13g2_inv_1
XFILLER_34_373 VPWR VGND sg13g2_fill_2
XFILLER_22_568 VPWR VGND sg13g2_decap_8
X_2977_ net743 sap_3_inst.alu.tmp\[7\] _0539_ VPWR VGND sg13g2_and2_1
X_3529_ _1054_ _1975_ _1053_ VPWR VGND sg13g2_nand2_1
XFILLER_38_690 VPWR VGND sg13g2_decap_8
XFILLER_26_863 VPWR VGND sg13g2_decap_8
XFILLER_41_822 VPWR VGND sg13g2_decap_8
XFILLER_13_502 VPWR VGND sg13g2_decap_8
XFILLER_41_899 VPWR VGND sg13g2_decap_8
XFILLER_13_579 VPWR VGND sg13g2_decap_8
XFILLER_21_590 VPWR VGND sg13g2_decap_8
XFILLER_5_712 VPWR VGND sg13g2_decap_8
XFILLER_5_789 VPWR VGND sg13g2_decap_8
XFILLER_45_1017 VPWR VGND sg13g2_decap_8
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_940 VPWR VGND sg13g2_decap_8
XFILLER_49_955 VPWR VGND sg13g2_decap_8
XFILLER_48_465 VPWR VGND sg13g2_decap_8
XFILLER_36_605 VPWR VGND sg13g2_decap_8
XFILLER_44_682 VPWR VGND sg13g2_decap_8
X_2900_ net543 _0454_ _0462_ _0464_ _0465_ VPWR VGND sg13g2_nor4_1
XFILLER_17_885 VPWR VGND sg13g2_decap_8
XFILLER_32_833 VPWR VGND sg13g2_decap_8
X_3880_ _1321_ net761 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\] _1312_
+ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2831_ VPWR VGND _0333_ _0397_ _0383_ net753 _0398_ net572 sg13g2_a221oi_1
X_2762_ _0199_ _0329_ net563 _0331_ VPWR VGND sg13g2_nor3_1
XFILLER_8_594 VPWR VGND sg13g2_decap_8
X_2693_ _1635_ _1744_ _0282_ _0004_ VPWR VGND sg13g2_nor3_1
X_3314_ VGND VPWR _0850_ _0820_ _0808_ sg13g2_or2_1
X_3245_ _0781_ _0779_ _0780_ VPWR VGND sg13g2_nand2_1
X_3176_ _0712_ _0691_ _0694_ _0711_ VPWR VGND sg13g2_and3_2
XFILLER_27_627 VPWR VGND sg13g2_decap_8
X_2127_ _1548_ _1547_ _1541_ VPWR VGND sg13g2_nand2b_1
XFILLER_42_608 VPWR VGND sg13g2_decap_8
XFILLER_35_660 VPWR VGND sg13g2_decap_8
X_2058_ VPWR _1481_ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_41_107 VPWR VGND sg13g2_fill_1
XFILLER_23_822 VPWR VGND sg13g2_decap_8
XFILLER_34_192 VPWR VGND sg13g2_fill_1
XFILLER_23_899 VPWR VGND sg13g2_decap_8
XFILLER_10_538 VPWR VGND sg13g2_decap_8
XFILLER_9_6 VPWR VGND sg13g2_fill_1
XFILLER_1_214 VPWR VGND sg13g2_fill_2
XFILLER_1_258 VPWR VGND sg13g2_fill_2
XFILLER_46_969 VPWR VGND sg13g2_decap_8
XFILLER_18_649 VPWR VGND sg13g2_decap_8
XFILLER_45_457 VPWR VGND sg13g2_decap_8
XFILLER_26_660 VPWR VGND sg13g2_decap_8
XFILLER_32_118 VPWR VGND sg13g2_fill_1
XFILLER_14_866 VPWR VGND sg13g2_decap_8
XFILLER_41_696 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_5_586 VPWR VGND sg13g2_decap_8
XFILLER_49_752 VPWR VGND sg13g2_decap_8
X_3030_ _0562_ _0581_ _0582_ _0583_ VPWR VGND sg13g2_nor3_1
XFILLER_37_947 VPWR VGND sg13g2_decap_8
XFILLER_17_682 VPWR VGND sg13g2_decap_8
XFILLER_32_630 VPWR VGND sg13g2_decap_8
X_3932_ net764 net55 _1367_ _0167_ VPWR VGND sg13g2_a21o_1
X_3863_ VGND VPWR _1304_ _1303_ _1497_ sg13g2_or2_1
XFILLER_20_814 VPWR VGND sg13g2_decap_8
X_2814_ net545 net616 _0381_ VPWR VGND sg13g2_nor2b_1
X_3794_ net598 _0952_ _1188_ _1254_ VPWR VGND sg13g2_nor3_1
XFILLER_8_391 VPWR VGND sg13g2_fill_2
X_2745_ _1822_ VPWR _0314_ VGND _0312_ _0313_ sg13g2_o21ai_1
X_2676_ _1587_ VPWR _0268_ VGND net696 _1646_ sg13g2_o21ai_1
XFILLER_28_1023 VPWR VGND sg13g2_decap_4
X_3228_ _0764_ net587 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] net613
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_28_925 VPWR VGND sg13g2_decap_8
X_3159_ _0695_ _0691_ _0694_ VPWR VGND sg13g2_nand2_2
XFILLER_15_619 VPWR VGND sg13g2_decap_8
XFILLER_11_858 VPWR VGND sg13g2_decap_8
XFILLER_23_696 VPWR VGND sg13g2_decap_8
XFILLER_7_818 VPWR VGND sg13g2_decap_8
XFILLER_2_567 VPWR VGND sg13g2_decap_8
XFILLER_18_424 VPWR VGND sg13g2_fill_1
XFILLER_19_936 VPWR VGND sg13g2_decap_8
XFILLER_46_766 VPWR VGND sg13g2_decap_8
XFILLER_27_991 VPWR VGND sg13g2_decap_8
XFILLER_34_928 VPWR VGND sg13g2_decap_8
XFILLER_42_972 VPWR VGND sg13g2_decap_8
XFILLER_14_663 VPWR VGND sg13g2_decap_8
XFILLER_41_493 VPWR VGND sg13g2_decap_8
XFILLER_9_188 VPWR VGND sg13g2_fill_1
XFILLER_6_862 VPWR VGND sg13g2_decap_8
X_2530_ _1941_ _1942_ _1943_ VPWR VGND sg13g2_and2_1
X_2461_ sap_3_inst.alu.flags\[6\] net675 _1879_ VPWR VGND sg13g2_nor2_1
X_4200_ net785 VGND VPWR net35 clk_div_out clknet_3_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_3_30 VPWR VGND sg13g2_fill_2
X_2392_ net709 _1812_ _1813_ VPWR VGND sg13g2_nor2_1
X_4131_ net786 VGND VPWR _0109_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[2\]
+ clknet_5_24__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4062_ net791 VGND VPWR _0040_ sap_3_inst.alu.acc\[6\] clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_3_1025 VPWR VGND sg13g2_decap_4
X_3013_ VGND VPWR _0543_ _0565_ _0566_ net564 sg13g2_a21oi_1
XFILLER_37_744 VPWR VGND sg13g2_decap_8
XFILLER_24_449 VPWR VGND sg13g2_decap_8
X_3915_ _1352_ net761 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[4\] _1305_
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_20_611 VPWR VGND sg13g2_decap_8
X_3846_ _0159_ _1287_ _1288_ VPWR VGND sg13g2_nand2_1
XFILLER_20_688 VPWR VGND sg13g2_decap_8
X_3777_ net15 net599 _1242_ _1243_ VPWR VGND sg13g2_nor3_1
X_2728_ net60 sap_3_inst.out\[7\] _0186_ _0025_ VPWR VGND sg13g2_mux2_1
X_2659_ sap_3_inst.alu.act\[5\] sap_3_inst.alu.act\[4\] sap_3_inst.alu.act\[7\] sap_3_inst.alu.act\[6\]
+ _0253_ VPWR VGND sg13g2_nor4_1
XFILLER_28_722 VPWR VGND sg13g2_decap_8
XFILLER_16_928 VPWR VGND sg13g2_decap_8
XFILLER_28_799 VPWR VGND sg13g2_decap_8
XFILLER_43_747 VPWR VGND sg13g2_decap_8
XFILLER_23_493 VPWR VGND sg13g2_decap_8
XFILLER_7_615 VPWR VGND sg13g2_decap_8
XFILLER_11_655 VPWR VGND sg13g2_decap_8
XFILLER_10_154 VPWR VGND sg13g2_fill_2
XFILLER_3_843 VPWR VGND sg13g2_decap_8
XFILLER_38_508 VPWR VGND sg13g2_decap_8
Xfanout690 _1552_ net690 VPWR VGND sg13g2_buf_1
XFILLER_19_733 VPWR VGND sg13g2_decap_8
XFILLER_46_563 VPWR VGND sg13g2_decap_8
XFILLER_34_725 VPWR VGND sg13g2_decap_8
X_3700_ VGND VPWR _1182_ _1190_ _0112_ _1189_ sg13g2_a21oi_1
XFILLER_14_460 VPWR VGND sg13g2_fill_1
XFILLER_15_983 VPWR VGND sg13g2_decap_8
XFILLER_30_920 VPWR VGND sg13g2_decap_8
XFILLER_30_997 VPWR VGND sg13g2_decap_8
X_3631_ VGND VPWR _1487_ net551 _0097_ _1136_ sg13g2_a21oi_1
X_3562_ _1082_ _1081_ _0828_ _1080_ _1079_ VPWR VGND sg13g2_a22oi_1
X_2513_ VPWR _1926_ _1925_ VGND sg13g2_inv_1
X_3493_ _1022_ net612 _1021_ VPWR VGND sg13g2_nand2b_1
X_2444_ _1863_ net625 sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] net629
+ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2375_ net662 _1761_ _1791_ _1796_ VPWR VGND sg13g2_nor3_2
XFILLER_38_0 VPWR VGND sg13g2_fill_1
X_4114_ net793 VGND VPWR _0092_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[1\]
+ clknet_5_25__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4045_ net783 VGND VPWR _0027_ sap_3_inst.alu.flags\[1\] net37 sg13g2_dfrbpq_1
XFILLER_37_541 VPWR VGND sg13g2_decap_8
XFILLER_25_758 VPWR VGND sg13g2_decap_8
XFILLER_40_739 VPWR VGND sg13g2_decap_8
XFILLER_21_975 VPWR VGND sg13g2_decap_8
XFILLER_32_1008 VPWR VGND sg13g2_decap_8
X_3829_ net578 _1173_ _1277_ _1278_ VPWR VGND sg13g2_nor3_1
XFILLER_20_485 VPWR VGND sg13g2_decap_8
XFILLER_4_607 VPWR VGND sg13g2_decap_8
XFILLER_0_813 VPWR VGND sg13g2_decap_8
XFILLER_16_725 VPWR VGND sg13g2_decap_8
XFILLER_43_544 VPWR VGND sg13g2_decap_8
XFILLER_15_224 VPWR VGND sg13g2_fill_2
XFILLER_28_596 VPWR VGND sg13g2_decap_8
XFILLER_12_931 VPWR VGND sg13g2_decap_8
XFILLER_8_902 VPWR VGND sg13g2_decap_8
XFILLER_8_979 VPWR VGND sg13g2_decap_8
XFILLER_48_1004 VPWR VGND sg13g2_decap_8
XFILLER_3_640 VPWR VGND sg13g2_decap_8
XFILLER_2_172 VPWR VGND sg13g2_fill_1
XFILLER_39_817 VPWR VGND sg13g2_decap_8
X_2160_ _1536_ _1557_ _1581_ VPWR VGND sg13g2_nor2_2
XFILLER_47_850 VPWR VGND sg13g2_decap_8
X_2091_ _1509_ _1511_ _1512_ VPWR VGND sg13g2_nor2_1
XFILLER_19_530 VPWR VGND sg13g2_decap_8
XFILLER_0_64 VPWR VGND sg13g2_decap_8
XFILLER_34_522 VPWR VGND sg13g2_decap_8
X_2993_ _0554_ VPWR _0555_ VGND _2007_ _0544_ sg13g2_o21ai_1
XFILLER_15_780 VPWR VGND sg13g2_decap_8
XFILLER_34_599 VPWR VGND sg13g2_decap_8
XFILLER_9_51 VPWR VGND sg13g2_fill_1
XFILLER_9_40 VPWR VGND sg13g2_fill_2
XFILLER_30_794 VPWR VGND sg13g2_decap_8
X_3614_ net640 _1078_ _1126_ VPWR VGND sg13g2_nor2_2
X_3545_ _1067_ net586 _1007_ VPWR VGND sg13g2_nand2_1
X_3476_ _1006_ _0971_ _0994_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_1020 VPWR VGND sg13g2_decap_8
X_2427_ _1848_ net8 _1847_ VPWR VGND sg13g2_nand2_1
X_2358_ _1685_ _1686_ _1777_ _1778_ _1779_ VPWR VGND sg13g2_and4_1
X_2289_ VGND VPWR _1707_ _1709_ _1710_ _1629_ sg13g2_a21oi_1
XFILLER_38_872 VPWR VGND sg13g2_decap_8
XFILLER_25_555 VPWR VGND sg13g2_decap_8
XFILLER_40_536 VPWR VGND sg13g2_decap_8
XFILLER_21_772 VPWR VGND sg13g2_decap_8
XFILLER_0_610 VPWR VGND sg13g2_decap_8
XFILLER_0_687 VPWR VGND sg13g2_decap_8
XFILLER_48_647 VPWR VGND sg13g2_decap_8
XFILLER_16_522 VPWR VGND sg13g2_decap_8
XFILLER_28_371 VPWR VGND sg13g2_decap_4
XFILLER_44_864 VPWR VGND sg13g2_decap_8
XFILLER_16_599 VPWR VGND sg13g2_decap_8
XFILLER_31_547 VPWR VGND sg13g2_decap_8
XFILLER_15_1025 VPWR VGND sg13g2_decap_4
XFILLER_8_776 VPWR VGND sg13g2_decap_8
XFILLER_4_971 VPWR VGND sg13g2_decap_8
X_3330_ _0865_ net645 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[1\] net648
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\] VPWR VGND sg13g2_a22oi_1
X_3261_ _0797_ net560 VPWR VGND sg13g2_inv_2
X_2212_ net717 net716 _1633_ VPWR VGND sg13g2_and2_1
X_3192_ VPWR VGND _0669_ _0655_ _0660_ net702 _0728_ _0652_ sg13g2_a221oi_1
XFILLER_39_614 VPWR VGND sg13g2_decap_8
X_2143_ _1564_ net740 net741 VPWR VGND sg13g2_nand2_1
XFILLER_27_809 VPWR VGND sg13g2_decap_8
X_2074_ net82 _1497_ VPWR VGND sg13g2_inv_4
XFILLER_35_842 VPWR VGND sg13g2_decap_8
XFILLER_22_547 VPWR VGND sg13g2_decap_8
X_2976_ VGND VPWR _0538_ sap_3_inst.alu.tmp\[7\] net743 sg13g2_or2_1
XFILLER_30_591 VPWR VGND sg13g2_decap_8
X_3528_ _0929_ _1052_ _1053_ VPWR VGND sg13g2_nor2_1
X_3459_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[6\] _0988_
+ net588 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] _0989_ net593 sg13g2_a221oi_1
XFILLER_45_639 VPWR VGND sg13g2_decap_8
XFILLER_26_842 VPWR VGND sg13g2_decap_8
XFILLER_41_801 VPWR VGND sg13g2_decap_8
XFILLER_13_558 VPWR VGND sg13g2_decap_8
XFILLER_41_878 VPWR VGND sg13g2_decap_8
XFILLER_5_768 VPWR VGND sg13g2_decap_8
XFILLER_49_934 VPWR VGND sg13g2_decap_8
XFILLER_1_996 VPWR VGND sg13g2_decap_8
XFILLER_48_444 VPWR VGND sg13g2_decap_8
XFILLER_0_484 VPWR VGND sg13g2_decap_8
XFILLER_17_864 VPWR VGND sg13g2_decap_8
XFILLER_44_661 VPWR VGND sg13g2_decap_8
XFILLER_32_812 VPWR VGND sg13g2_decap_8
X_2830_ _0397_ net755 sap_3_inst.alu.tmp\[2\] _0340_ VPWR VGND sg13g2_and3_1
XFILLER_32_889 VPWR VGND sg13g2_decap_8
X_2761_ _1946_ _0201_ _0330_ VPWR VGND sg13g2_and2_1
XFILLER_8_573 VPWR VGND sg13g2_decap_8
X_2692_ _1535_ _0282_ _0003_ VPWR VGND sg13g2_nor2_1
X_3313_ _0849_ _0814_ _0819_ _0807_ _0802_ VPWR VGND sg13g2_a22oi_1
X_3244_ _0780_ net645 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[3\] net653
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_1023 VPWR VGND sg13g2_decap_4
X_3175_ _0708_ _0709_ _1830_ _0711_ VPWR VGND sg13g2_nand3_1
XFILLER_27_606 VPWR VGND sg13g2_decap_8
X_2126_ _1547_ net698 _1546_ VPWR VGND sg13g2_nand2_1
XFILLER_39_488 VPWR VGND sg13g2_decap_8
XFILLER_26_149 VPWR VGND sg13g2_fill_1
X_2057_ VPWR _1480_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[6\] VGND
+ sg13g2_inv_1
XFILLER_23_801 VPWR VGND sg13g2_decap_8
XFILLER_10_517 VPWR VGND sg13g2_decap_8
XFILLER_23_878 VPWR VGND sg13g2_decap_8
X_2959_ VPWR VGND net744 _0521_ net572 net748 _0522_ net573 sg13g2_a221oi_1
XFILLER_2_749 VPWR VGND sg13g2_decap_8
XFILLER_46_948 VPWR VGND sg13g2_decap_8
XFILLER_45_436 VPWR VGND sg13g2_decap_8
XFILLER_18_628 VPWR VGND sg13g2_decap_8
XFILLER_13_300 VPWR VGND sg13g2_fill_2
XFILLER_14_845 VPWR VGND sg13g2_decap_8
XFILLER_41_675 VPWR VGND sg13g2_decap_8
XFILLER_5_565 VPWR VGND sg13g2_decap_8
XFILLER_49_731 VPWR VGND sg13g2_decap_8
XFILLER_1_793 VPWR VGND sg13g2_decap_8
XFILLER_37_926 VPWR VGND sg13g2_decap_8
XFILLER_17_661 VPWR VGND sg13g2_decap_8
X_3931_ VPWR VGND _1366_ net765 _1360_ _1475_ _1367_ net763 sg13g2_a221oi_1
XFILLER_16_171 VPWR VGND sg13g2_fill_2
XFILLER_16_193 VPWR VGND sg13g2_fill_2
X_3862_ _1303_ sap_3_inst.reg_file.array_serializer_inst.word_index\[2\] VPWR VGND
+ sap_3_inst.reg_file.array_serializer_inst.word_index\[3\] sg13g2_nand2b_2
X_2813_ net555 net757 _0380_ _0035_ VPWR VGND sg13g2_a21o_1
XFILLER_32_686 VPWR VGND sg13g2_decap_8
X_3793_ VPWR _0142_ _1253_ VGND sg13g2_inv_1
X_2744_ net683 VPWR _0313_ VGND _1551_ _1814_ sg13g2_o21ai_1
X_2675_ _1750_ _0265_ _1659_ _0267_ VPWR VGND _0266_ sg13g2_nand4_1
XFILLER_28_1002 VPWR VGND sg13g2_decap_8
X_3227_ net659 _0719_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[5\] _0763_
+ VPWR VGND sg13g2_nand3_1
XFILLER_28_904 VPWR VGND sg13g2_decap_8
X_3158_ _0694_ _0692_ _0693_ VPWR VGND sg13g2_nand2_2
X_2109_ _1530_ _1499_ _1527_ VPWR VGND sg13g2_nand2_2
XFILLER_43_929 VPWR VGND sg13g2_decap_8
XFILLER_14_108 VPWR VGND sg13g2_fill_2
XFILLER_14_119 VPWR VGND sg13g2_fill_1
X_3089_ VGND VPWR _0625_ _0624_ _0622_ sg13g2_or2_1
XFILLER_23_675 VPWR VGND sg13g2_decap_8
XFILLER_35_1017 VPWR VGND sg13g2_decap_8
XFILLER_35_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_837 VPWR VGND sg13g2_decap_8
XFILLER_2_546 VPWR VGND sg13g2_decap_8
Xclkbuf_5_22__f_sap_3_inst.alu.clk_regs clknet_4_11_0_sap_3_inst.alu.clk_regs clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_19_915 VPWR VGND sg13g2_decap_8
XFILLER_46_745 VPWR VGND sg13g2_decap_8
XFILLER_34_907 VPWR VGND sg13g2_decap_8
XFILLER_27_970 VPWR VGND sg13g2_decap_8
XFILLER_42_951 VPWR VGND sg13g2_decap_8
XFILLER_14_642 VPWR VGND sg13g2_decap_8
XFILLER_41_472 VPWR VGND sg13g2_decap_8
XFILLER_9_123 VPWR VGND sg13g2_fill_2
XFILLER_9_112 VPWR VGND sg13g2_fill_1
XFILLER_10_881 VPWR VGND sg13g2_decap_8
XFILLER_6_841 VPWR VGND sg13g2_decap_8
X_2460_ net23 net547 VPWR VGND sg13g2_inv_2
X_2391_ _1812_ net712 net685 VPWR VGND sg13g2_nand2_1
X_4130_ net773 VGND VPWR _0108_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[1\]
+ clknet_5_7__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_3_64 VPWR VGND sg13g2_decap_8
XFILLER_3_75 VPWR VGND sg13g2_fill_1
XFILLER_1_590 VPWR VGND sg13g2_decap_8
X_4061_ net790 VGND VPWR _0039_ sap_3_inst.alu.acc\[5\] clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_3_1004 VPWR VGND sg13g2_decap_8
X_3012_ _0564_ VPWR _0565_ VGND _0541_ _0563_ sg13g2_o21ai_1
XFILLER_37_723 VPWR VGND sg13g2_decap_8
XFILLER_18_992 VPWR VGND sg13g2_decap_8
XFILLER_24_428 VPWR VGND sg13g2_decap_8
X_3914_ net764 net51 _1351_ _0165_ VPWR VGND sg13g2_a21o_1
XFILLER_32_461 VPWR VGND sg13g2_fill_2
XFILLER_33_984 VPWR VGND sg13g2_decap_8
X_3845_ _1286_ _1289_ _0158_ VPWR VGND sg13g2_nor2_1
XFILLER_20_667 VPWR VGND sg13g2_decap_8
X_3776_ net574 _0997_ _1241_ _1242_ VPWR VGND sg13g2_nor3_1
X_2727_ net56 sap_3_inst.out\[6\] _0186_ _0024_ VPWR VGND sg13g2_mux2_1
X_2658_ sap_3_inst.alu.act\[1\] sap_3_inst.alu.act\[0\] sap_3_inst.alu.act\[3\] sap_3_inst.alu.act\[2\]
+ _0252_ VPWR VGND sg13g2_nor4_1
X_2589_ net760 net757 _1999_ VPWR VGND sg13g2_xor2_1
XFILLER_27_200 VPWR VGND sg13g2_fill_1
XFILLER_28_701 VPWR VGND sg13g2_decap_8
XFILLER_16_907 VPWR VGND sg13g2_decap_8
XFILLER_43_726 VPWR VGND sg13g2_decap_8
XFILLER_28_778 VPWR VGND sg13g2_decap_8
XFILLER_30_409 VPWR VGND sg13g2_decap_4
XFILLER_23_472 VPWR VGND sg13g2_decap_8
XFILLER_24_995 VPWR VGND sg13g2_decap_8
XFILLER_10_133 VPWR VGND sg13g2_fill_2
XFILLER_10_122 VPWR VGND sg13g2_fill_1
XFILLER_11_634 VPWR VGND sg13g2_decap_8
XFILLER_10_166 VPWR VGND sg13g2_fill_2
XFILLER_10_188 VPWR VGND sg13g2_fill_2
XFILLER_12_62 VPWR VGND sg13g2_fill_1
XFILLER_3_822 VPWR VGND sg13g2_decap_8
XFILLER_12_73 VPWR VGND sg13g2_fill_2
XFILLER_3_899 VPWR VGND sg13g2_decap_8
Xfanout680 net681 net680 VPWR VGND sg13g2_buf_8
XFILLER_19_712 VPWR VGND sg13g2_decap_8
Xfanout691 net692 net691 VPWR VGND sg13g2_buf_8
XFILLER_46_542 VPWR VGND sg13g2_decap_8
XFILLER_19_789 VPWR VGND sg13g2_decap_8
XFILLER_34_704 VPWR VGND sg13g2_decap_8
XFILLER_15_962 VPWR VGND sg13g2_decap_8
XFILLER_33_269 VPWR VGND sg13g2_fill_2
X_3630_ _1002_ _1068_ net550 _1136_ VPWR VGND sg13g2_nor3_1
XFILLER_30_976 VPWR VGND sg13g2_decap_8
X_3561_ VGND VPWR net590 net561 _1081_ _0830_ sg13g2_a21oi_1
X_2512_ net728 _1924_ _1925_ VPWR VGND sg13g2_nor2_1
X_3492_ _1021_ _0998_ _1020_ VPWR VGND sg13g2_xnor2_1
X_2443_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\] net639
+ net636 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[6\] _1862_ net677 sg13g2_a221oi_1
X_2374_ _1795_ _1746_ _1762_ _1792_ VPWR VGND sg13g2_and3_2
X_4113_ net796 VGND VPWR _0091_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[0\]
+ clknet_5_31__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
X_4044_ net786 VGND VPWR _0026_ sap_3_inst.alu.flags\[0\] net36 sg13g2_dfrbpq_1
XFILLER_37_520 VPWR VGND sg13g2_decap_8
XFILLER_25_737 VPWR VGND sg13g2_decap_8
XFILLER_37_597 VPWR VGND sg13g2_decap_8
XFILLER_40_718 VPWR VGND sg13g2_decap_8
XFILLER_33_781 VPWR VGND sg13g2_decap_8
XFILLER_21_954 VPWR VGND sg13g2_decap_8
X_3828_ net16 _0687_ _1277_ VPWR VGND sg13g2_nor2b_1
X_3759_ net11 net599 _1228_ _1229_ VPWR VGND sg13g2_nor3_1
XFILLER_3_129 VPWR VGND sg13g2_decap_8
XFILLER_0_869 VPWR VGND sg13g2_decap_8
XFILLER_48_829 VPWR VGND sg13g2_decap_8
XFILLER_47_339 VPWR VGND sg13g2_decap_8
XFILLER_16_704 VPWR VGND sg13g2_decap_8
XFILLER_28_575 VPWR VGND sg13g2_decap_8
XFILLER_43_523 VPWR VGND sg13g2_decap_8
XFILLER_12_910 VPWR VGND sg13g2_decap_8
XFILLER_30_228 VPWR VGND sg13g2_fill_1
XFILLER_31_729 VPWR VGND sg13g2_decap_8
XFILLER_11_420 VPWR VGND sg13g2_fill_2
XFILLER_24_792 VPWR VGND sg13g2_decap_8
XFILLER_12_987 VPWR VGND sg13g2_decap_8
XFILLER_8_958 VPWR VGND sg13g2_decap_8
Xclkbuf_4_1_0_sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs clknet_4_1_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_3_696 VPWR VGND sg13g2_decap_8
Xclkbuf_5_19__f_sap_3_inst.alu.clk_regs clknet_4_9_0_sap_3_inst.alu.clk_regs clknet_5_19__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2090_ _1511_ net727 VPWR VGND net725 sg13g2_nand2b_2
XFILLER_0_43 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_fill_2
XFILLER_34_501 VPWR VGND sg13g2_decap_8
XFILLER_19_586 VPWR VGND sg13g2_decap_8
X_2992_ _0554_ _0324_ _0553_ VPWR VGND sg13g2_nand2_1
XFILLER_22_729 VPWR VGND sg13g2_decap_8
XFILLER_34_578 VPWR VGND sg13g2_decap_8
XFILLER_30_773 VPWR VGND sg13g2_decap_8
X_3613_ _0090_ _1124_ _1125_ net591 _1496_ VPWR VGND sg13g2_a22oi_1
X_3544_ _0080_ _1064_ _1066_ net558 _1478_ VPWR VGND sg13g2_a22oi_1
X_3475_ _0931_ _0945_ _0969_ _0994_ _1005_ VPWR VGND sg13g2_nor4_1
X_2426_ net693 VPWR _1847_ VGND _1831_ _1846_ sg13g2_o21ai_1
X_2357_ _1778_ _1634_ _1656_ net688 _1555_ VPWR VGND sg13g2_a22oi_1
X_2288_ _1606_ _1708_ _1709_ VPWR VGND sg13g2_nor2_1
XFILLER_38_851 VPWR VGND sg13g2_decap_8
XFILLER_25_534 VPWR VGND sg13g2_decap_8
XFILLER_40_515 VPWR VGND sg13g2_decap_8
XFILLER_12_228 VPWR VGND sg13g2_fill_2
XFILLER_21_751 VPWR VGND sg13g2_decap_8
XFILLER_4_449 VPWR VGND sg13g2_fill_1
XFILLER_48_626 VPWR VGND sg13g2_decap_8
XFILLER_0_666 VPWR VGND sg13g2_decap_8
XFILLER_44_843 VPWR VGND sg13g2_decap_8
XFILLER_29_895 VPWR VGND sg13g2_decap_8
XFILLER_16_578 VPWR VGND sg13g2_decap_8
XFILLER_31_526 VPWR VGND sg13g2_decap_8
XFILLER_15_1004 VPWR VGND sg13g2_decap_8
XFILLER_34_93 VPWR VGND sg13g2_fill_2
XFILLER_8_755 VPWR VGND sg13g2_decap_8
XFILLER_11_261 VPWR VGND sg13g2_fill_1
XFILLER_12_784 VPWR VGND sg13g2_decap_8
XFILLER_4_950 VPWR VGND sg13g2_decap_8
XFILLER_3_493 VPWR VGND sg13g2_decap_8
X_3260_ _0792_ _0793_ _0794_ _0795_ _0796_ VPWR VGND sg13g2_and4_1
X_2211_ net680 _1629_ _1630_ _1632_ VPWR VGND sg13g2_or3_1
X_3191_ _0727_ _0672_ _0710_ VPWR VGND sg13g2_nand2_2
X_2142_ net740 net741 _1563_ VPWR VGND sg13g2_and2_1
X_2073_ VPWR _1496_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_35_821 VPWR VGND sg13g2_decap_8
XFILLER_22_526 VPWR VGND sg13g2_decap_8
XFILLER_35_898 VPWR VGND sg13g2_decap_8
X_2975_ VGND VPWR _0534_ _0535_ _0537_ _0536_ sg13g2_a21oi_1
XFILLER_30_570 VPWR VGND sg13g2_decap_8
X_3527_ net583 _0935_ _1052_ VPWR VGND sg13g2_nor2_1
X_3458_ sap_3_inst.reg_file.array_serializer_inst.data\[3\]\[6\] net641 _0988_ VPWR
+ VGND sg13g2_and2_1
X_2409_ VGND VPWR net713 _1675_ _1830_ _1526_ sg13g2_a21oi_1
X_3389_ _0922_ _0797_ _0851_ VPWR VGND sg13g2_nand2b_1
XFILLER_45_618 VPWR VGND sg13g2_decap_8
XFILLER_44_106 VPWR VGND sg13g2_fill_1
XFILLER_26_821 VPWR VGND sg13g2_decap_8
XFILLER_40_301 VPWR VGND sg13g2_fill_2
XFILLER_25_375 VPWR VGND sg13g2_decap_8
XFILLER_26_898 VPWR VGND sg13g2_decap_8
XFILLER_38_1026 VPWR VGND sg13g2_fill_2
XFILLER_41_857 VPWR VGND sg13g2_decap_8
XFILLER_13_537 VPWR VGND sg13g2_decap_8
XFILLER_5_747 VPWR VGND sg13g2_decap_8
XFILLER_49_913 VPWR VGND sg13g2_decap_8
XFILLER_0_463 VPWR VGND sg13g2_decap_8
XFILLER_1_975 VPWR VGND sg13g2_decap_8
XFILLER_48_423 VPWR VGND sg13g2_decap_8
XFILLER_29_60 VPWR VGND sg13g2_fill_1
XFILLER_29_692 VPWR VGND sg13g2_decap_8
XFILLER_44_640 VPWR VGND sg13g2_decap_8
XFILLER_17_843 VPWR VGND sg13g2_decap_8
XFILLER_32_868 VPWR VGND sg13g2_decap_8
X_2760_ _0329_ _0326_ _0328_ VPWR VGND sg13g2_nand2_1
XFILLER_12_581 VPWR VGND sg13g2_decap_8
XFILLER_8_552 VPWR VGND sg13g2_decap_8
X_2691_ net719 _0282_ _0002_ VPWR VGND sg13g2_nor2_1
X_3312_ _0841_ _0846_ _0848_ VPWR VGND sg13g2_nor2_1
XFILLER_6_1002 VPWR VGND sg13g2_decap_8
X_3243_ _0779_ net648 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[3\] net650
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[3\] VPWR VGND sg13g2_a22oi_1
X_3174_ _0710_ _1830_ _0708_ _0709_ VPWR VGND sg13g2_and3_2
XFILLER_39_467 VPWR VGND sg13g2_decap_8
XFILLER_48_990 VPWR VGND sg13g2_decap_8
X_2125_ _1509_ _1543_ _1546_ VPWR VGND sg13g2_nor2_2
X_2056_ _1479_ sap_3_inst.reg_file.array_serializer_inst.data\[0\]\[6\] VPWR VGND
+ sg13g2_inv_2
XFILLER_23_857 VPWR VGND sg13g2_decap_8
XFILLER_35_695 VPWR VGND sg13g2_decap_8
X_2958_ net618 _0197_ _0506_ _0521_ VPWR VGND sg13g2_nor3_1
XFILLER_31_890 VPWR VGND sg13g2_decap_8
X_2889_ _0453_ VPWR _0454_ VGND net750 _0327_ sg13g2_o21ai_1
XFILLER_2_728 VPWR VGND sg13g2_decap_8
XFILLER_46_927 VPWR VGND sg13g2_decap_8
XFILLER_18_607 VPWR VGND sg13g2_decap_8
XFILLER_45_415 VPWR VGND sg13g2_decap_8
XFILLER_14_824 VPWR VGND sg13g2_decap_8
XFILLER_26_695 VPWR VGND sg13g2_decap_8
XFILLER_41_654 VPWR VGND sg13g2_decap_8
XFILLER_22_890 VPWR VGND sg13g2_decap_8
XFILLER_5_544 VPWR VGND sg13g2_decap_8
XFILLER_1_772 VPWR VGND sg13g2_decap_8
XFILLER_49_710 VPWR VGND sg13g2_decap_8
XFILLER_0_282 VPWR VGND sg13g2_fill_2
XFILLER_37_905 VPWR VGND sg13g2_decap_8
XFILLER_49_787 VPWR VGND sg13g2_decap_8
XFILLER_17_640 VPWR VGND sg13g2_decap_8
XFILLER_36_437 VPWR VGND sg13g2_fill_2
XFILLER_45_982 VPWR VGND sg13g2_decap_8
X_3930_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] _1365_
+ _1317_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[5\] _1366_ _1312_ sg13g2_a221oi_1
X_3861_ net768 _1301_ _1302_ VPWR VGND sg13g2_nor2_2
XFILLER_32_665 VPWR VGND sg13g2_decap_8
X_2812_ VPWR VGND _0379_ net555 _0378_ _0225_ _0380_ net617 sg13g2_a221oi_1
XFILLER_20_849 VPWR VGND sg13g2_decap_8
X_3792_ _1253_ _1054_ _1252_ net600 sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\]
+ VPWR VGND sg13g2_a22oi_1
X_2743_ VGND VPWR _1611_ _1639_ _0312_ net689 sg13g2_a21oi_1
XFILLER_9_894 VPWR VGND sg13g2_decap_8
X_2674_ _1626_ VPWR _0266_ VGND _1589_ _1596_ sg13g2_o21ai_1
X_3226_ _0762_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[5\] net640 VPWR
+ VGND sg13g2_nand2_1
X_3157_ _0693_ net724 _1534_ VPWR VGND sg13g2_nand2_1
XFILLER_43_908 VPWR VGND sg13g2_decap_8
X_2108_ _1500_ _1528_ _1529_ VPWR VGND sg13g2_nor2_1
XFILLER_27_459 VPWR VGND sg13g2_decap_8
X_3088_ _1534_ VPWR _0624_ VGND net733 _0623_ sg13g2_o21ai_1
X_2039_ VPWR _1462_ sap_3_inst.alu.act\[0\] VGND sg13g2_inv_1
XFILLER_35_492 VPWR VGND sg13g2_decap_8
XFILLER_11_816 VPWR VGND sg13g2_decap_8
XFILLER_23_654 VPWR VGND sg13g2_decap_8
XFILLER_2_525 VPWR VGND sg13g2_decap_8
XFILLER_46_724 VPWR VGND sg13g2_decap_8
XFILLER_42_930 VPWR VGND sg13g2_decap_8
XFILLER_14_621 VPWR VGND sg13g2_decap_8
XFILLER_26_492 VPWR VGND sg13g2_decap_8
XFILLER_41_451 VPWR VGND sg13g2_decap_8
XFILLER_14_698 VPWR VGND sg13g2_decap_8
XFILLER_6_820 VPWR VGND sg13g2_decap_8
XFILLER_10_860 VPWR VGND sg13g2_decap_8
XFILLER_6_897 VPWR VGND sg13g2_decap_8
X_2390_ _1723_ _1810_ _1811_ VPWR VGND sg13g2_and2_1
X_4060_ net790 VGND VPWR _0038_ sap_3_inst.alu.acc\[4\] clknet_5_22__leaf_sap_3_inst.alu.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_49_584 VPWR VGND sg13g2_decap_8
X_3011_ _0564_ net744 sap_3_inst.alu.tmp\[7\] VPWR VGND sg13g2_nand2b_1
XFILLER_37_702 VPWR VGND sg13g2_decap_8
XFILLER_18_971 VPWR VGND sg13g2_decap_8
XFILLER_24_407 VPWR VGND sg13g2_decap_8
XFILLER_25_919 VPWR VGND sg13g2_decap_8
XFILLER_37_779 VPWR VGND sg13g2_decap_8
X_3913_ VPWR VGND _1350_ net764 _1344_ _1440_ _1351_ net762 sg13g2_a221oi_1
XFILLER_33_963 VPWR VGND sg13g2_decap_8
X_3844_ _1281_ VPWR _1289_ VGND net63 _1288_ sg13g2_o21ai_1
XFILLER_20_646 VPWR VGND sg13g2_decap_8
X_3775_ VGND VPWR _0955_ _0969_ _1241_ _0994_ sg13g2_a21oi_1
X_2726_ net65 sap_3_inst.out\[5\] net766 _0023_ VPWR VGND sg13g2_mux2_1
XFILLER_9_691 VPWR VGND sg13g2_decap_8
X_2657_ _0249_ _0250_ _1954_ _0251_ VPWR VGND sg13g2_nand3_1
X_2588_ _1858_ net545 _1998_ VPWR VGND sg13g2_nor2_1
XFILLER_47_27 VPWR VGND sg13g2_fill_2
XFILLER_41_1011 VPWR VGND sg13g2_decap_8
X_3209_ _0745_ net646 sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] net649
+ sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_28_757 VPWR VGND sg13g2_decap_8
X_4189_ net800 VGND VPWR _0167_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[5\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_43_705 VPWR VGND sg13g2_decap_8
XFILLER_24_974 VPWR VGND sg13g2_decap_8
XFILLER_11_613 VPWR VGND sg13g2_decap_8
XFILLER_3_801 VPWR VGND sg13g2_decap_8
XFILLER_3_878 VPWR VGND sg13g2_decap_8
Xfanout681 _1617_ net681 VPWR VGND sg13g2_buf_2
Xfanout670 _0314_ net670 VPWR VGND sg13g2_buf_8
Xfanout692 net693 net692 VPWR VGND sg13g2_buf_8
XFILLER_46_521 VPWR VGND sg13g2_decap_8
XFILLER_19_768 VPWR VGND sg13g2_decap_8
XFILLER_46_598 VPWR VGND sg13g2_decap_8
XFILLER_15_941 VPWR VGND sg13g2_decap_8
XFILLER_18_1013 VPWR VGND sg13g2_decap_8
XFILLER_14_495 VPWR VGND sg13g2_decap_8
XFILLER_30_955 VPWR VGND sg13g2_decap_8
X_3560_ VGND VPWR net9 _1078_ _1080_ _0829_ sg13g2_a21oi_1
X_2511_ VGND VPWR net725 net685 _1924_ _1821_ sg13g2_a21oi_1
X_3491_ _1020_ _1018_ _1019_ net612 _1490_ VPWR VGND sg13g2_a22oi_1
XFILLER_6_694 VPWR VGND sg13g2_decap_8
X_2442_ _1859_ _1860_ _1861_ VPWR VGND sg13g2_and2_1
X_2373_ _1746_ _1761_ _1793_ _1794_ VPWR VGND sg13g2_nor3_2
X_4112_ net775 VGND VPWR _0090_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\]
+ clknet_5_10__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_25_1017 VPWR VGND sg13g2_decap_8
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
X_4043_ net788 VGND VPWR _0025_ u_ser.shadow_reg\[7\] clknet_3_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_49_381 VPWR VGND sg13g2_decap_8
XFILLER_25_716 VPWR VGND sg13g2_decap_8
XFILLER_37_576 VPWR VGND sg13g2_decap_8
XFILLER_33_760 VPWR VGND sg13g2_decap_8
XFILLER_21_933 VPWR VGND sg13g2_decap_8
X_3827_ _1276_ net585 _1027_ VPWR VGND sg13g2_nand2_1
X_3758_ VGND VPWR _0873_ _0894_ _1228_ _1227_ sg13g2_a21oi_1
X_2709_ _1578_ _1642_ net694 _0288_ VPWR VGND sg13g2_nand3_1
X_3689_ _1046_ _1086_ _1184_ VPWR VGND sg13g2_nor2_2
XFILLER_0_848 VPWR VGND sg13g2_decap_8
XFILLER_48_808 VPWR VGND sg13g2_decap_8
XFILLER_43_502 VPWR VGND sg13g2_decap_8
XFILLER_28_554 VPWR VGND sg13g2_decap_8
XFILLER_15_226 VPWR VGND sg13g2_fill_1
XFILLER_31_708 VPWR VGND sg13g2_decap_8
XFILLER_43_579 VPWR VGND sg13g2_decap_8
XFILLER_24_771 VPWR VGND sg13g2_decap_8
XFILLER_8_937 VPWR VGND sg13g2_decap_8
XFILLER_11_465 VPWR VGND sg13g2_fill_1
XFILLER_12_966 VPWR VGND sg13g2_decap_8
XFILLER_3_675 VPWR VGND sg13g2_decap_8
XFILLER_2_141 VPWR VGND sg13g2_fill_2
XFILLER_24_8 VPWR VGND sg13g2_fill_1
XFILLER_46_351 VPWR VGND sg13g2_decap_8
XFILLER_19_565 VPWR VGND sg13g2_decap_8
XFILLER_47_885 VPWR VGND sg13g2_decap_8
XFILLER_46_395 VPWR VGND sg13g2_decap_8
XFILLER_22_708 VPWR VGND sg13g2_decap_8
XFILLER_34_557 VPWR VGND sg13g2_decap_8
X_2991_ _0553_ _0518_ _0552_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_752 VPWR VGND sg13g2_decap_8
X_3612_ _1125_ net579 VPWR VGND _1021_ sg13g2_nand2b_2
X_3543_ net558 _1065_ _1066_ VPWR VGND sg13g2_nor2_1
XFILLER_43_0 VPWR VGND sg13g2_fill_2
XFILLER_6_491 VPWR VGND sg13g2_decap_8
X_3474_ _1003_ VPWR _1004_ VGND net611 _0999_ sg13g2_o21ai_1
X_2425_ _1512_ _1844_ _1845_ _1846_ VPWR VGND sg13g2_nor3_1
X_2356_ _1777_ _1774_ _1544_ _1655_ net687 VPWR VGND sg13g2_a22oi_1
X_2287_ net695 _1622_ _1708_ VPWR VGND sg13g2_nor2_1
XFILLER_38_830 VPWR VGND sg13g2_decap_8
XFILLER_25_513 VPWR VGND sg13g2_decap_8
XFILLER_13_719 VPWR VGND sg13g2_decap_8
XFILLER_21_730 VPWR VGND sg13g2_decap_8
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_5_929 VPWR VGND sg13g2_decap_8
XFILLER_0_645 VPWR VGND sg13g2_decap_8
XFILLER_48_605 VPWR VGND sg13g2_decap_8
XFILLER_47_115 VPWR VGND sg13g2_fill_2
XFILLER_29_874 VPWR VGND sg13g2_decap_8
XFILLER_44_822 VPWR VGND sg13g2_decap_8
XFILLER_16_557 VPWR VGND sg13g2_decap_8
XFILLER_44_899 VPWR VGND sg13g2_decap_8
XFILLER_31_505 VPWR VGND sg13g2_decap_8
XFILLER_12_763 VPWR VGND sg13g2_decap_8
XFILLER_8_734 VPWR VGND sg13g2_decap_8
XFILLER_3_472 VPWR VGND sg13g2_decap_8
X_2210_ net680 _1629_ _1630_ _1631_ VPWR VGND sg13g2_nor3_1
X_3190_ _0657_ net665 _0711_ _0726_ VPWR VGND sg13g2_nor3_1
X_2141_ _1562_ net726 net728 VPWR VGND sg13g2_nand2_2
XFILLER_22_1009 VPWR VGND sg13g2_decap_8
XFILLER_39_649 VPWR VGND sg13g2_decap_8
X_2072_ VPWR _1495_ sap_3_inst.reg_file.array_serializer_inst.data\[4\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_35_800 VPWR VGND sg13g2_decap_8
XFILLER_47_682 VPWR VGND sg13g2_decap_8
XFILLER_22_505 VPWR VGND sg13g2_decap_8
XFILLER_35_877 VPWR VGND sg13g2_decap_8
X_2974_ _1936_ VPWR _0536_ VGND _0534_ _0535_ sg13g2_o21ai_1
X_3526_ _0077_ _1049_ _1051_ net557 _1454_ VPWR VGND sg13g2_a22oi_1
X_3457_ _0072_ _0981_ _0985_ net562 _1475_ VPWR VGND sg13g2_a22oi_1
X_2408_ _1829_ _1828_ sap_3_inst.alu.flags\[7\] _1827_ net743 VPWR VGND sg13g2_a22oi_1
X_3388_ _0921_ net577 _0920_ VPWR VGND sg13g2_nand2_2
X_2339_ _1752_ _1755_ _1756_ _1759_ _1760_ VPWR VGND sg13g2_and4_1
X_4009_ net68 u_ser.state\[1\] net766 _0189_ VPWR VGND sg13g2_a21o_1
XFILLER_26_800 VPWR VGND sg13g2_decap_8
XFILLER_38_1005 VPWR VGND sg13g2_decap_8
XFILLER_13_516 VPWR VGND sg13g2_decap_8
XFILLER_26_877 VPWR VGND sg13g2_decap_8
XFILLER_41_836 VPWR VGND sg13g2_decap_8
XFILLER_40_357 VPWR VGND sg13g2_fill_1
XFILLER_9_509 VPWR VGND sg13g2_decap_8
XFILLER_5_726 VPWR VGND sg13g2_decap_8
XFILLER_1_954 VPWR VGND sg13g2_decap_8
XFILLER_48_402 VPWR VGND sg13g2_decap_8
XFILLER_0_442 VPWR VGND sg13g2_decap_8
XFILLER_49_969 VPWR VGND sg13g2_decap_8
XFILLER_36_619 VPWR VGND sg13g2_decap_8
XFILLER_48_479 VPWR VGND sg13g2_decap_8
XFILLER_17_822 VPWR VGND sg13g2_decap_8
XFILLER_29_671 VPWR VGND sg13g2_decap_8
XFILLER_17_899 VPWR VGND sg13g2_decap_8
XFILLER_44_696 VPWR VGND sg13g2_decap_8
XFILLER_32_847 VPWR VGND sg13g2_decap_8
XFILLER_8_531 VPWR VGND sg13g2_decap_8
XFILLER_12_560 VPWR VGND sg13g2_decap_8
X_2690_ VPWR VGND _1499_ _0281_ _1528_ _1508_ _0282_ net712 sg13g2_a221oi_1
X_3311_ VPWR _0847_ _0846_ VGND sg13g2_inv_1
X_3242_ sap_3_inst.reg_file.array_serializer_inst.data\[9\]\[3\] net656 _0778_ VPWR
+ VGND sg13g2_and2_1
X_3173_ net702 VPWR _0709_ VGND _0706_ _0707_ sg13g2_o21ai_1
X_2124_ _1545_ net698 _1542_ VPWR VGND sg13g2_nand2_1
X_2055_ VPWR _1478_ sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[5\] VGND
+ sg13g2_inv_1
Xclkbuf_5_30__f_sap_3_inst.alu.clk_regs clknet_4_15_0_sap_3_inst.alu.clk_regs clknet_5_30__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_35_674 VPWR VGND sg13g2_decap_8
XFILLER_23_836 VPWR VGND sg13g2_decap_8
XFILLER_22_346 VPWR VGND sg13g2_fill_1
X_2957_ VGND VPWR _0333_ _0506_ _0520_ net563 sg13g2_a21oi_1
X_2888_ _0324_ _0451_ _0453_ VPWR VGND _0452_ sg13g2_nand3b_1
XFILLER_2_707 VPWR VGND sg13g2_decap_8
X_3509_ _1036_ net571 _0635_ _1037_ VPWR VGND sg13g2_a21o_1
XFILLER_46_906 VPWR VGND sg13g2_decap_8
XFILLER_14_803 VPWR VGND sg13g2_decap_8
XFILLER_25_151 VPWR VGND sg13g2_fill_2
XFILLER_26_674 VPWR VGND sg13g2_decap_8
XFILLER_41_633 VPWR VGND sg13g2_decap_8
XFILLER_13_302 VPWR VGND sg13g2_fill_1
XFILLER_13_368 VPWR VGND sg13g2_fill_1
XFILLER_40_132 VPWR VGND sg13g2_fill_1
XFILLER_9_339 VPWR VGND sg13g2_fill_1
XFILLER_40_176 VPWR VGND sg13g2_fill_2
XFILLER_12_1008 VPWR VGND sg13g2_decap_8
XFILLER_5_523 VPWR VGND sg13g2_decap_8
XFILLER_1_751 VPWR VGND sg13g2_decap_8
XFILLER_49_766 VPWR VGND sg13g2_decap_8
XFILLER_45_961 VPWR VGND sg13g2_decap_8
XFILLER_16_140 VPWR VGND sg13g2_fill_1
XFILLER_44_493 VPWR VGND sg13g2_decap_8
XFILLER_16_173 VPWR VGND sg13g2_fill_1
XFILLER_17_696 VPWR VGND sg13g2_decap_8
X_3860_ VGND VPWR _1301_ _1300_ _1497_ sg13g2_or2_1
XFILLER_32_644 VPWR VGND sg13g2_decap_8
X_2811_ VGND VPWR sap_3_inst.alu.act\[1\] net670 _0379_ net617 sg13g2_a21oi_1
XFILLER_13_880 VPWR VGND sg13g2_decap_8
XFILLER_20_828 VPWR VGND sg13g2_decap_8
X_3791_ net656 _1055_ _1252_ VPWR VGND sg13g2_and2_1
X_2742_ VGND VPWR _0311_ net617 _1938_ sg13g2_or2_1
XFILLER_9_873 VPWR VGND sg13g2_decap_8
X_2673_ _0265_ _1646_ _1592_ _1637_ net707 VPWR VGND sg13g2_a22oi_1
X_3225_ _0761_ net643 sap_3_inst.reg_file.array_serializer_inst.data\[7\]\[5\] net646
+ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_243 VPWR VGND sg13g2_fill_2
X_3156_ _0692_ _1534_ _0623_ VPWR VGND sg13g2_nand2_1
XFILLER_28_939 VPWR VGND sg13g2_decap_8
X_3087_ _0623_ net698 _1712_ VPWR VGND sg13g2_nand2_1
X_2107_ _1528_ net719 sap_3_inst.controller.stage\[1\] VPWR VGND sg13g2_nand2_2
XFILLER_27_438 VPWR VGND sg13g2_decap_8
X_2038_ VPWR _1461_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[0\] VGND
+ sg13g2_inv_1
XFILLER_36_983 VPWR VGND sg13g2_decap_8
XFILLER_23_633 VPWR VGND sg13g2_decap_8
X_3989_ _1407_ sap_3_inst.alu.act\[7\] net548 VPWR VGND sg13g2_nand2_1
XFILLER_2_504 VPWR VGND sg13g2_decap_8
XFILLER_46_703 VPWR VGND sg13g2_decap_8
XFILLER_14_600 VPWR VGND sg13g2_decap_8
XFILLER_26_471 VPWR VGND sg13g2_decap_8
XFILLER_42_986 VPWR VGND sg13g2_decap_8
XFILLER_14_677 VPWR VGND sg13g2_decap_8
XFILLER_6_876 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_fill_2
XFILLER_3_11 VPWR VGND sg13g2_fill_2
XFILLER_49_563 VPWR VGND sg13g2_decap_8
XFILLER_3_99 VPWR VGND sg13g2_decap_4
X_3010_ sap_3_inst.alu.acc\[7\] sap_3_inst.alu.tmp\[7\] _0563_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_758 VPWR VGND sg13g2_decap_8
XFILLER_18_950 VPWR VGND sg13g2_decap_8
XFILLER_17_460 VPWR VGND sg13g2_fill_2
X_3912_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[3\] _1349_
+ _1308_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[3\] _1350_ _1305_ sg13g2_a221oi_1
XFILLER_33_942 VPWR VGND sg13g2_decap_8
X_3843_ net769 _1282_ sap_3_inst.reg_file.array_serializer_inst.bit_pos\[1\] _1288_
+ VPWR VGND sg13g2_nand3_1
XFILLER_20_625 VPWR VGND sg13g2_decap_8
X_3774_ _0136_ _0984_ _1240_ net598 _1476_ VPWR VGND sg13g2_a22oi_1
XFILLER_9_670 VPWR VGND sg13g2_decap_8
X_2725_ net74 sap_3_inst.out\[4\] net766 _0022_ VPWR VGND sg13g2_mux2_1
X_2656_ net757 net759 net749 net752 _0250_ VPWR VGND sg13g2_nor4_1
X_2587_ _1986_ _1723_ _1997_ net545 VPWR VGND sg13g2_a21o_2
X_4188_ net794 VGND VPWR _0166_ sap_3_inst.reg_file.array_serializer_inst.shadow_reg\[4\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
X_3208_ _0743_ VPWR _0744_ VGND _0736_ _0742_ sg13g2_o21ai_1
X_3139_ _0675_ _1535_ _1633_ VPWR VGND sg13g2_nand2_1
XFILLER_28_736 VPWR VGND sg13g2_decap_8
Xclkbuf_5_27__f_sap_3_inst.alu.clk_regs clknet_4_13_0_sap_3_inst.alu.clk_regs clknet_5_27__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_36_780 VPWR VGND sg13g2_decap_8
XFILLER_24_953 VPWR VGND sg13g2_decap_8
XFILLER_23_452 VPWR VGND sg13g2_fill_2
XFILLER_10_168 VPWR VGND sg13g2_fill_1
XFILLER_7_629 VPWR VGND sg13g2_decap_8
XFILLER_11_669 VPWR VGND sg13g2_decap_8
XFILLER_12_75 VPWR VGND sg13g2_fill_1
XFILLER_3_857 VPWR VGND sg13g2_decap_8
Xfanout660 _0625_ net660 VPWR VGND sg13g2_buf_8
XFILLER_46_500 VPWR VGND sg13g2_decap_8
Xfanout682 _1714_ net682 VPWR VGND sg13g2_buf_8
Xfanout693 _1532_ net693 VPWR VGND sg13g2_buf_8
Xfanout671 net672 net671 VPWR VGND sg13g2_buf_8
XFILLER_19_747 VPWR VGND sg13g2_decap_8
XFILLER_46_577 VPWR VGND sg13g2_decap_8
XFILLER_15_920 VPWR VGND sg13g2_decap_8
XFILLER_34_739 VPWR VGND sg13g2_decap_8
XFILLER_42_783 VPWR VGND sg13g2_decap_8
XFILLER_15_997 VPWR VGND sg13g2_decap_8
XFILLER_41_282 VPWR VGND sg13g2_fill_2
XFILLER_30_934 VPWR VGND sg13g2_decap_8
X_3490_ VPWR VGND sap_3_inst.reg_file.array_serializer_inst.data\[1\]\[7\] _1017_
+ net587 sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[7\] _1019_ net592 sg13g2_a221oi_1
X_2510_ _1923_ _1546_ net688 VPWR VGND sg13g2_nand2_1
XFILLER_6_673 VPWR VGND sg13g2_decap_8
X_2441_ _1860_ _1801_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[6\] _1797_
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[6\] VPWR VGND sg13g2_a22oi_1
X_2372_ VGND VPWR _1793_ _1790_ _1772_ sg13g2_or2_1
X_4111_ net780 VGND VPWR _0089_ sap_3_inst.reg_file.array_serializer_inst.data\[2\]\[6\]
+ clknet_5_13__leaf_sap_3_inst.alu.clk_regs sg13g2_dfrbpq_2
XFILLER_49_360 VPWR VGND sg13g2_decap_8
X_4042_ net788 VGND VPWR _0024_ u_ser.shadow_reg\[6\] clknet_3_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_37_555 VPWR VGND sg13g2_decap_8
XFILLER_21_912 VPWR VGND sg13g2_decap_8
XFILLER_21_989 VPWR VGND sg13g2_decap_8
X_3826_ _0153_ _1114_ _1275_ net605 _1481_ VPWR VGND sg13g2_a22oi_1
XFILLER_20_499 VPWR VGND sg13g2_decap_8
X_3757_ _0844_ VPWR _1227_ VGND _0873_ _0894_ sg13g2_o21ai_1
X_2708_ VPWR VGND _1655_ net681 net687 net700 _0287_ _1553_ sg13g2_a221oi_1
XFILLER_3_109 VPWR VGND sg13g2_fill_1
X_3688_ _1181_ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[0\] _1183_ _0107_
+ VPWR VGND sg13g2_a21o_1
X_2639_ _0234_ net619 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[0\] net632
+ sap_3_inst.reg_file.array_serializer_inst.data\[10\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_0_827 VPWR VGND sg13g2_decap_8
XFILLER_28_533 VPWR VGND sg13g2_decap_8
XFILLER_16_739 VPWR VGND sg13g2_decap_8
XFILLER_43_558 VPWR VGND sg13g2_decap_8
XFILLER_24_750 VPWR VGND sg13g2_decap_8
XFILLER_12_945 VPWR VGND sg13g2_decap_8
XFILLER_23_282 VPWR VGND sg13g2_fill_1
XFILLER_8_916 VPWR VGND sg13g2_decap_8
XFILLER_23_52 VPWR VGND sg13g2_fill_2
XFILLER_48_1018 VPWR VGND sg13g2_decap_8
XFILLER_3_654 VPWR VGND sg13g2_decap_8
XFILLER_2_131 VPWR VGND sg13g2_decap_4
XFILLER_47_864 VPWR VGND sg13g2_decap_8
XFILLER_0_23 VPWR VGND sg13g2_fill_1
XFILLER_0_1009 VPWR VGND sg13g2_decap_8
XFILLER_19_544 VPWR VGND sg13g2_decap_8
XFILLER_46_374 VPWR VGND sg13g2_decap_8
XFILLER_0_89 VPWR VGND sg13g2_decap_8
XFILLER_34_536 VPWR VGND sg13g2_decap_8
X_2990_ _0552_ _0540_ _0551_ VPWR VGND sg13g2_xnor2_1
XFILLER_42_580 VPWR VGND sg13g2_decap_8
XFILLER_14_271 VPWR VGND sg13g2_fill_2
XFILLER_15_794 VPWR VGND sg13g2_decap_8
XFILLER_30_731 VPWR VGND sg13g2_decap_8
X_3611_ net591 _1123_ _1124_ VPWR VGND sg13g2_nor2_1
X_3542_ net576 _0987_ _1065_ VPWR VGND sg13g2_nor2_1
XFILLER_7_993 VPWR VGND sg13g2_decap_8
X_3473_ VGND VPWR net611 _1001_ _1003_ net575 sg13g2_a21oi_1
X_2424_ _1540_ net685 _1845_ VPWR VGND sg13g2_and2_1
X_2355_ _1614_ VPWR _1776_ VGND _1698_ _1728_ sg13g2_o21ai_1
X_2286_ net696 _1687_ _1688_ _1707_ VPWR VGND sg13g2_or3_1
XFILLER_38_886 VPWR VGND sg13g2_decap_8
XFILLER_25_569 VPWR VGND sg13g2_decap_8
XFILLER_21_786 VPWR VGND sg13g2_decap_8
X_3809_ net11 net603 _1263_ VPWR VGND sg13g2_nor2_1
XFILLER_5_908 VPWR VGND sg13g2_decap_8
XFILLER_0_624 VPWR VGND sg13g2_decap_8
XFILLER_29_853 VPWR VGND sg13g2_decap_8
XFILLER_44_801 VPWR VGND sg13g2_decap_8
XFILLER_16_536 VPWR VGND sg13g2_decap_8
XFILLER_44_878 VPWR VGND sg13g2_decap_8
XFILLER_8_713 VPWR VGND sg13g2_decap_8
XFILLER_12_742 VPWR VGND sg13g2_decap_8
XFILLER_4_985 VPWR VGND sg13g2_decap_8
XFILLER_3_451 VPWR VGND sg13g2_decap_8
X_2140_ net726 net728 _1561_ VPWR VGND sg13g2_and2_1
XFILLER_39_628 VPWR VGND sg13g2_decap_8
X_2071_ VPWR _1494_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_47_661 VPWR VGND sg13g2_decap_8
XFILLER_35_856 VPWR VGND sg13g2_decap_8
X_2973_ _0535_ net743 net671 VPWR VGND sg13g2_xnor2_1
XFILLER_15_591 VPWR VGND sg13g2_decap_8
XFILLER_7_790 VPWR VGND sg13g2_decap_8
X_3525_ net557 _1050_ _1051_ VPWR VGND sg13g2_nor2_1
X_3456_ _0986_ VPWR _0987_ VGND net559 _0854_ sg13g2_o21ai_1
X_2407_ net723 _1584_ _1647_ _1828_ VPWR VGND sg13g2_nor3_2
X_3387_ _0916_ _0897_ _0919_ _0920_ VPWR VGND sg13g2_a21o_1
X_2338_ _1751_ net679 _1758_ _1759_ VPWR VGND sg13g2_nor3_1
X_2269_ _1528_ _1557_ _1690_ VPWR VGND sg13g2_nor2_2
XFILLER_44_119 VPWR VGND sg13g2_fill_2
X_4008_ VPWR _0188_ _1423_ VGND sg13g2_inv_1
XFILLER_38_683 VPWR VGND sg13g2_decap_8
XFILLER_26_856 VPWR VGND sg13g2_decap_8
XFILLER_41_815 VPWR VGND sg13g2_decap_8
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_21_583 VPWR VGND sg13g2_decap_8
XFILLER_5_705 VPWR VGND sg13g2_decap_8
XFILLER_1_933 VPWR VGND sg13g2_decap_8
XFILLER_49_948 VPWR VGND sg13g2_decap_8
XFILLER_0_498 VPWR VGND sg13g2_decap_8
XFILLER_48_458 VPWR VGND sg13g2_decap_8
XFILLER_21_1010 VPWR VGND sg13g2_decap_8
XFILLER_17_801 VPWR VGND sg13g2_decap_8
XFILLER_29_650 VPWR VGND sg13g2_decap_8
XFILLER_44_675 VPWR VGND sg13g2_decap_8
XFILLER_17_878 VPWR VGND sg13g2_decap_8
XFILLER_16_377 VPWR VGND sg13g2_fill_1
XFILLER_31_303 VPWR VGND sg13g2_fill_1
XFILLER_32_826 VPWR VGND sg13g2_decap_8
XFILLER_8_510 VPWR VGND sg13g2_decap_8
Xclkbuf_5_1__f_sap_3_inst.alu.clk_regs clknet_4_0_0_sap_3_inst.alu.clk_regs clknet_5_1__leaf_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_8_587 VPWR VGND sg13g2_decap_8
X_3310_ net575 VPWR _0846_ VGND net561 net574 sg13g2_o21ai_1
XFILLER_4_782 VPWR VGND sg13g2_decap_8
X_3241_ sap_3_inst.reg_file.array_serializer_inst.data\[11\]\[3\] net608 _0777_ VPWR
+ VGND sg13g2_and2_1
X_3172_ _0708_ net713 _1782_ VPWR VGND sg13g2_nand2b_1
X_2123_ _1500_ _1528_ _1543_ _1544_ VPWR VGND sg13g2_nor3_1
X_2054_ VPWR _1477_ sap_3_inst.reg_file.array_serializer_inst.data\[6\]\[5\] VGND
+ sg13g2_inv_1
XFILLER_23_815 VPWR VGND sg13g2_decap_8
XFILLER_35_653 VPWR VGND sg13g2_decap_8
X_2956_ _0325_ _0517_ _0518_ _0519_ VPWR VGND sg13g2_nor3_1
X_2887_ _0426_ _0450_ _0452_ VPWR VGND sg13g2_nor2_1
Xclkbuf_0_sap_3_inst.alu.clk_regs sap_3_inst.alu.clk_regs clknet_0_sap_3_inst.alu.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3508_ VGND VPWR _0610_ net614 _1036_ net587 sg13g2_a21oi_1
X_3439_ _0970_ _0967_ _0968_ VPWR VGND sg13g2_nand2_2
XFILLER_38_480 VPWR VGND sg13g2_decap_8
XFILLER_39_992 VPWR VGND sg13g2_decap_8
XFILLER_26_653 VPWR VGND sg13g2_decap_8
XFILLER_41_612 VPWR VGND sg13g2_decap_8
XFILLER_14_859 VPWR VGND sg13g2_decap_8
XFILLER_41_689 VPWR VGND sg13g2_decap_8
XFILLER_5_502 VPWR VGND sg13g2_decap_8
XFILLER_5_579 VPWR VGND sg13g2_decap_8
Xoutput30 net30 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_730 VPWR VGND sg13g2_decap_8
XFILLER_49_745 VPWR VGND sg13g2_decap_8
XFILLER_45_940 VPWR VGND sg13g2_decap_8
XFILLER_44_472 VPWR VGND sg13g2_decap_8
XFILLER_17_675 VPWR VGND sg13g2_decap_8
XFILLER_32_623 VPWR VGND sg13g2_decap_8
XFILLER_20_807 VPWR VGND sg13g2_decap_8
X_2810_ _0377_ VPWR _0378_ VGND net544 _0376_ sg13g2_o21ai_1
X_3790_ _0141_ _1049_ _1251_ net600 _1447_ VPWR VGND sg13g2_a22oi_1
XFILLER_31_155 VPWR VGND sg13g2_fill_2
XFILLER_9_852 VPWR VGND sg13g2_decap_8
X_2741_ _0309_ VPWR _0310_ VGND _1675_ _0298_ sg13g2_o21ai_1
XFILLER_8_384 VPWR VGND sg13g2_fill_2
X_2672_ _0262_ _0263_ _0264_ VPWR VGND sg13g2_nor2_1
XFILLER_28_1016 VPWR VGND sg13g2_decap_8
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
X_3224_ _0760_ net649 sap_3_inst.reg_file.array_serializer_inst.data\[8\]\[5\] net651
+ sap_3_inst.reg_file.array_serializer_inst.data\[5\]\[5\] VPWR VGND sg13g2_a22oi_1
.ends

