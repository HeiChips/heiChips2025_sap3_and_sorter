* NGSPICE file created from heichips25_sap3.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_lgcp_1 abstract view
.subckt sg13g2_lgcp_1 GATE CLK GCLK VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

.subckt heichips25_sap3 VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
X_3155_ VGND VPWR net718 _1941_ _0064_ _0627_ sg13g2_a21oi_1
XFILLER_28_918 VPWR VGND sg13g2_decap_8
X_3086_ net772 _0334_ _0583_ VPWR VGND sg13g2_nor2_1
X_2106_ VPWR _1524_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[0\]
+ VGND sg13g2_inv_1
XFILLER_36_995 VPWR VGND sg13g2_decap_8
XFILLER_23_634 VPWR VGND sg13g2_decap_8
XFILLER_35_1009 VPWR VGND sg13g2_decap_8
X_3988_ _1364_ net48 net798 VPWR VGND sg13g2_nand2_1
X_2939_ VPWR _0440_ _0439_ VGND sg13g2_inv_1
XFILLER_11_1020 VPWR VGND sg13g2_decap_8
XFILLER_2_505 VPWR VGND sg13g2_decap_8
Xfanout820 net826 net820 VPWR VGND sg13g2_buf_8
Xfanout831 net832 net831 VPWR VGND sg13g2_buf_8
XFILLER_46_748 VPWR VGND sg13g2_decap_8
XFILLER_27_973 VPWR VGND sg13g2_decap_8
XFILLER_42_954 VPWR VGND sg13g2_decap_8
XFILLER_41_453 VPWR VGND sg13g2_decap_8
XFILLER_14_667 VPWR VGND sg13g2_decap_8
XFILLER_9_126 VPWR VGND sg13g2_fill_2
XFILLER_9_159 VPWR VGND sg13g2_fill_1
XFILLER_6_855 VPWR VGND sg13g2_decap_8
XFILLER_10_884 VPWR VGND sg13g2_decap_8
XFILLER_3_56 VPWR VGND sg13g2_fill_2
XFILLER_49_531 VPWR VGND sg13g2_decap_8
XFILLER_3_67 VPWR VGND sg13g2_fill_1
XFILLER_37_726 VPWR VGND sg13g2_decap_8
XFILLER_24_409 VPWR VGND sg13g2_decap_8
XFILLER_45_792 VPWR VGND sg13g2_decap_8
XFILLER_18_984 VPWR VGND sg13g2_decap_8
XFILLER_33_932 VPWR VGND sg13g2_decap_8
X_3911_ net593 VPWR _1298_ VGND net647 _0969_ sg13g2_o21ai_1
X_3842_ _1243_ VPWR _0130_ VGND _1244_ _1248_ sg13g2_o21ai_1
XFILLER_20_637 VPWR VGND sg13g2_decap_8
XFILLER_32_497 VPWR VGND sg13g2_decap_8
X_3773_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[7\] net675 _1205_
+ VPWR VGND sg13g2_nor2_1
X_2724_ VGND VPWR net1 _1884_ _0254_ _0253_ sg13g2_a21oi_1
X_2655_ _2062_ _1864_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[3\]
+ net625 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2586_ VPWR VGND _1496_ _1994_ _1894_ _1595_ _1995_ net722 sg13g2_a221oi_1
X_4325_ net823 VGND VPWR _0182_ sap_3_inst.alu_inst.act\[5\] clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4256_ net809 VGND VPWR _0113_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[7\]
+ clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_41_1013 VPWR VGND sg13g2_decap_8
X_3207_ _0678_ _0677_ _0672_ _0676_ _1670_ VPWR VGND sg13g2_a22oi_1
X_4187_ net821 VGND VPWR _0044_ sap_3_inst.out\[3\] clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_28_715 VPWR VGND sg13g2_decap_8
X_3138_ _0619_ VPWR _0055_ VGND _1967_ net701 sg13g2_o21ai_1
X_3069_ VPWR _0039_ _0566_ VGND sg13g2_inv_1
XFILLER_23_431 VPWR VGND sg13g2_decap_8
XFILLER_36_792 VPWR VGND sg13g2_decap_8
XFILLER_24_976 VPWR VGND sg13g2_decap_8
XFILLER_3_847 VPWR VGND sg13g2_decap_8
Xfanout650 net651 net650 VPWR VGND sg13g2_buf_1
Xfanout694 _0330_ net694 VPWR VGND sg13g2_buf_2
Xclkbuf_5_21__f_sap_3_inst.alu_inst.clk_regs clknet_4_10_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
Xfanout672 net673 net672 VPWR VGND sg13g2_buf_8
Xfanout683 net685 net683 VPWR VGND sg13g2_buf_8
Xfanout661 net662 net661 VPWR VGND sg13g2_buf_8
XFILLER_46_545 VPWR VGND sg13g2_decap_8
XFILLER_37_73 VPWR VGND sg13g2_fill_2
XFILLER_15_910 VPWR VGND sg13g2_decap_8
XFILLER_27_770 VPWR VGND sg13g2_decap_8
XFILLER_42_751 VPWR VGND sg13g2_decap_8
XFILLER_15_987 VPWR VGND sg13g2_decap_8
XFILLER_18_1026 VPWR VGND sg13g2_fill_2
XFILLER_30_924 VPWR VGND sg13g2_decap_8
XFILLER_10_681 VPWR VGND sg13g2_decap_8
XFILLER_6_652 VPWR VGND sg13g2_decap_8
X_2440_ VPWR _1857_ net621 VGND sg13g2_inv_1
XFILLER_5_195 VPWR VGND sg13g2_fill_1
X_2371_ _1783_ _1784_ _1774_ _1788_ VPWR VGND _1787_ sg13g2_nand4_1
Xclkbuf_5_10__f_sap_3_inst.alu_inst.clk_regs clknet_4_5_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
X_4110_ _1463_ _0578_ net698 VPWR VGND sg13g2_nand2_1
X_4041_ _1313_ net51 _1411_ _0166_ VPWR VGND sg13g2_a21o_1
XFILLER_37_523 VPWR VGND sg13g2_decap_8
XFILLER_18_781 VPWR VGND sg13g2_decap_8
XFILLER_17_280 VPWR VGND sg13g2_fill_1
XFILLER_21_902 VPWR VGND sg13g2_decap_8
XFILLER_20_434 VPWR VGND sg13g2_fill_1
XFILLER_21_979 VPWR VGND sg13g2_decap_8
X_3825_ _1216_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[3\] net635
+ _0125_ VPWR VGND sg13g2_mux2_1
X_3756_ VGND VPWR _1188_ _1190_ _1191_ net656 sg13g2_a21oi_1
X_2707_ _0237_ VPWR _0026_ VGND _2057_ _0236_ sg13g2_o21ai_1
X_3687_ net15 _1097_ _1136_ VPWR VGND sg13g2_nor2_1
X_2638_ net696 net627 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[1\]
+ _2047_ VPWR VGND sg13g2_nand3_1
X_2569_ _1980_ _1509_ _1900_ VPWR VGND sg13g2_nand2_1
X_4308_ net835 VGND VPWR _0165_ sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[4\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
X_4239_ net814 VGND VPWR _0096_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[6\]
+ clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_28_512 VPWR VGND sg13g2_decap_8
XFILLER_28_589 VPWR VGND sg13g2_decap_8
XFILLER_23_250 VPWR VGND sg13g2_fill_1
XFILLER_24_773 VPWR VGND sg13g2_decap_8
XFILLER_8_906 VPWR VGND sg13g2_decap_8
XFILLER_12_968 VPWR VGND sg13g2_decap_8
XFILLER_3_644 VPWR VGND sg13g2_decap_8
XFILLER_47_865 VPWR VGND sg13g2_decap_8
XFILLER_46_342 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_567 VPWR VGND sg13g2_decap_8
XFILLER_15_784 VPWR VGND sg13g2_decap_8
XFILLER_30_721 VPWR VGND sg13g2_decap_8
XFILLER_9_88 VPWR VGND sg13g2_decap_8
XFILLER_9_55 VPWR VGND sg13g2_fill_2
XFILLER_9_99 VPWR VGND sg13g2_fill_1
XFILLER_30_798 VPWR VGND sg13g2_decap_8
X_3610_ VGND VPWR _1069_ _1070_ _0957_ _0861_ sg13g2_a21oi_2
X_3541_ net586 _1006_ _1007_ VPWR VGND sg13g2_nor2_2
XFILLER_7_961 VPWR VGND sg13g2_decap_8
X_3472_ _0939_ VPWR _0940_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[3\]
+ net662 sg13g2_o21ai_1
XFILLER_43_2 VPWR VGND sg13g2_fill_1
X_2423_ net713 _1833_ _1836_ _1839_ _1840_ VPWR VGND sg13g2_nor4_1
X_2354_ _1759_ _1770_ _1771_ VPWR VGND sg13g2_nor2_1
X_2285_ VGND VPWR _1630_ _1685_ _1702_ net735 sg13g2_a21oi_1
XFILLER_38_832 VPWR VGND sg13g2_decap_8
X_4024_ _1396_ _1349_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[4\]
+ _1346_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_37_320 VPWR VGND sg13g2_fill_2
Xheichips25_sap3_34 VPWR VGND uo_out[7] sg13g2_tielo
XFILLER_25_548 VPWR VGND sg13g2_decap_8
XFILLER_20_242 VPWR VGND sg13g2_fill_2
X_3808_ net657 _1074_ _1227_ VPWR VGND sg13g2_nor2_1
XFILLER_20_275 VPWR VGND sg13g2_fill_1
XFILLER_21_776 VPWR VGND sg13g2_decap_8
X_3739_ VPWR _0099_ _1176_ VGND sg13g2_inv_1
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_29_810 VPWR VGND sg13g2_decap_8
XFILLER_44_813 VPWR VGND sg13g2_decap_8
XFILLER_29_887 VPWR VGND sg13g2_decap_8
XFILLER_16_548 VPWR VGND sg13g2_decap_8
XFILLER_24_570 VPWR VGND sg13g2_decap_8
XFILLER_8_703 VPWR VGND sg13g2_decap_8
XFILLER_12_765 VPWR VGND sg13g2_decap_8
XFILLER_7_224 VPWR VGND sg13g2_fill_2
XFILLER_4_942 VPWR VGND sg13g2_decap_8
X_2070_ VPWR _1488_ u_ser.state\[0\] VGND sg13g2_inv_1
XFILLER_47_662 VPWR VGND sg13g2_decap_8
XFILLER_46_150 VPWR VGND sg13g2_fill_1
XFILLER_35_813 VPWR VGND sg13g2_decap_8
X_2972_ _0472_ net704 _0470_ VPWR VGND sg13g2_nand2_1
XFILLER_15_581 VPWR VGND sg13g2_decap_8
XFILLER_22_529 VPWR VGND sg13g2_decap_8
XFILLER_30_595 VPWR VGND sg13g2_decap_8
X_3524_ _0989_ VPWR _0990_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[5\]
+ net661 sg13g2_o21ai_1
X_3455_ _0719_ net648 _0924_ VPWR VGND sg13g2_nor2_1
X_2406_ _1823_ net759 _1762_ VPWR VGND sg13g2_nand2_1
X_3386_ _0720_ net659 _0857_ VPWR VGND sg13g2_nor2_2
X_2337_ _1636_ _1642_ net720 _1754_ VPWR VGND sg13g2_nor3_1
X_2268_ _1685_ _1679_ net738 net732 net737 VPWR VGND sg13g2_a22oi_1
XFILLER_26_824 VPWR VGND sg13g2_decap_8
X_4007_ VGND VPWR _1501_ net795 _1381_ _1313_ sg13g2_a21oi_1
X_2199_ _1616_ net767 net770 VPWR VGND sg13g2_nand2_2
XFILLER_37_161 VPWR VGND sg13g2_fill_1
XFILLER_38_1007 VPWR VGND sg13g2_decap_8
XFILLER_41_838 VPWR VGND sg13g2_decap_8
XFILLER_13_529 VPWR VGND sg13g2_decap_8
XFILLER_21_573 VPWR VGND sg13g2_decap_8
XFILLER_1_912 VPWR VGND sg13g2_decap_8
XFILLER_49_916 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
Xhold30 sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[0\] VPWR VGND net77
+ sg13g2_dlygate4sd3_1
XFILLER_1_989 VPWR VGND sg13g2_decap_8
XFILLER_48_437 VPWR VGND sg13g2_decap_8
XFILLER_21_1000 VPWR VGND sg13g2_decap_8
XFILLER_44_610 VPWR VGND sg13g2_decap_8
XFILLER_17_835 VPWR VGND sg13g2_decap_8
XFILLER_29_684 VPWR VGND sg13g2_decap_8
XFILLER_32_805 VPWR VGND sg13g2_decap_8
XFILLER_44_687 VPWR VGND sg13g2_decap_8
XFILLER_31_304 VPWR VGND sg13g2_fill_1
XFILLER_8_500 VPWR VGND sg13g2_decap_8
XFILLER_12_562 VPWR VGND sg13g2_decap_8
XFILLER_8_577 VPWR VGND sg13g2_decap_8
X_3240_ _0707_ _0710_ _0711_ VPWR VGND sg13g2_and2_1
X_3171_ VPWR VGND net715 net719 _0632_ net759 _0642_ _1886_ sg13g2_a221oi_1
XFILLER_6_1027 VPWR VGND sg13g2_fill_2
XFILLER_6_1016 VPWR VGND sg13g2_decap_8
X_2122_ VPWR _1540_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[6\]
+ VGND sg13g2_inv_1
XFILLER_35_610 VPWR VGND sg13g2_decap_8
XFILLER_23_816 VPWR VGND sg13g2_decap_8
XFILLER_35_687 VPWR VGND sg13g2_decap_8
X_2955_ _0456_ _0453_ _0455_ VPWR VGND sg13g2_xnor2_1
X_2886_ VPWR _0389_ _0388_ VGND sg13g2_inv_1
X_3507_ _0974_ _0862_ _0973_ VPWR VGND sg13g2_nand2_1
X_3438_ _0907_ net677 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[2\]
+ net688 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[2\] VPWR VGND sg13g2_a22oi_1
X_3369_ _0840_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[1\] net671
+ VPWR VGND sg13g2_nand2_1
XFILLER_45_407 VPWR VGND sg13g2_decap_8
XFILLER_26_621 VPWR VGND sg13g2_decap_8
XFILLER_14_849 VPWR VGND sg13g2_decap_8
XFILLER_26_698 VPWR VGND sg13g2_decap_8
XFILLER_41_635 VPWR VGND sg13g2_decap_8
XFILLER_15_43 VPWR VGND sg13g2_fill_2
XFILLER_22_893 VPWR VGND sg13g2_decap_8
XFILLER_5_569 VPWR VGND sg13g2_decap_8
Xoutput20 net32 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_49_713 VPWR VGND sg13g2_decap_8
XFILLER_1_786 VPWR VGND sg13g2_decap_8
XFILLER_37_908 VPWR VGND sg13g2_decap_8
XFILLER_17_632 VPWR VGND sg13g2_decap_8
XFILLER_29_481 VPWR VGND sg13g2_decap_8
XFILLER_45_974 VPWR VGND sg13g2_decap_8
XFILLER_44_484 VPWR VGND sg13g2_decap_8
XFILLER_32_602 VPWR VGND sg13g2_decap_8
XFILLER_20_819 VPWR VGND sg13g2_decap_8
XFILLER_32_679 VPWR VGND sg13g2_decap_8
XFILLER_13_893 VPWR VGND sg13g2_decap_8
X_2740_ _0265_ VPWR _0269_ VGND _2056_ _0268_ sg13g2_o21ai_1
XFILLER_9_886 VPWR VGND sg13g2_decap_8
X_2671_ _0205_ sap_3_inst.alu_flags\[3\] _1902_ VPWR VGND sg13g2_nand2_1
X_4341_ mem_ram_we net25 VPWR VGND sg13g2_buf_1
X_4272_ net811 VGND VPWR _0129_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[7\]
+ clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3223_ _1633_ VPWR _0694_ VGND _0692_ _0693_ sg13g2_o21ai_1
XFILLER_39_201 VPWR VGND sg13g2_fill_1
XFILLER_39_223 VPWR VGND sg13g2_fill_2
X_3154_ net756 net718 _0627_ VPWR VGND sg13g2_nor2_1
X_3085_ _0355_ _0572_ _0582_ VPWR VGND sg13g2_nor2_1
X_2105_ VPWR _1523_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[0\]
+ VGND sg13g2_inv_1
XFILLER_36_974 VPWR VGND sg13g2_decap_8
XFILLER_23_613 VPWR VGND sg13g2_decap_8
XFILLER_22_156 VPWR VGND sg13g2_fill_1
X_3987_ _0154_ VPWR _1363_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[0\]
+ _1344_ sg13g2_o21ai_1
X_2938_ _0439_ _0438_ VPWR VGND _0437_ sg13g2_nand2b_2
X_2869_ _0372_ net703 sap_3_inst.alu_inst.act\[1\] VPWR VGND sg13g2_nand2b_1
Xfanout810 net812 net810 VPWR VGND sg13g2_buf_8
Xfanout821 net825 net821 VPWR VGND sg13g2_buf_8
Xfanout832 net836 net832 VPWR VGND sg13g2_buf_8
XFILLER_46_727 VPWR VGND sg13g2_decap_8
XFILLER_27_952 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_42_933 VPWR VGND sg13g2_decap_8
XFILLER_14_646 VPWR VGND sg13g2_decap_8
XFILLER_26_495 VPWR VGND sg13g2_decap_8
XFILLER_9_138 VPWR VGND sg13g2_fill_2
XFILLER_10_863 VPWR VGND sg13g2_decap_8
XFILLER_22_690 VPWR VGND sg13g2_decap_8
XFILLER_6_834 VPWR VGND sg13g2_decap_8
XFILLER_49_510 VPWR VGND sg13g2_decap_8
XFILLER_1_583 VPWR VGND sg13g2_decap_8
XFILLER_3_1008 VPWR VGND sg13g2_decap_8
XFILLER_37_705 VPWR VGND sg13g2_decap_8
XFILLER_49_587 VPWR VGND sg13g2_decap_8
XFILLER_18_963 VPWR VGND sg13g2_decap_8
XFILLER_45_771 VPWR VGND sg13g2_decap_8
XFILLER_33_911 VPWR VGND sg13g2_decap_8
X_3910_ net647 VPWR _1297_ VGND net586 _0979_ sg13g2_o21ai_1
XFILLER_20_616 VPWR VGND sg13g2_decap_8
X_3841_ VPWR VGND _0719_ _1055_ _1247_ _1245_ _1248_ _1246_ sg13g2_a221oi_1
XFILLER_33_988 VPWR VGND sg13g2_decap_8
X_3772_ _1198_ VPWR _0104_ VGND _1202_ _1203_ sg13g2_o21ai_1
XFILLER_13_690 VPWR VGND sg13g2_decap_8
X_2723_ VGND VPWR _1899_ _0252_ _0253_ _0251_ sg13g2_a21oi_1
XFILLER_8_171 VPWR VGND sg13g2_fill_1
XFILLER_9_683 VPWR VGND sg13g2_decap_8
X_2654_ _1809_ net626 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[3\]
+ _2061_ VPWR VGND sg13g2_nand3_1
X_2585_ _1605_ net725 _1994_ VPWR VGND sg13g2_nor2_1
X_4324_ net823 VGND VPWR _0181_ sap_3_inst.alu_inst.act\[4\] clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4255_ net811 VGND VPWR _0112_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[6\]
+ clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4186_ net821 VGND VPWR _0043_ sap_3_inst.out\[2\] clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3206_ _1652_ _1666_ _1644_ _0677_ VPWR VGND sg13g2_nand3_1
X_3137_ _0619_ sap_3_inst.alu_inst.tmp\[5\] net700 VPWR VGND sg13g2_nand2_1
XFILLER_27_215 VPWR VGND sg13g2_fill_1
X_3068_ _0566_ _0564_ _0565_ net598 net776 VPWR VGND sg13g2_a22oi_1
XFILLER_36_771 VPWR VGND sg13g2_decap_8
XFILLER_24_955 VPWR VGND sg13g2_decap_8
XFILLER_11_649 VPWR VGND sg13g2_decap_8
XFILLER_23_487 VPWR VGND sg13g2_decap_8
XFILLER_6_119 VPWR VGND sg13g2_fill_1
XFILLER_12_33 VPWR VGND sg13g2_fill_2
XFILLER_3_826 VPWR VGND sg13g2_decap_8
Xfanout651 _0759_ net651 VPWR VGND sg13g2_buf_8
Xfanout640 _0765_ net640 VPWR VGND sg13g2_buf_8
Xfanout684 net685 net684 VPWR VGND sg13g2_buf_8
Xfanout673 net674 net673 VPWR VGND sg13g2_buf_8
Xfanout662 _0713_ net662 VPWR VGND sg13g2_buf_8
XFILLER_46_524 VPWR VGND sg13g2_decap_8
Xfanout695 _1899_ net695 VPWR VGND sg13g2_buf_8
XFILLER_19_749 VPWR VGND sg13g2_decap_8
XFILLER_42_730 VPWR VGND sg13g2_decap_8
XFILLER_15_966 VPWR VGND sg13g2_decap_8
XFILLER_18_1005 VPWR VGND sg13g2_decap_8
XFILLER_30_903 VPWR VGND sg13g2_decap_8
XFILLER_41_284 VPWR VGND sg13g2_fill_1
XFILLER_10_660 VPWR VGND sg13g2_decap_8
XFILLER_6_631 VPWR VGND sg13g2_decap_8
X_2370_ _1704_ _1730_ _1772_ _1786_ _1787_ VPWR VGND sg13g2_nor4_1
XFILLER_1_380 VPWR VGND sg13g2_fill_1
X_4040_ VGND VPWR _1404_ _1409_ _1411_ _1410_ sg13g2_a21oi_1
XFILLER_49_384 VPWR VGND sg13g2_decap_8
XFILLER_37_502 VPWR VGND sg13g2_decap_8
XFILLER_18_760 VPWR VGND sg13g2_decap_8
XFILLER_37_579 VPWR VGND sg13g2_decap_8
XFILLER_33_785 VPWR VGND sg13g2_decap_8
XFILLER_21_958 VPWR VGND sg13g2_decap_8
X_3824_ _0124_ _1236_ _1065_ net635 _1503_ VPWR VGND sg13g2_a22oi_1
X_3755_ _1189_ VPWR _1190_ VGND _1991_ net602 sg13g2_o21ai_1
XFILLER_9_480 VPWR VGND sg13g2_decap_8
X_3686_ _1027_ _1134_ _1135_ VPWR VGND sg13g2_nor2_1
X_2706_ _0237_ sap_3_inst.alu_flags\[2\] _2057_ VPWR VGND sg13g2_nand2_1
X_2637_ _2046_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[1\] net623
+ VPWR VGND sg13g2_nand2_1
X_2568_ _1969_ _1978_ _1979_ VPWR VGND _1768_ sg13g2_nand3b_1
X_2499_ net752 _1628_ net721 _1915_ VPWR VGND sg13g2_nor3_2
X_4307_ net834 VGND VPWR _0164_ sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[3\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_1
X_4238_ net830 VGND VPWR _0095_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[5\]
+ clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4169_ net807 VGND VPWR _0002_ sap_3_inst.controller_inst.stage\[1\] net41 sg13g2_dfrbpq_2
XFILLER_28_568 VPWR VGND sg13g2_decap_8
XFILLER_43_549 VPWR VGND sg13g2_decap_8
XFILLER_24_752 VPWR VGND sg13g2_decap_8
XFILLER_12_947 VPWR VGND sg13g2_decap_8
XFILLER_23_295 VPWR VGND sg13g2_decap_4
XFILLER_20_980 VPWR VGND sg13g2_decap_8
XFILLER_3_623 VPWR VGND sg13g2_decap_8
XFILLER_47_844 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_4
XFILLER_19_546 VPWR VGND sg13g2_decap_8
XFILLER_46_398 VPWR VGND sg13g2_decap_8
XFILLER_34_549 VPWR VGND sg13g2_decap_8
XFILLER_15_763 VPWR VGND sg13g2_decap_8
XFILLER_9_34 VPWR VGND sg13g2_fill_1
XFILLER_30_700 VPWR VGND sg13g2_decap_8
XFILLER_30_777 VPWR VGND sg13g2_decap_8
XFILLER_31_1013 VPWR VGND sg13g2_decap_8
XFILLER_7_940 VPWR VGND sg13g2_decap_8
X_3540_ _1006_ _0978_ _0990_ VPWR VGND sg13g2_xnor2_1
X_3471_ _0936_ _0937_ _0935_ _0939_ VPWR VGND _0938_ sg13g2_nand4_1
X_2422_ _1729_ VPWR _1839_ VGND net726 net733 sg13g2_o21ai_1
X_2353_ net727 _1769_ _1770_ VPWR VGND sg13g2_nor2_1
X_4023_ _1395_ _1340_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[4\]
+ net796 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[4\] VPWR VGND sg13g2_a22oi_1
X_2284_ VGND VPWR net724 _1673_ _1701_ _1700_ sg13g2_a21oi_1
XFILLER_38_811 VPWR VGND sg13g2_decap_8
XFILLER_38_888 VPWR VGND sg13g2_decap_8
XFILLER_25_527 VPWR VGND sg13g2_decap_8
XFILLER_33_582 VPWR VGND sg13g2_decap_8
XFILLER_21_755 VPWR VGND sg13g2_decap_8
X_3807_ net658 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[3\] _1226_
+ _0117_ VPWR VGND sg13g2_a21o_1
X_3738_ _1176_ _1174_ _1175_ net655 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[1\]
+ VPWR VGND sg13g2_a22oi_1
X_3669_ _1120_ net609 _0979_ VPWR VGND sg13g2_nand2_1
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_48_619 VPWR VGND sg13g2_decap_8
XFILLER_28_310 VPWR VGND sg13g2_fill_2
XFILLER_29_866 VPWR VGND sg13g2_decap_8
XFILLER_16_527 VPWR VGND sg13g2_decap_8
XFILLER_44_869 VPWR VGND sg13g2_decap_8
XFILLER_12_744 VPWR VGND sg13g2_decap_8
XFILLER_15_1008 VPWR VGND sg13g2_decap_8
XFILLER_8_759 VPWR VGND sg13g2_decap_8
XFILLER_7_236 VPWR VGND sg13g2_fill_2
XFILLER_4_921 VPWR VGND sg13g2_decap_8
XFILLER_4_998 VPWR VGND sg13g2_decap_8
XFILLER_3_497 VPWR VGND sg13g2_decap_8
XFILLER_47_641 VPWR VGND sg13g2_decap_8
XFILLER_22_508 VPWR VGND sg13g2_decap_8
XFILLER_35_869 VPWR VGND sg13g2_decap_8
X_2971_ VGND VPWR _0454_ _0469_ _0471_ _0468_ sg13g2_a21oi_1
XFILLER_15_560 VPWR VGND sg13g2_decap_8
XFILLER_30_574 VPWR VGND sg13g2_decap_8
X_3523_ _0987_ _0988_ _0986_ _0989_ VPWR VGND sg13g2_nand3_1
X_3454_ _0923_ _0836_ _0847_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_0 VPWR VGND sg13g2_fill_1
X_2405_ net759 _1762_ _1822_ VPWR VGND sg13g2_and2_1
X_3385_ net612 _0855_ _0856_ VPWR VGND sg13g2_nor2_1
X_2336_ _1753_ net725 _1693_ VPWR VGND sg13g2_nand2_1
XFILLER_29_107 VPWR VGND sg13g2_fill_1
X_2267_ sap_3_inst.controller_inst.stage\[0\] _1683_ _1684_ VPWR VGND sg13g2_nor2_2
XFILLER_26_803 VPWR VGND sg13g2_decap_8
X_4006_ _1374_ _1378_ _1373_ _1380_ VPWR VGND _1379_ sg13g2_nand4_1
X_2198_ VGND VPWR _1608_ _1614_ _1615_ _1606_ sg13g2_a21oi_1
XFILLER_38_685 VPWR VGND sg13g2_decap_8
XFILLER_41_817 VPWR VGND sg13g2_decap_8
XFILLER_13_508 VPWR VGND sg13g2_decap_8
XFILLER_21_552 VPWR VGND sg13g2_decap_8
XFILLER_0_412 VPWR VGND sg13g2_fill_1
XFILLER_1_968 VPWR VGND sg13g2_decap_8
XFILLER_48_416 VPWR VGND sg13g2_decap_8
Xhold20 u_ser.shadow_reg\[4\] VPWR VGND net67 sg13g2_dlygate4sd3_1
Xhold31 sap_3_inst.reg_file_inst.array_serializer_inst.state\[0\] VPWR VGND net78
+ sg13g2_dlygate4sd3_1
XFILLER_17_814 VPWR VGND sg13g2_decap_8
XFILLER_29_663 VPWR VGND sg13g2_decap_8
XFILLER_44_666 VPWR VGND sg13g2_decap_8
XFILLER_25_891 VPWR VGND sg13g2_decap_8
XFILLER_12_541 VPWR VGND sg13g2_decap_8
XFILLER_8_556 VPWR VGND sg13g2_decap_8
XFILLER_4_795 VPWR VGND sg13g2_decap_8
X_3170_ _0633_ _0634_ _0637_ _0640_ _0641_ VPWR VGND sg13g2_nor4_1
X_2121_ _1539_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[6\] VPWR
+ VGND sg13g2_inv_2
XFILLER_48_983 VPWR VGND sg13g2_decap_8
XFILLER_35_666 VPWR VGND sg13g2_decap_8
XFILLER_16_891 VPWR VGND sg13g2_decap_8
X_2954_ _0455_ net783 net708 VPWR VGND sg13g2_xnor2_1
X_2885_ _2000_ VPWR _0388_ VGND net792 _0386_ sg13g2_o21ai_1
XFILLER_31_894 VPWR VGND sg13g2_decap_8
X_3506_ VGND VPWR _0802_ _0861_ _0973_ net585 sg13g2_a21oi_1
X_3437_ _0906_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[2\] net596
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_1023 VPWR VGND sg13g2_decap_4
X_3368_ _0839_ net677 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[1\]
+ net683 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2319_ VGND VPWR _1554_ _1679_ _1736_ _1735_ sg13g2_a21oi_1
XFILLER_46_909 VPWR VGND sg13g2_decap_8
X_3299_ _0768_ _0769_ _0770_ VPWR VGND sg13g2_and2_1
XFILLER_26_600 VPWR VGND sg13g2_decap_8
XFILLER_38_482 VPWR VGND sg13g2_decap_8
XFILLER_41_614 VPWR VGND sg13g2_decap_8
XFILLER_14_828 VPWR VGND sg13g2_decap_8
XFILLER_26_677 VPWR VGND sg13g2_decap_8
XFILLER_40_168 VPWR VGND sg13g2_fill_2
XFILLER_40_146 VPWR VGND sg13g2_fill_2
XFILLER_22_872 VPWR VGND sg13g2_decap_8
XFILLER_31_76 VPWR VGND sg13g2_fill_2
XFILLER_5_548 VPWR VGND sg13g2_decap_8
Xoutput21 net21 uio_out[4] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_oe[1] VPWR VGND sg13g2_buf_1
XFILLER_1_765 VPWR VGND sg13g2_decap_8
XFILLER_49_769 VPWR VGND sg13g2_decap_8
XFILLER_17_611 VPWR VGND sg13g2_decap_8
XFILLER_45_953 VPWR VGND sg13g2_decap_8
XFILLER_44_463 VPWR VGND sg13g2_decap_8
XFILLER_17_688 VPWR VGND sg13g2_decap_8
XFILLER_16_198 VPWR VGND sg13g2_fill_1
XFILLER_31_102 VPWR VGND sg13g2_fill_2
XFILLER_32_658 VPWR VGND sg13g2_decap_8
XFILLER_13_872 VPWR VGND sg13g2_decap_8
XFILLER_12_382 VPWR VGND sg13g2_fill_2
XFILLER_9_865 VPWR VGND sg13g2_decap_8
X_2670_ net577 VPWR _0204_ VGND _0199_ _0203_ sg13g2_o21ai_1
X_4271_ net811 VGND VPWR _0128_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[6\]
+ clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_4_592 VPWR VGND sg13g2_decap_8
X_3222_ _1650_ _1652_ _1640_ _0693_ VPWR VGND _1691_ sg13g2_nand4_1
X_3153_ VGND VPWR net717 net569 _0063_ _0626_ sg13g2_a21oi_1
X_2104_ VPWR _1522_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[0\]
+ VGND sg13g2_inv_1
XFILLER_48_780 VPWR VGND sg13g2_decap_8
X_3084_ _0581_ _0361_ _0570_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_953 VPWR VGND sg13g2_decap_8
XFILLER_23_669 VPWR VGND sg13g2_decap_8
X_3986_ _1359_ _1361_ _1362_ VPWR VGND sg13g2_nor2_1
X_2937_ _0438_ net784 sap_3_inst.alu_inst.tmp\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_31_691 VPWR VGND sg13g2_decap_8
X_2868_ VGND VPWR _1508_ net599 _0033_ _0371_ sg13g2_a21oi_1
X_2799_ net714 _1697_ _1704_ _1802_ _0313_ VPWR VGND sg13g2_nor4_1
Xfanout800 u_ser.bit_pos\[0\] net800 VPWR VGND sg13g2_buf_2
Xfanout811 net812 net811 VPWR VGND sg13g2_buf_8
Xfanout822 net825 net822 VPWR VGND sg13g2_buf_8
Xfanout833 net834 net833 VPWR VGND sg13g2_buf_8
XFILLER_46_706 VPWR VGND sg13g2_decap_8
XFILLER_27_931 VPWR VGND sg13g2_decap_8
XFILLER_42_912 VPWR VGND sg13g2_decap_8
XFILLER_26_474 VPWR VGND sg13g2_decap_8
XFILLER_14_625 VPWR VGND sg13g2_decap_8
XFILLER_42_989 VPWR VGND sg13g2_decap_8
XFILLER_41_488 VPWR VGND sg13g2_decap_8
XFILLER_9_128 VPWR VGND sg13g2_fill_1
XFILLER_10_842 VPWR VGND sg13g2_decap_8
XFILLER_6_813 VPWR VGND sg13g2_decap_8
XFILLER_1_562 VPWR VGND sg13g2_decap_8
XFILLER_3_58 VPWR VGND sg13g2_fill_1
XFILLER_49_566 VPWR VGND sg13g2_decap_8
XFILLER_18_942 VPWR VGND sg13g2_decap_8
XFILLER_36_227 VPWR VGND sg13g2_fill_2
XFILLER_45_750 VPWR VGND sg13g2_decap_8
XFILLER_17_485 VPWR VGND sg13g2_decap_8
X_3840_ _1247_ _0301_ _0730_ VPWR VGND sg13g2_nand2_1
XFILLER_33_967 VPWR VGND sg13g2_decap_8
X_3771_ VGND VPWR _1204_ _1021_ net586 sg13g2_or2_1
XFILLER_34_1011 VPWR VGND sg13g2_decap_8
XFILLER_9_662 VPWR VGND sg13g2_decap_8
X_2722_ _0252_ sap_3_inst.alu_flags\[0\] _1902_ VPWR VGND sg13g2_nand2_1
X_2653_ net697 net626 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[3\]
+ _2060_ VPWR VGND sg13g2_nand3_1
X_2584_ _1993_ _1598_ _1612_ VPWR VGND sg13g2_nand2_1
X_4323_ net825 VGND VPWR _0180_ sap_3_inst.alu_inst.act\[3\] clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4254_ net830 VGND VPWR _0111_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[5\]
+ clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3205_ VGND VPWR net727 net720 _0676_ _1691_ sg13g2_a21oi_1
X_4185_ net821 VGND VPWR _0042_ sap_3_inst.out\[1\] clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3136_ _0618_ VPWR _0054_ VGND _1991_ net701 sg13g2_o21ai_1
X_3067_ VGND VPWR _1941_ net693 _0565_ net598 sg13g2_a21oi_1
XFILLER_36_750 VPWR VGND sg13g2_decap_8
XFILLER_24_934 VPWR VGND sg13g2_decap_8
XFILLER_23_466 VPWR VGND sg13g2_decap_8
XFILLER_11_628 VPWR VGND sg13g2_decap_8
X_3969_ _1345_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[0\] VPWR
+ VGND sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[1\] sg13g2_nand2b_2
XFILLER_3_805 VPWR VGND sg13g2_decap_8
Xfanout630 net633 net630 VPWR VGND sg13g2_buf_8
Xfanout641 _0762_ net641 VPWR VGND sg13g2_buf_8
Xfanout663 net664 net663 VPWR VGND sg13g2_buf_8
Xfanout674 _0757_ net674 VPWR VGND sg13g2_buf_8
Xfanout685 _0747_ net685 VPWR VGND sg13g2_buf_8
Xfanout652 net654 net652 VPWR VGND sg13g2_buf_8
XFILLER_46_503 VPWR VGND sg13g2_decap_8
XFILLER_19_728 VPWR VGND sg13g2_decap_8
Xfanout696 _1792_ net696 VPWR VGND sg13g2_buf_8
XFILLER_37_86 VPWR VGND sg13g2_fill_2
XFILLER_15_945 VPWR VGND sg13g2_decap_8
XFILLER_33_219 VPWR VGND sg13g2_fill_2
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_26_293 VPWR VGND sg13g2_fill_2
XFILLER_42_786 VPWR VGND sg13g2_decap_8
XFILLER_14_499 VPWR VGND sg13g2_decap_8
XFILLER_30_959 VPWR VGND sg13g2_decap_8
XFILLER_6_610 VPWR VGND sg13g2_decap_8
XFILLER_6_687 VPWR VGND sg13g2_decap_8
XFILLER_5_153 VPWR VGND sg13g2_fill_1
X_4152__10 VPWR net44 clknet_leaf_0_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
XFILLER_49_363 VPWR VGND sg13g2_decap_8
Xclkbuf_5_1__f_sap_3_inst.alu_inst.clk_regs clknet_4_0_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_37_558 VPWR VGND sg13g2_decap_8
XFILLER_25_709 VPWR VGND sg13g2_decap_8
XFILLER_33_764 VPWR VGND sg13g2_decap_8
X_3823_ _1066_ net634 _1236_ VPWR VGND sg13g2_nor2_1
XFILLER_21_937 VPWR VGND sg13g2_decap_8
X_3754_ VGND VPWR net13 net602 _1189_ net593 sg13g2_a21oi_1
X_3685_ net592 VPWR _1134_ VGND net638 _1028_ sg13g2_o21ai_1
X_2705_ _0235_ VPWR _0236_ VGND _1916_ net19 sg13g2_o21ai_1
X_2636_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[1\] net620
+ net629 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[1\] _2045_ net713
+ sg13g2_a221oi_1
X_2567_ _1972_ _1974_ _1970_ _1978_ VPWR VGND _1977_ sg13g2_nand4_1
XFILLER_0_819 VPWR VGND sg13g2_decap_8
X_2498_ net24 _1914_ VPWR VGND sg13g2_inv_4
X_4306_ net833 VGND VPWR _0163_ sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[2\]
+ clknet_3_3__leaf_clk sg13g2_dfrbpq_1
X_4237_ net814 VGND VPWR _0094_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[4\]
+ clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4168_ net804 VGND VPWR _0001_ sap_3_inst.controller_inst.stage\[0\] net40 sg13g2_dfrbpq_2
XFILLER_28_547 VPWR VGND sg13g2_decap_8
X_3119_ VGND VPWR _0350_ _0600_ _0607_ _0606_ sg13g2_a21oi_1
X_4099_ _1509_ _0480_ net698 _1455_ VPWR VGND sg13g2_mux2_1
XFILLER_16_709 VPWR VGND sg13g2_decap_8
XFILLER_43_528 VPWR VGND sg13g2_decap_8
XFILLER_24_731 VPWR VGND sg13g2_decap_8
XFILLER_12_926 VPWR VGND sg13g2_decap_8
XFILLER_3_602 VPWR VGND sg13g2_decap_8
XFILLER_2_101 VPWR VGND sg13g2_decap_4
XFILLER_3_679 VPWR VGND sg13g2_decap_8
XFILLER_47_823 VPWR VGND sg13g2_decap_8
XFILLER_19_525 VPWR VGND sg13g2_decap_8
XFILLER_46_377 VPWR VGND sg13g2_decap_8
XFILLER_34_528 VPWR VGND sg13g2_decap_8
XFILLER_15_742 VPWR VGND sg13g2_decap_8
XFILLER_42_583 VPWR VGND sg13g2_decap_8
XFILLER_9_57 VPWR VGND sg13g2_fill_1
XFILLER_30_756 VPWR VGND sg13g2_decap_8
XFILLER_11_992 VPWR VGND sg13g2_decap_8
XFILLER_7_996 VPWR VGND sg13g2_decap_8
XFILLER_6_484 VPWR VGND sg13g2_decap_8
X_3470_ _0938_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[3\] _0763_
+ VPWR VGND sg13g2_nand2_1
X_2421_ net728 _1600_ _1837_ _1838_ VPWR VGND sg13g2_nor3_1
X_2352_ _1769_ net765 _1616_ VPWR VGND sg13g2_nand2_1
XFILLER_9_1026 VPWR VGND sg13g2_fill_2
X_2283_ _1561_ _1572_ _1557_ _1700_ VPWR VGND sg13g2_nand3_1
X_4022_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[4\] _1347_
+ _1394_ net794 sg13g2_a21oi_1
XFILLER_25_506 VPWR VGND sg13g2_decap_8
XFILLER_37_366 VPWR VGND sg13g2_fill_1
XFILLER_38_867 VPWR VGND sg13g2_decap_8
XFILLER_37_377 VPWR VGND sg13g2_fill_2
XFILLER_33_561 VPWR VGND sg13g2_decap_8
XFILLER_21_734 VPWR VGND sg13g2_decap_8
X_3806_ VGND VPWR _1070_ _1183_ _1226_ net658 sg13g2_a21oi_1
XFILLER_20_288 VPWR VGND sg13g2_decap_8
X_3737_ VGND VPWR net607 _0900_ _1175_ net655 sg13g2_a21oi_1
X_3668_ net609 _0979_ _1119_ VPWR VGND sg13g2_and2_1
X_3599_ net583 _1060_ _1061_ VPWR VGND sg13g2_nor2_1
X_2619_ net667 net627 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[1\]
+ _2028_ VPWR VGND sg13g2_nand3_1
XFILLER_0_616 VPWR VGND sg13g2_decap_8
XFILLER_29_845 VPWR VGND sg13g2_decap_8
XFILLER_16_506 VPWR VGND sg13g2_decap_8
XFILLER_18_55 VPWR VGND sg13g2_fill_1
XFILLER_44_848 VPWR VGND sg13g2_decap_8
XFILLER_31_509 VPWR VGND sg13g2_decap_8
XFILLER_12_723 VPWR VGND sg13g2_decap_8
XFILLER_8_738 VPWR VGND sg13g2_decap_8
XFILLER_4_900 VPWR VGND sg13g2_decap_8
XFILLER_4_977 VPWR VGND sg13g2_decap_8
XFILLER_3_476 VPWR VGND sg13g2_decap_8
XFILLER_47_620 VPWR VGND sg13g2_decap_8
XFILLER_47_697 VPWR VGND sg13g2_decap_8
XFILLER_35_848 VPWR VGND sg13g2_decap_8
X_2970_ _0468_ _0469_ _0454_ _0470_ VPWR VGND sg13g2_nand3_1
XFILLER_43_892 VPWR VGND sg13g2_decap_8
XFILLER_30_553 VPWR VGND sg13g2_decap_8
XFILLER_7_793 VPWR VGND sg13g2_decap_8
X_3522_ _0988_ net640 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[5\]
+ net642 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[5\] VPWR VGND sg13g2_a22oi_1
X_3453_ _0922_ _0875_ net11 VPWR VGND sg13g2_nand2b_1
X_2404_ VGND VPWR net769 _1750_ _1821_ _1748_ sg13g2_a21oi_1
X_3384_ _0855_ _0854_ VPWR VGND _0853_ sg13g2_nand2b_2
X_2335_ _1752_ net732 _1553_ net736 net738 VPWR VGND sg13g2_a22oi_1
X_2266_ sap_3_inst.controller_inst.stage\[3\] net746 _1683_ VPWR VGND net745 sg13g2_nand3b_1
X_2197_ _1614_ net729 net725 VPWR VGND sg13g2_nand2_1
X_4005_ _1379_ _1350_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[2\]
+ _1346_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_38_664 VPWR VGND sg13g2_decap_8
XFILLER_26_859 VPWR VGND sg13g2_decap_8
XFILLER_40_306 VPWR VGND sg13g2_fill_1
XFILLER_21_531 VPWR VGND sg13g2_decap_8
XFILLER_34_892 VPWR VGND sg13g2_decap_8
XFILLER_1_947 VPWR VGND sg13g2_decap_8
Xhold10 u_ser.shadow_reg\[7\] VPWR VGND net57 sg13g2_dlygate4sd3_1
Xhold21 u_ser.state\[0\] VPWR VGND net68 sg13g2_dlygate4sd3_1
Xhold32 sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[0\] VPWR VGND net79
+ sg13g2_dlygate4sd3_1
XFILLER_29_642 VPWR VGND sg13g2_decap_8
XFILLER_44_645 VPWR VGND sg13g2_decap_8
XFILLER_25_870 VPWR VGND sg13g2_decap_8
XFILLER_12_520 VPWR VGND sg13g2_decap_8
XFILLER_40_884 VPWR VGND sg13g2_decap_8
XFILLER_8_535 VPWR VGND sg13g2_decap_8
XFILLER_12_597 VPWR VGND sg13g2_decap_8
XFILLER_4_774 VPWR VGND sg13g2_decap_8
X_2120_ VPWR _1538_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[5\]
+ VGND sg13g2_inv_1
XFILLER_0_980 VPWR VGND sg13g2_decap_8
XFILLER_48_962 VPWR VGND sg13g2_decap_8
XFILLER_19_174 VPWR VGND sg13g2_fill_1
XFILLER_47_494 VPWR VGND sg13g2_decap_8
XFILLER_35_645 VPWR VGND sg13g2_decap_8
XFILLER_16_870 VPWR VGND sg13g2_decap_8
X_2953_ _0454_ net783 net708 VPWR VGND sg13g2_nand2_1
XFILLER_37_1020 VPWR VGND sg13g2_decap_8
XFILLER_31_873 VPWR VGND sg13g2_decap_8
X_2884_ _0387_ net792 _0386_ VPWR VGND sg13g2_nand2_1
X_3505_ net21 net13 _0875_ _0972_ VPWR VGND sg13g2_mux2_1
XFILLER_7_590 VPWR VGND sg13g2_decap_8
XFILLER_44_1002 VPWR VGND sg13g2_decap_8
X_3436_ _0067_ _0896_ _0905_ net596 _1510_ VPWR VGND sg13g2_a22oi_1
X_3367_ _0838_ net680 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[1\]
+ net688 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2318_ _1735_ _1630_ _1683_ VPWR VGND sg13g2_nand2_1
X_3298_ _0769_ net664 sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[0\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_39_984 VPWR VGND sg13g2_decap_8
X_2249_ VGND VPWR _1666_ net749 _1576_ sg13g2_or2_1
XFILLER_26_656 VPWR VGND sg13g2_decap_8
XFILLER_14_807 VPWR VGND sg13g2_decap_8
XFILLER_22_851 VPWR VGND sg13g2_decap_8
XFILLER_5_527 VPWR VGND sg13g2_decap_8
Xoutput22 net22 uio_out[5] VPWR VGND sg13g2_buf_1
Xoutput9 net9 uio_oe[0] VPWR VGND sg13g2_buf_1
Xoutput11 net11 uio_oe[2] VPWR VGND sg13g2_buf_1
XFILLER_1_744 VPWR VGND sg13g2_decap_8
XFILLER_49_748 VPWR VGND sg13g2_decap_8
XFILLER_45_932 VPWR VGND sg13g2_decap_8
XFILLER_44_442 VPWR VGND sg13g2_decap_8
XFILLER_17_667 VPWR VGND sg13g2_decap_8
XFILLER_32_637 VPWR VGND sg13g2_decap_8
XFILLER_13_851 VPWR VGND sg13g2_decap_8
XFILLER_40_681 VPWR VGND sg13g2_decap_8
XFILLER_9_844 VPWR VGND sg13g2_decap_8
X_4270_ net815 VGND VPWR _0127_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[5\]
+ clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_4_571 VPWR VGND sg13g2_decap_8
X_3221_ _1666_ _1700_ _1644_ _0692_ VPWR VGND sg13g2_nand3_1
X_3152_ net758 net717 _0626_ VPWR VGND sg13g2_nor2_1
X_2103_ VPWR _1521_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[0\]
+ VGND sg13g2_inv_1
XFILLER_39_247 VPWR VGND sg13g2_fill_1
X_3083_ _0580_ _0358_ net691 net692 net776 VPWR VGND sg13g2_a22oi_1
XFILLER_35_420 VPWR VGND sg13g2_fill_1
XFILLER_36_932 VPWR VGND sg13g2_decap_8
XFILLER_23_648 VPWR VGND sg13g2_decap_8
X_3985_ _1361_ _1355_ _1360_ VPWR VGND sg13g2_nand2_1
X_2936_ net784 sap_3_inst.alu_inst.tmp\[3\] _0437_ VPWR VGND sg13g2_nor2_1
XFILLER_31_670 VPWR VGND sg13g2_decap_8
X_2867_ VPWR VGND _0370_ net599 _0369_ net31 _0371_ net694 sg13g2_a221oi_1
X_2798_ _0312_ _1744_ _0311_ VPWR VGND sg13g2_nand2_1
XFILLER_2_519 VPWR VGND sg13g2_decap_8
Xclkbuf_1_0__f_clk_div_out clknet_0_clk_div_out clknet_1_0__leaf_clk_div_out VPWR
+ VGND sg13g2_buf_8
Xfanout812 net813 net812 VPWR VGND sg13g2_buf_8
Xfanout801 sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[3\] net801 VPWR
+ VGND sg13g2_buf_8
Xfanout823 net825 net823 VPWR VGND sg13g2_buf_8
X_3419_ _1518_ net637 _0889_ VPWR VGND sg13g2_nor2_1
Xfanout834 net835 net834 VPWR VGND sg13g2_buf_8
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_39_781 VPWR VGND sg13g2_decap_8
XFILLER_14_604 VPWR VGND sg13g2_decap_8
XFILLER_26_453 VPWR VGND sg13g2_decap_8
XFILLER_27_987 VPWR VGND sg13g2_decap_8
XFILLER_42_968 VPWR VGND sg13g2_decap_8
XFILLER_41_467 VPWR VGND sg13g2_decap_8
XFILLER_10_821 VPWR VGND sg13g2_decap_8
XFILLER_6_869 VPWR VGND sg13g2_decap_8
XFILLER_10_898 VPWR VGND sg13g2_decap_8
XFILLER_1_541 VPWR VGND sg13g2_decap_8
XFILLER_3_48 VPWR VGND sg13g2_fill_2
XFILLER_49_545 VPWR VGND sg13g2_decap_8
XFILLER_18_921 VPWR VGND sg13g2_decap_8
XFILLER_18_998 VPWR VGND sg13g2_decap_8
XFILLER_33_946 VPWR VGND sg13g2_decap_8
X_3770_ _1203_ net676 _1132_ VPWR VGND sg13g2_nand2_1
XFILLER_9_641 VPWR VGND sg13g2_decap_8
X_2721_ net793 net695 _0251_ VPWR VGND sg13g2_nor2_1
XFILLER_8_140 VPWR VGND sg13g2_fill_2
X_2652_ _2059_ _1497_ net632 VPWR VGND sg13g2_nand2_1
X_2583_ VGND VPWR net710 _1991_ _0029_ _1992_ sg13g2_a21oi_1
XFILLER_5_891 VPWR VGND sg13g2_decap_8
X_4322_ net824 VGND VPWR _0179_ sap_3_inst.alu_inst.act\[2\] clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4253_ net814 VGND VPWR _0110_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[4\]
+ clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3204_ _1670_ _0674_ _1649_ _0675_ VPWR VGND sg13g2_nand3_1
XFILLER_41_1027 VPWR VGND sg13g2_fill_2
X_4184_ net817 VGND VPWR _0041_ sap_3_inst.out\[0\] clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3135_ _0618_ sap_3_inst.alu_inst.tmp\[4\] net700 VPWR VGND sg13g2_nand2_1
XFILLER_28_729 VPWR VGND sg13g2_decap_8
X_3066_ _0564_ _0563_ _0562_ VPWR VGND sg13g2_nand2b_1
XFILLER_24_913 VPWR VGND sg13g2_decap_8
XFILLER_23_445 VPWR VGND sg13g2_decap_8
X_3968_ VGND VPWR _1342_ _1344_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[2\]
+ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[3\] sg13g2_a21oi_2
XFILLER_11_607 VPWR VGND sg13g2_decap_8
X_2919_ _0421_ _0420_ _0344_ _0413_ _0348_ VPWR VGND sg13g2_a22oi_1
X_3899_ _1289_ net659 net648 VPWR VGND sg13g2_nand2_1
XFILLER_2_327 VPWR VGND sg13g2_fill_1
Xfanout631 net632 net631 VPWR VGND sg13g2_buf_8
Xfanout620 _1856_ net620 VPWR VGND sg13g2_buf_8
Xfanout642 _0762_ net642 VPWR VGND sg13g2_buf_8
Xfanout653 net654 net653 VPWR VGND sg13g2_buf_1
Xfanout675 net679 net675 VPWR VGND sg13g2_buf_8
Xfanout664 net665 net664 VPWR VGND sg13g2_buf_8
XFILLER_19_707 VPWR VGND sg13g2_decap_8
Xfanout697 _1792_ net697 VPWR VGND sg13g2_buf_2
Xfanout686 net688 net686 VPWR VGND sg13g2_buf_8
XFILLER_46_559 VPWR VGND sg13g2_decap_8
XFILLER_15_924 VPWR VGND sg13g2_decap_8
XFILLER_27_784 VPWR VGND sg13g2_decap_8
XFILLER_42_765 VPWR VGND sg13g2_decap_8
XFILLER_30_938 VPWR VGND sg13g2_decap_8
XFILLER_10_695 VPWR VGND sg13g2_decap_8
XFILLER_6_666 VPWR VGND sg13g2_decap_8
XFILLER_2_883 VPWR VGND sg13g2_decap_8
XFILLER_49_342 VPWR VGND sg13g2_decap_8
XFILLER_37_537 VPWR VGND sg13g2_decap_8
XFILLER_18_795 VPWR VGND sg13g2_decap_8
XFILLER_33_743 VPWR VGND sg13g2_decap_8
XFILLER_21_916 VPWR VGND sg13g2_decap_8
X_3822_ _0123_ _1235_ _1063_ net635 _1514_ VPWR VGND sg13g2_a22oi_1
X_3753_ net592 VPWR _1188_ VGND _0968_ _1187_ sg13g2_o21ai_1
X_3684_ _1133_ net638 _1132_ VPWR VGND sg13g2_nand2_1
X_2704_ _0235_ _1916_ _0234_ VPWR VGND sg13g2_nand2_1
X_2635_ _2044_ _2041_ _2042_ _2043_ VPWR VGND sg13g2_and3_1
X_2566_ _1971_ _1973_ _1975_ _1976_ _1977_ VPWR VGND sg13g2_and4_1
X_4305_ net833 VGND VPWR _0162_ sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[1\]
+ clknet_3_3__leaf_clk sg13g2_dfrbpq_1
X_2497_ _1905_ _1913_ _1868_ net24 VPWR VGND sg13g2_nand3_1
X_4236_ net830 VGND VPWR _0093_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[3\]
+ clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4167_ net817 VGND VPWR _0028_ sap_3_inst.alu_flags\[1\] net39 sg13g2_dfrbpq_1
X_3118_ _0605_ VPWR _0606_ VGND _0345_ _0602_ sg13g2_o21ai_1
XFILLER_28_526 VPWR VGND sg13g2_decap_8
XFILLER_43_507 VPWR VGND sg13g2_decap_8
X_4098_ _1454_ VPWR _0180_ VGND net578 _1453_ sg13g2_o21ai_1
X_3049_ _0545_ _0542_ _0547_ VPWR VGND sg13g2_xor2_1
XFILLER_24_710 VPWR VGND sg13g2_decap_8
XFILLER_12_905 VPWR VGND sg13g2_decap_8
XFILLER_24_787 VPWR VGND sg13g2_decap_8
Xclkbuf_5_25__f_sap_3_inst.alu_inst.clk_regs clknet_4_12_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_3_658 VPWR VGND sg13g2_decap_8
XFILLER_24_1011 VPWR VGND sg13g2_decap_8
XFILLER_47_802 VPWR VGND sg13g2_decap_8
XFILLER_19_504 VPWR VGND sg13g2_decap_8
XFILLER_47_879 VPWR VGND sg13g2_decap_8
XFILLER_46_356 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_4
XFILLER_34_507 VPWR VGND sg13g2_decap_8
XFILLER_15_721 VPWR VGND sg13g2_decap_8
XFILLER_27_581 VPWR VGND sg13g2_decap_8
Xclkbuf_5_14__f_sap_3_inst.alu_inst.clk_regs clknet_4_7_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_42_562 VPWR VGND sg13g2_decap_8
XFILLER_14_264 VPWR VGND sg13g2_fill_2
XFILLER_9_69 VPWR VGND sg13g2_fill_2
XFILLER_15_798 VPWR VGND sg13g2_decap_8
XFILLER_30_735 VPWR VGND sg13g2_decap_8
XFILLER_11_971 VPWR VGND sg13g2_decap_8
XFILLER_7_975 VPWR VGND sg13g2_decap_8
XFILLER_6_463 VPWR VGND sg13g2_decap_8
XFILLER_10_492 VPWR VGND sg13g2_decap_8
X_2420_ _1837_ net763 net752 VPWR VGND sg13g2_nand2_1
XFILLER_9_1005 VPWR VGND sg13g2_decap_8
X_2351_ _1588_ _1720_ _1578_ _1768_ VPWR VGND _1767_ sg13g2_nand4_1
X_2282_ _1558_ _1562_ _1573_ _1699_ VPWR VGND sg13g2_nor3_2
XFILLER_2_680 VPWR VGND sg13g2_decap_8
X_4021_ _1393_ VPWR _0164_ VGND _1391_ _1392_ sg13g2_o21ai_1
XFILLER_38_846 VPWR VGND sg13g2_decap_8
XFILLER_18_592 VPWR VGND sg13g2_decap_8
XFILLER_33_540 VPWR VGND sg13g2_decap_8
XFILLER_21_713 VPWR VGND sg13g2_decap_8
X_3805_ _1224_ VPWR _0116_ VGND _0929_ _1225_ sg13g2_o21ai_1
X_3736_ _1170_ _1172_ _1149_ _1174_ VPWR VGND _1173_ sg13g2_nand4_1
X_3667_ _0968_ _1117_ _1118_ VPWR VGND sg13g2_nor2_1
X_2618_ net696 net627 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[1\]
+ _2027_ VPWR VGND sg13g2_nand3_1
X_3598_ net588 _0883_ _1060_ VPWR VGND sg13g2_nor2_2
X_2549_ _1962_ net622 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[5\]
+ net632 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4219_ net819 VGND VPWR _0076_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[2\]
+ clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_29_824 VPWR VGND sg13g2_decap_8
XFILLER_44_827 VPWR VGND sg13g2_decap_8
XFILLER_12_702 VPWR VGND sg13g2_decap_8
XFILLER_24_584 VPWR VGND sg13g2_decap_8
XFILLER_8_717 VPWR VGND sg13g2_decap_8
XFILLER_12_779 VPWR VGND sg13g2_decap_8
XFILLER_4_956 VPWR VGND sg13g2_decap_8
XFILLER_3_455 VPWR VGND sg13g2_decap_8
XFILLER_47_676 VPWR VGND sg13g2_decap_8
XFILLER_35_827 VPWR VGND sg13g2_decap_8
XFILLER_28_890 VPWR VGND sg13g2_decap_8
XFILLER_34_337 VPWR VGND sg13g2_fill_2
XFILLER_43_871 VPWR VGND sg13g2_decap_8
XFILLER_15_595 VPWR VGND sg13g2_decap_8
XFILLER_30_532 VPWR VGND sg13g2_decap_8
X_3521_ _0987_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[5\] _0763_
+ VPWR VGND sg13g2_nand2_1
XFILLER_7_772 VPWR VGND sg13g2_decap_8
X_3452_ _0921_ _0227_ net605 VPWR VGND sg13g2_nand2_1
X_2403_ _1813_ VPWR _1820_ VGND _1678_ _1819_ sg13g2_o21ai_1
X_3383_ _0770_ VPWR _0854_ VGND _0780_ _0852_ sg13g2_o21ai_1
X_2334_ _1602_ _1697_ _1748_ _1750_ _1751_ VPWR VGND sg13g2_nor4_1
X_2265_ _1682_ _1580_ _1679_ VPWR VGND sg13g2_nand2_2
X_2196_ _1613_ net738 _1610_ VPWR VGND sg13g2_nand2_2
X_4004_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[2\] _1351_
+ _1378_ net795 sg13g2_a21oi_1
XFILLER_38_643 VPWR VGND sg13g2_decap_8
XFILLER_26_838 VPWR VGND sg13g2_decap_8
X_4145__3 VPWR net37 clknet_leaf_1_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
XFILLER_34_871 VPWR VGND sg13g2_decap_8
XFILLER_21_510 VPWR VGND sg13g2_decap_8
XFILLER_14_1010 VPWR VGND sg13g2_decap_8
XFILLER_21_587 VPWR VGND sg13g2_decap_8
XFILLER_5_709 VPWR VGND sg13g2_decap_8
X_3719_ _1161_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[5\] net582
+ VPWR VGND sg13g2_nand2_1
XFILLER_1_926 VPWR VGND sg13g2_decap_8
Xhold11 u_ser.shadow_reg\[0\] VPWR VGND net58 sg13g2_dlygate4sd3_1
Xhold22 _0195_ VPWR VGND net69 sg13g2_dlygate4sd3_1
XFILLER_0_469 VPWR VGND sg13g2_decap_8
XFILLER_29_66 VPWR VGND sg13g2_fill_2
XFILLER_29_621 VPWR VGND sg13g2_decap_8
XFILLER_21_1014 VPWR VGND sg13g2_decap_8
XFILLER_44_624 VPWR VGND sg13g2_decap_8
XFILLER_16_304 VPWR VGND sg13g2_fill_2
XFILLER_29_698 VPWR VGND sg13g2_decap_8
XFILLER_17_849 VPWR VGND sg13g2_decap_8
XFILLER_32_819 VPWR VGND sg13g2_decap_8
XFILLER_40_863 VPWR VGND sg13g2_decap_8
XFILLER_8_514 VPWR VGND sg13g2_decap_8
XFILLER_12_576 VPWR VGND sg13g2_decap_8
XFILLER_4_753 VPWR VGND sg13g2_decap_8
XFILLER_10_90 VPWR VGND sg13g2_decap_4
XFILLER_48_941 VPWR VGND sg13g2_decap_8
XFILLER_47_473 VPWR VGND sg13g2_decap_8
XFILLER_35_624 VPWR VGND sg13g2_decap_8
XFILLER_22_307 VPWR VGND sg13g2_decap_8
X_2952_ _0453_ _0422_ _0425_ VPWR VGND sg13g2_nand2_1
XFILLER_31_852 VPWR VGND sg13g2_decap_8
X_2883_ net709 net789 _0386_ VPWR VGND sg13g2_xor2_1
XFILLER_30_373 VPWR VGND sg13g2_fill_1
X_3504_ VGND VPWR net663 _0968_ _0971_ _0970_ sg13g2_a21oi_1
X_3435_ net596 _0902_ _0904_ _0905_ VPWR VGND sg13g2_nor3_1
X_3366_ _0690_ _0748_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[1\]
+ _0837_ VPWR VGND sg13g2_nand3_1
X_2317_ VGND VPWR _1732_ _1733_ _1734_ net733 sg13g2_a21oi_1
X_3297_ _0761_ _0764_ _0756_ _0768_ VPWR VGND _0767_ sg13g2_nand4_1
XFILLER_39_963 VPWR VGND sg13g2_decap_8
X_2248_ _1665_ _1637_ net714 VPWR VGND sg13g2_nand2_1
X_2179_ _1596_ net753 _1496_ VPWR VGND sg13g2_nand2_2
XFILLER_26_635 VPWR VGND sg13g2_decap_8
XFILLER_41_649 VPWR VGND sg13g2_decap_8
XFILLER_15_35 VPWR VGND sg13g2_fill_1
XFILLER_15_57 VPWR VGND sg13g2_fill_2
XFILLER_25_178 VPWR VGND sg13g2_fill_2
XFILLER_40_148 VPWR VGND sg13g2_fill_1
XFILLER_22_830 VPWR VGND sg13g2_decap_8
XFILLER_5_506 VPWR VGND sg13g2_decap_8
XFILLER_31_67 VPWR VGND sg13g2_fill_1
Xoutput23 net23 uio_out[6] VPWR VGND sg13g2_buf_1
Xoutput12 net12 uio_oe[3] VPWR VGND sg13g2_buf_1
XFILLER_1_723 VPWR VGND sg13g2_decap_8
XFILLER_49_727 VPWR VGND sg13g2_decap_8
XFILLER_45_911 VPWR VGND sg13g2_decap_8
XFILLER_44_421 VPWR VGND sg13g2_decap_8
XFILLER_17_646 VPWR VGND sg13g2_decap_8
XFILLER_29_495 VPWR VGND sg13g2_decap_8
XFILLER_45_988 VPWR VGND sg13g2_decap_8
XFILLER_44_498 VPWR VGND sg13g2_decap_8
XFILLER_31_104 VPWR VGND sg13g2_fill_1
XFILLER_32_616 VPWR VGND sg13g2_decap_8
XFILLER_13_830 VPWR VGND sg13g2_decap_8
XFILLER_40_660 VPWR VGND sg13g2_decap_8
XFILLER_9_823 VPWR VGND sg13g2_decap_8
XFILLER_4_550 VPWR VGND sg13g2_decap_8
XFILLER_28_1009 VPWR VGND sg13g2_decap_8
X_3220_ _1699_ _1782_ _0691_ VPWR VGND sg13g2_nor2_1
X_3151_ VGND VPWR net717 _1991_ _0062_ _0625_ sg13g2_a21oi_1
X_2102_ VPWR _1520_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[0\]
+ VGND sg13g2_inv_1
X_3082_ sap_3_inst.alu_inst.tmp\[7\] _0363_ net772 _0579_ VPWR VGND sg13g2_nand3_1
XFILLER_36_911 VPWR VGND sg13g2_decap_8
XFILLER_36_988 VPWR VGND sg13g2_decap_8
XFILLER_23_627 VPWR VGND sg13g2_decap_8
XFILLER_35_498 VPWR VGND sg13g2_decap_8
X_3984_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[0\] _1353_
+ _1360_ net794 sg13g2_a21oi_1
X_2935_ net32 net693 _0436_ VPWR VGND sg13g2_nor2b_1
X_2866_ VGND VPWR _1525_ net703 _0370_ net694 sg13g2_a21oi_1
XFILLER_11_1013 VPWR VGND sg13g2_decap_8
X_2797_ _1794_ _0310_ _0311_ VPWR VGND sg13g2_nor2b_1
Xfanout802 sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[2\] net802 VPWR
+ VGND sg13g2_buf_8
Xfanout824 net825 net824 VPWR VGND sg13g2_buf_8
X_3418_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[1\] _0887_
+ net648 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[1\] _0888_ net671
+ sg13g2_a221oi_1
Xfanout813 net836 net813 VPWR VGND sg13g2_buf_8
X_3349_ _1522_ net690 _0749_ _0820_ VPWR VGND sg13g2_nor3_1
Xfanout835 net836 net835 VPWR VGND sg13g2_buf_8
XFILLER_39_760 VPWR VGND sg13g2_decap_8
XFILLER_26_432 VPWR VGND sg13g2_decap_8
XFILLER_27_966 VPWR VGND sg13g2_decap_8
XFILLER_42_947 VPWR VGND sg13g2_decap_8
XFILLER_13_126 VPWR VGND sg13g2_fill_1
XFILLER_42_33 VPWR VGND sg13g2_fill_1
XFILLER_10_800 VPWR VGND sg13g2_decap_8
XFILLER_10_877 VPWR VGND sg13g2_decap_8
XFILLER_6_848 VPWR VGND sg13g2_decap_8
XFILLER_1_520 VPWR VGND sg13g2_decap_8
XFILLER_49_524 VPWR VGND sg13g2_decap_8
XFILLER_1_597 VPWR VGND sg13g2_decap_8
XFILLER_18_900 VPWR VGND sg13g2_decap_8
XFILLER_37_719 VPWR VGND sg13g2_decap_8
XFILLER_18_977 VPWR VGND sg13g2_decap_8
XFILLER_45_785 VPWR VGND sg13g2_decap_8
XFILLER_33_925 VPWR VGND sg13g2_decap_8
XFILLER_9_620 VPWR VGND sg13g2_decap_8
X_2720_ VGND VPWR _0250_ _0249_ _1768_ sg13g2_or2_1
X_2651_ _2058_ sap_3_inst.alu_flags\[3\] _2057_ VPWR VGND sg13g2_nand2_1
XFILLER_9_697 VPWR VGND sg13g2_decap_8
X_2582_ sap_3_inst.alu_flags\[4\] net710 _1992_ VPWR VGND sg13g2_nor2_1
XFILLER_5_870 VPWR VGND sg13g2_decap_8
X_4321_ net824 VGND VPWR _0178_ sap_3_inst.alu_inst.act\[1\] clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4252_ net831 VGND VPWR _0109_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[3\]
+ clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3203_ _1673_ net720 net726 _0674_ VPWR VGND _0671_ sg13g2_nand4_1
XFILLER_41_1006 VPWR VGND sg13g2_decap_8
X_4183_ net820 VGND VPWR _0040_ sap_3_inst.alu_inst.acc\[7\] clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3134_ net32 sap_3_inst.alu_inst.tmp\[3\] net700 _0053_ VPWR VGND sg13g2_mux2_1
XFILLER_28_708 VPWR VGND sg13g2_decap_8
X_3065_ VGND VPWR sap_3_inst.alu_inst.act\[6\] net702 _0563_ net693 sg13g2_a21oi_1
XFILLER_36_785 VPWR VGND sg13g2_decap_8
XFILLER_23_424 VPWR VGND sg13g2_decap_8
XFILLER_24_969 VPWR VGND sg13g2_decap_8
X_3967_ net802 net801 _1342_ _1343_ VPWR VGND sg13g2_a21o_1
X_2918_ _0420_ _0393_ _0417_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_980 VPWR VGND sg13g2_decap_8
X_3898_ _1288_ VPWR _0146_ VGND _1520_ net649 sg13g2_o21ai_1
X_2849_ _2055_ _0337_ _0351_ _0352_ _0353_ VPWR VGND sg13g2_and4_1
XFILLER_5_8 VPWR VGND sg13g2_fill_2
Xfanout610 net611 net610 VPWR VGND sg13g2_buf_1
Xfanout621 _1856_ net621 VPWR VGND sg13g2_buf_8
Xfanout632 net633 net632 VPWR VGND sg13g2_buf_8
Xfanout643 net646 net643 VPWR VGND sg13g2_buf_8
Xfanout654 _0758_ net654 VPWR VGND sg13g2_buf_8
Xfanout665 _0712_ net665 VPWR VGND sg13g2_buf_8
Xfanout676 net679 net676 VPWR VGND sg13g2_buf_1
Xfanout698 _1438_ net698 VPWR VGND sg13g2_buf_8
Xfanout687 net688 net687 VPWR VGND sg13g2_buf_1
XFILLER_46_538 VPWR VGND sg13g2_decap_8
XFILLER_15_903 VPWR VGND sg13g2_decap_8
XFILLER_27_763 VPWR VGND sg13g2_decap_8
XFILLER_14_402 VPWR VGND sg13g2_fill_2
XFILLER_42_744 VPWR VGND sg13g2_decap_8
XFILLER_18_1019 VPWR VGND sg13g2_decap_8
XFILLER_26_295 VPWR VGND sg13g2_fill_1
XFILLER_30_917 VPWR VGND sg13g2_decap_8
XFILLER_23_991 VPWR VGND sg13g2_decap_8
XFILLER_6_645 VPWR VGND sg13g2_decap_8
XFILLER_10_674 VPWR VGND sg13g2_decap_8
XFILLER_2_862 VPWR VGND sg13g2_decap_8
XFILLER_49_321 VPWR VGND sg13g2_decap_8
XFILLER_37_516 VPWR VGND sg13g2_decap_8
XFILLER_49_398 VPWR VGND sg13g2_decap_8
XFILLER_45_582 VPWR VGND sg13g2_decap_8
XFILLER_18_774 VPWR VGND sg13g2_decap_8
XFILLER_33_722 VPWR VGND sg13g2_decap_8
X_3821_ _1060_ net635 _1235_ VPWR VGND sg13g2_nor2_1
XFILLER_33_799 VPWR VGND sg13g2_decap_8
X_3752_ net676 _0969_ _1187_ VPWR VGND sg13g2_nor2_1
X_3683_ _1132_ net609 _1021_ VPWR VGND sg13g2_nand2_1
XFILLER_9_494 VPWR VGND sg13g2_decap_8
X_2703_ _0234_ _0230_ _0233_ VPWR VGND sg13g2_xnor2_1
X_2634_ _2043_ net617 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[1\]
+ net619 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[1\] VPWR VGND
+ sg13g2_a22oi_1
X_2565_ _1976_ net618 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[4\]
+ net711 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4304_ net833 VGND VPWR _0161_ sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[0\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
X_2496_ net576 VPWR _1913_ VGND _1908_ _1912_ sg13g2_o21ai_1
X_4235_ net820 VGND VPWR _0092_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[2\]
+ clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4166_ net819 VGND VPWR _0027_ sap_3_inst.alu_flags\[3\] net38 sg13g2_dfrbpq_1
XFILLER_28_505 VPWR VGND sg13g2_decap_8
X_3117_ VPWR VGND net792 _0604_ net691 net772 _0605_ net692 sg13g2_a221oi_1
X_4097_ _1454_ sap_3_inst.alu_inst.act\[3\] net578 VPWR VGND sg13g2_nand2_1
X_3048_ _0542_ _0545_ _0546_ VPWR VGND sg13g2_nor2_1
XFILLER_36_582 VPWR VGND sg13g2_decap_8
XFILLER_24_766 VPWR VGND sg13g2_decap_8
XFILLER_20_994 VPWR VGND sg13g2_decap_8
XFILLER_3_637 VPWR VGND sg13g2_decap_8
XFILLER_2_169 VPWR VGND sg13g2_fill_2
XFILLER_47_858 VPWR VGND sg13g2_decap_8
XFILLER_46_335 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_15_700 VPWR VGND sg13g2_decap_8
XFILLER_27_560 VPWR VGND sg13g2_decap_8
XFILLER_42_541 VPWR VGND sg13g2_decap_8
XFILLER_15_777 VPWR VGND sg13g2_decap_8
XFILLER_30_714 VPWR VGND sg13g2_decap_8
XFILLER_11_950 VPWR VGND sg13g2_decap_8
XFILLER_6_420 VPWR VGND sg13g2_fill_2
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_7_954 VPWR VGND sg13g2_decap_8
Xsap_3_inst.clock.clock_gate_inst _0000_ clknet_1_0__leaf_clk_div_out sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_lgcp_1
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
X_2350_ _1567_ VPWR _1767_ VGND _1724_ _1766_ sg13g2_o21ai_1
X_2281_ VGND VPWR net726 _1682_ _1698_ net735 sg13g2_a21oi_1
X_4020_ _1393_ net49 net798 VPWR VGND sg13g2_nand2_1
XFILLER_38_825 VPWR VGND sg13g2_decap_8
XFILLER_18_571 VPWR VGND sg13g2_decap_8
XFILLER_33_596 VPWR VGND sg13g2_decap_8
XFILLER_21_769 VPWR VGND sg13g2_decap_8
X_3804_ _1225_ net681 _1154_ VPWR VGND sg13g2_nand2_1
XFILLER_20_279 VPWR VGND sg13g2_decap_4
X_3735_ _1173_ net655 _1062_ VPWR VGND sg13g2_nand2_1
X_3666_ net592 VPWR _1117_ VGND net638 _0969_ sg13g2_o21ai_1
XFILLER_47_1012 VPWR VGND sg13g2_decap_8
X_2617_ _2026_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[1\] net623
+ VPWR VGND sg13g2_nand2_1
X_3597_ _1059_ VPWR _0074_ VGND _1524_ _1054_ sg13g2_o21ai_1
X_2548_ _1961_ net625 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[5\]
+ net712 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[5\] VPWR VGND
+ sg13g2_a22oi_1
X_2479_ _1896_ net719 _1895_ VPWR VGND sg13g2_nand2_1
X_4218_ net808 VGND VPWR _0075_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[1\]
+ clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_29_803 VPWR VGND sg13g2_decap_8
XFILLER_44_806 VPWR VGND sg13g2_decap_8
XFILLER_37_880 VPWR VGND sg13g2_decap_8
XFILLER_24_563 VPWR VGND sg13g2_decap_8
XFILLER_11_224 VPWR VGND sg13g2_fill_2
XFILLER_12_758 VPWR VGND sg13g2_decap_8
Xclkload0 VPWR clkload0/Y clknet_3_1__leaf_clk VGND sg13g2_inv_1
XFILLER_20_791 VPWR VGND sg13g2_decap_8
XFILLER_4_935 VPWR VGND sg13g2_decap_8
XFILLER_47_655 VPWR VGND sg13g2_decap_8
XFILLER_35_806 VPWR VGND sg13g2_decap_8
XFILLER_43_850 VPWR VGND sg13g2_decap_8
XFILLER_15_574 VPWR VGND sg13g2_decap_8
XFILLER_30_511 VPWR VGND sg13g2_fill_1
XFILLER_30_588 VPWR VGND sg13g2_decap_8
XFILLER_7_751 VPWR VGND sg13g2_decap_8
X_3520_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[5\] _0985_
+ net649 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[5\] _0986_ net672
+ sg13g2_a221oi_1
X_3451_ VGND VPWR net661 _0919_ _0920_ _0918_ sg13g2_a21oi_1
X_2402_ _1784_ _1817_ _1708_ _1819_ VPWR VGND _1818_ sg13g2_nand4_1
X_3382_ _0770_ _0780_ _0852_ _0853_ VPWR VGND sg13g2_nor3_1
X_2333_ _1596_ _1749_ _1750_ VPWR VGND sg13g2_nor2_1
X_2264_ _1681_ net745 _1580_ VPWR VGND sg13g2_nand2_1
XFILLER_38_622 VPWR VGND sg13g2_decap_8
X_2195_ net738 net736 _1612_ VPWR VGND sg13g2_and2_1
X_4003_ _1377_ _1375_ _1376_ VPWR VGND sg13g2_nand2_1
XFILLER_26_817 VPWR VGND sg13g2_decap_8
XFILLER_38_699 VPWR VGND sg13g2_decap_8
XFILLER_34_850 VPWR VGND sg13g2_decap_8
XFILLER_40_319 VPWR VGND sg13g2_fill_2
XFILLER_21_566 VPWR VGND sg13g2_decap_8
X_3718_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[4\] _1160_ _1147_
+ _0094_ VPWR VGND sg13g2_mux2_1
X_3649_ _1103_ net594 _0894_ VPWR VGND sg13g2_nand2_1
XFILLER_1_905 VPWR VGND sg13g2_decap_8
XFILLER_49_909 VPWR VGND sg13g2_decap_8
Xhold12 u_ser.shadow_reg\[3\] VPWR VGND net59 sg13g2_dlygate4sd3_1
XFILLER_0_448 VPWR VGND sg13g2_decap_8
Xhold23 regFile_serial VPWR VGND net70 sg13g2_dlygate4sd3_1
XFILLER_29_600 VPWR VGND sg13g2_decap_8
XFILLER_44_603 VPWR VGND sg13g2_decap_8
XFILLER_17_828 VPWR VGND sg13g2_decap_8
XFILLER_29_677 VPWR VGND sg13g2_decap_8
XFILLER_28_187 VPWR VGND sg13g2_fill_2
XFILLER_40_842 VPWR VGND sg13g2_decap_8
XFILLER_12_555 VPWR VGND sg13g2_decap_8
XFILLER_6_38 VPWR VGND sg13g2_fill_2
XFILLER_4_732 VPWR VGND sg13g2_decap_8
XFILLER_3_231 VPWR VGND sg13g2_fill_2
XFILLER_6_1009 VPWR VGND sg13g2_decap_8
XFILLER_48_920 VPWR VGND sg13g2_decap_8
XFILLER_48_997 VPWR VGND sg13g2_decap_8
XFILLER_47_452 VPWR VGND sg13g2_decap_8
XFILLER_35_603 VPWR VGND sg13g2_decap_8
XFILLER_23_809 VPWR VGND sg13g2_decap_8
X_2951_ _0346_ VPWR _0452_ VGND _0349_ _0413_ sg13g2_o21ai_1
XFILLER_31_831 VPWR VGND sg13g2_decap_8
X_2882_ _0385_ net789 net709 VPWR VGND sg13g2_nand2_1
X_3503_ net592 VPWR _0970_ VGND net663 _0969_ sg13g2_o21ai_1
X_3434_ VGND VPWR _2051_ net605 _0904_ _0903_ sg13g2_a21oi_1
X_3365_ _0830_ _0835_ _0836_ VPWR VGND sg13g2_and2_1
X_2316_ _1733_ _1587_ net732 VPWR VGND sg13g2_nand2_1
X_3296_ _0767_ net639 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[0\]
+ net642 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_942 VPWR VGND sg13g2_decap_8
X_2247_ _1648_ _1654_ _1657_ _1663_ _1664_ VPWR VGND sg13g2_nor4_1
XFILLER_26_614 VPWR VGND sg13g2_decap_8
X_2178_ net755 net753 _1595_ VPWR VGND sg13g2_nor2b_2
XFILLER_38_496 VPWR VGND sg13g2_decap_8
XFILLER_41_628 VPWR VGND sg13g2_decap_8
XFILLER_22_886 VPWR VGND sg13g2_decap_8
XFILLER_1_702 VPWR VGND sg13g2_decap_8
Xoutput24 net24 uio_out[7] VPWR VGND sg13g2_buf_1
Xoutput13 net13 uio_oe[4] VPWR VGND sg13g2_buf_1
XFILLER_49_706 VPWR VGND sg13g2_decap_8
XFILLER_1_779 VPWR VGND sg13g2_decap_8
XFILLER_16_102 VPWR VGND sg13g2_fill_1
XFILLER_17_625 VPWR VGND sg13g2_decap_8
XFILLER_29_474 VPWR VGND sg13g2_decap_8
XFILLER_45_967 VPWR VGND sg13g2_decap_8
XFILLER_44_477 VPWR VGND sg13g2_decap_8
XFILLER_9_802 VPWR VGND sg13g2_decap_8
XFILLER_12_341 VPWR VGND sg13g2_fill_1
XFILLER_13_886 VPWR VGND sg13g2_decap_8
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_9_879 VPWR VGND sg13g2_decap_8
X_3150_ net759 net717 _0625_ VPWR VGND sg13g2_nor2_1
X_3081_ _0578_ _0572_ _0577_ VPWR VGND sg13g2_xnor2_1
X_2101_ VPWR _1519_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[1\]
+ VGND sg13g2_inv_1
XFILLER_48_794 VPWR VGND sg13g2_decap_8
XFILLER_23_606 VPWR VGND sg13g2_decap_8
XFILLER_36_967 VPWR VGND sg13g2_decap_8
X_3983_ _1356_ _1357_ _1354_ _1359_ VPWR VGND _1358_ sg13g2_nand4_1
X_2934_ net598 net787 _0435_ _0035_ VPWR VGND sg13g2_a21o_1
X_2865_ _0368_ VPWR _0369_ VGND net792 _0337_ sg13g2_o21ai_1
XFILLER_30_160 VPWR VGND sg13g2_fill_1
X_2796_ net724 VPWR _0310_ VGND _1650_ _1685_ sg13g2_o21ai_1
Xfanout814 net816 net814 VPWR VGND sg13g2_buf_8
Xfanout825 net826 net825 VPWR VGND sg13g2_buf_8
X_3417_ _0885_ _0886_ net660 _0887_ VPWR VGND sg13g2_nand3_1
Xfanout803 net79 net803 VPWR VGND sg13g2_buf_8
Xfanout836 rst_n net836 VPWR VGND sg13g2_buf_8
X_3348_ _0819_ _0817_ _0818_ VPWR VGND sg13g2_nand2_1
X_3279_ _0653_ _0665_ _0708_ _0750_ VPWR VGND sg13g2_nor3_1
XFILLER_27_945 VPWR VGND sg13g2_decap_8
XFILLER_42_926 VPWR VGND sg13g2_decap_8
XFILLER_14_639 VPWR VGND sg13g2_decap_8
XFILLER_26_488 VPWR VGND sg13g2_decap_8
XFILLER_22_683 VPWR VGND sg13g2_decap_8
XFILLER_6_827 VPWR VGND sg13g2_decap_8
XFILLER_10_856 VPWR VGND sg13g2_decap_8
XFILLER_49_503 VPWR VGND sg13g2_decap_8
XFILLER_1_576 VPWR VGND sg13g2_decap_8
XFILLER_29_282 VPWR VGND sg13g2_decap_4
XFILLER_45_764 VPWR VGND sg13g2_decap_8
XFILLER_18_956 VPWR VGND sg13g2_decap_8
XFILLER_33_904 VPWR VGND sg13g2_decap_8
XFILLER_17_499 VPWR VGND sg13g2_decap_8
XFILLER_20_609 VPWR VGND sg13g2_decap_8
XFILLER_41_992 VPWR VGND sg13g2_decap_8
XFILLER_13_683 VPWR VGND sg13g2_decap_8
XFILLER_34_1025 VPWR VGND sg13g2_decap_4
XFILLER_9_676 VPWR VGND sg13g2_decap_8
XFILLER_12_193 VPWR VGND sg13g2_fill_2
X_2650_ _2057_ _2003_ _2056_ VPWR VGND sg13g2_nand2_2
X_2581_ net21 _1991_ VPWR VGND sg13g2_inv_4
X_4320_ net824 VGND VPWR _0177_ sap_3_inst.alu_inst.act\[0\] clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4251_ net827 VGND VPWR _0108_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[2\]
+ clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3202_ VGND VPWR _0673_ _0671_ net735 sg13g2_or2_1
X_4182_ net825 VGND VPWR _0039_ sap_3_inst.alu_inst.acc\[6\] clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3133_ _0617_ VPWR _0052_ VGND _0227_ net700 sg13g2_o21ai_1
X_3064_ VPWR VGND _0539_ net702 _0561_ _0353_ _0562_ _0556_ sg13g2_a221oi_1
XFILLER_48_591 VPWR VGND sg13g2_decap_8
XFILLER_36_764 VPWR VGND sg13g2_decap_8
XFILLER_35_263 VPWR VGND sg13g2_fill_1
XFILLER_24_948 VPWR VGND sg13g2_decap_8
X_3966_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[0\] sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[1\]
+ net801 net802 _1342_ VPWR VGND sg13g2_nor4_1
X_2917_ VPWR _0419_ _0418_ VGND sg13g2_inv_1
X_3897_ _0870_ _1287_ net649 _1288_ VPWR VGND sg13g2_nand3_1
X_2848_ _0352_ _2005_ _2008_ VPWR VGND sg13g2_nand2_1
XFILLER_3_819 VPWR VGND sg13g2_decap_8
X_2779_ VPWR net9 _0301_ VGND sg13g2_inv_1
Xfanout633 _1845_ net633 VPWR VGND sg13g2_buf_8
Xfanout611 _0857_ net611 VPWR VGND sg13g2_buf_8
Xfanout622 net623 net622 VPWR VGND sg13g2_buf_8
Xfanout600 _1862_ net600 VPWR VGND sg13g2_buf_8
Xfanout644 net646 net644 VPWR VGND sg13g2_buf_1
Xfanout655 _0754_ net655 VPWR VGND sg13g2_buf_8
Xfanout666 _1828_ net666 VPWR VGND sg13g2_buf_2
Xfanout699 _1438_ net699 VPWR VGND sg13g2_buf_2
Xfanout688 _0711_ net688 VPWR VGND sg13g2_buf_8
Xfanout677 net679 net677 VPWR VGND sg13g2_buf_8
XFILLER_46_517 VPWR VGND sg13g2_decap_8
XFILLER_2_1023 VPWR VGND sg13g2_decap_4
XFILLER_27_742 VPWR VGND sg13g2_decap_8
XFILLER_42_723 VPWR VGND sg13g2_decap_8
XFILLER_14_447 VPWR VGND sg13g2_fill_1
XFILLER_15_959 VPWR VGND sg13g2_decap_8
XFILLER_23_970 VPWR VGND sg13g2_decap_8
XFILLER_22_480 VPWR VGND sg13g2_decap_8
XFILLER_10_653 VPWR VGND sg13g2_decap_8
XFILLER_6_624 VPWR VGND sg13g2_decap_8
XFILLER_2_841 VPWR VGND sg13g2_decap_8
XFILLER_49_300 VPWR VGND sg13g2_decap_8
XFILLER_49_377 VPWR VGND sg13g2_decap_8
XFILLER_18_753 VPWR VGND sg13g2_decap_8
XFILLER_45_561 VPWR VGND sg13g2_decap_8
XFILLER_33_701 VPWR VGND sg13g2_decap_8
XFILLER_17_285 VPWR VGND sg13g2_fill_1
X_3820_ net635 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[0\] _1234_
+ _0122_ VPWR VGND sg13g2_a21o_1
XFILLER_33_778 VPWR VGND sg13g2_decap_8
X_3751_ _1181_ _1186_ _0101_ VPWR VGND sg13g2_nor2b_1
XFILLER_9_462 VPWR VGND sg13g2_fill_1
XFILLER_13_480 VPWR VGND sg13g2_decap_8
X_2702_ _0233_ _0231_ _0232_ VPWR VGND sg13g2_xnor2_1
X_3682_ _1131_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[6\] net637
+ VPWR VGND sg13g2_nand2_1
X_2633_ net667 net627 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[1\]
+ _2042_ VPWR VGND sg13g2_nand3_1
X_2564_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[4\] net614
+ _1975_ net631 sg13g2_a21oi_1
X_4303_ net833 VGND VPWR _0160_ regFile_serial clknet_3_6__leaf_clk sg13g2_dfrbpq_1
X_2495_ _1910_ _1911_ _1909_ _1912_ VPWR VGND sg13g2_nand3_1
X_4234_ net808 VGND VPWR _0091_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[1\]
+ clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4165_ net819 VGND VPWR _0026_ sap_3_inst.alu_flags\[2\] net37 sg13g2_dfrbpq_1
X_3116_ VGND VPWR sap_3_inst.alu_flags\[1\] _2017_ _0604_ _0603_ sg13g2_a21oi_1
X_4096_ _1452_ VPWR _1453_ VGND net784 net699 sg13g2_o21ai_1
X_3047_ VGND VPWR net778 _1527_ _0545_ _0514_ sg13g2_a21oi_1
XFILLER_36_561 VPWR VGND sg13g2_decap_8
XFILLER_24_745 VPWR VGND sg13g2_decap_8
XFILLER_11_439 VPWR VGND sg13g2_fill_2
XFILLER_23_288 VPWR VGND sg13g2_decap_4
XFILLER_23_58 VPWR VGND sg13g2_fill_2
X_3949_ _1325_ VPWR _1326_ VGND net803 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[1\]
+ sg13g2_o21ai_1
XFILLER_20_973 VPWR VGND sg13g2_decap_8
XFILLER_3_616 VPWR VGND sg13g2_decap_8
XFILLER_2_115 VPWR VGND sg13g2_fill_2
XFILLER_48_22 VPWR VGND sg13g2_fill_2
XFILLER_47_837 VPWR VGND sg13g2_decap_8
XFILLER_19_539 VPWR VGND sg13g2_decap_8
XFILLER_0_18 VPWR VGND sg13g2_fill_1
XFILLER_42_520 VPWR VGND sg13g2_decap_8
XFILLER_15_756 VPWR VGND sg13g2_decap_8
XFILLER_42_597 VPWR VGND sg13g2_decap_8
Xclkbuf_5_5__f_sap_3_inst.alu_inst.clk_regs clknet_4_2_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_31_1006 VPWR VGND sg13g2_decap_8
XFILLER_7_933 VPWR VGND sg13g2_decap_8
XFILLER_6_498 VPWR VGND sg13g2_decap_8
X_2280_ net726 _1607_ _1697_ VPWR VGND sg13g2_nor2_2
XFILLER_38_804 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_2_sap_3_inst.alu_inst.clk clknet_1_0__leaf_sap_3_inst.alu_inst.clk clknet_leaf_2_sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_18_550 VPWR VGND sg13g2_decap_8
XFILLER_46_881 VPWR VGND sg13g2_decap_8
X_3803_ _1224_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[2\] net658
+ VPWR VGND sg13g2_nand2_1
XFILLER_33_575 VPWR VGND sg13g2_decap_8
XFILLER_21_748 VPWR VGND sg13g2_decap_8
X_3734_ _1171_ VPWR _1172_ VGND net18 net602 sg13g2_o21ai_1
X_3665_ VPWR _0085_ _1116_ VGND sg13g2_inv_1
X_2616_ _2025_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[1\] net629
+ VPWR VGND sg13g2_nand2_1
X_3596_ net583 _1057_ _1058_ _1059_ VPWR VGND sg13g2_or3_1
X_2547_ _1960_ _1862_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[5\]
+ net617 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[5\] VPWR VGND sg13g2_a22oi_1
X_2478_ _1895_ _1592_ _1629_ VPWR VGND sg13g2_nand2_1
X_4217_ net828 VGND VPWR _0074_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[0\]
+ clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_29_859 VPWR VGND sg13g2_decap_8
X_4079_ _1439_ net698 VPWR VGND sg13g2_inv_2
XFILLER_24_542 VPWR VGND sg13g2_decap_8
XFILLER_12_737 VPWR VGND sg13g2_decap_8
Xclkload1 clknet_3_2__leaf_clk clkload1/X VPWR VGND sg13g2_buf_1
XFILLER_20_770 VPWR VGND sg13g2_decap_8
XFILLER_4_914 VPWR VGND sg13g2_decap_8
XFILLER_47_634 VPWR VGND sg13g2_decap_8
XFILLER_34_339 VPWR VGND sg13g2_fill_1
XFILLER_15_553 VPWR VGND sg13g2_decap_8
XFILLER_30_567 VPWR VGND sg13g2_decap_8
XFILLER_7_730 VPWR VGND sg13g2_decap_8
X_3450_ _0919_ _0836_ _0848_ VPWR VGND sg13g2_xnor2_1
X_2401_ _1818_ _1692_ _1777_ _1688_ _1654_ VPWR VGND sg13g2_a22oi_1
X_3381_ _0793_ _0802_ _0786_ _0852_ VPWR VGND _0850_ sg13g2_nand4_1
X_2332_ _1749_ net731 _1617_ VPWR VGND sg13g2_nand2_1
XFILLER_3_980 VPWR VGND sg13g2_decap_8
X_2263_ _1680_ sap_3_inst.controller_inst.stage\[2\] net744 VPWR VGND sg13g2_nand2_1
X_4002_ _1376_ _1352_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[2\]
+ _1340_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_38_601 VPWR VGND sg13g2_decap_8
X_2194_ _1611_ net745 VPWR VGND net744 sg13g2_nand2b_2
XFILLER_37_111 VPWR VGND sg13g2_fill_2
XFILLER_38_678 VPWR VGND sg13g2_decap_8
XFILLER_37_188 VPWR VGND sg13g2_fill_2
XFILLER_33_361 VPWR VGND sg13g2_fill_1
XFILLER_21_545 VPWR VGND sg13g2_decap_8
X_3717_ _1075_ _0974_ _1160_ VPWR VGND _1074_ sg13g2_nand3b_1
X_3648_ _1102_ VPWR _0082_ VGND _1523_ net639 sg13g2_o21ai_1
X_3579_ _1043_ _0779_ _0852_ VPWR VGND sg13g2_xnor2_1
XFILLER_48_409 VPWR VGND sg13g2_decap_8
Xhold13 u_ser.shadow_reg\[1\] VPWR VGND net60 sg13g2_dlygate4sd3_1
Xhold24 u_ser.bit_pos\[1\] VPWR VGND net71 sg13g2_dlygate4sd3_1
XFILLER_29_656 VPWR VGND sg13g2_decap_8
XFILLER_17_807 VPWR VGND sg13g2_decap_8
XFILLER_44_659 VPWR VGND sg13g2_decap_8
XFILLER_40_821 VPWR VGND sg13g2_decap_8
XFILLER_24_372 VPWR VGND sg13g2_fill_1
XFILLER_25_884 VPWR VGND sg13g2_decap_8
XFILLER_12_534 VPWR VGND sg13g2_decap_8
XFILLER_40_898 VPWR VGND sg13g2_decap_8
XFILLER_8_549 VPWR VGND sg13g2_decap_8
XFILLER_4_711 VPWR VGND sg13g2_decap_8
XFILLER_4_788 VPWR VGND sg13g2_decap_8
XFILLER_47_431 VPWR VGND sg13g2_decap_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
XFILLER_48_976 VPWR VGND sg13g2_decap_8
XFILLER_35_659 VPWR VGND sg13g2_decap_8
X_2950_ _0445_ _0447_ _0450_ _0451_ VPWR VGND sg13g2_nor3_1
XFILLER_16_884 VPWR VGND sg13g2_decap_8
XFILLER_31_810 VPWR VGND sg13g2_decap_8
X_2881_ _0384_ net792 net692 VPWR VGND sg13g2_nand2_1
XFILLER_31_887 VPWR VGND sg13g2_decap_8
X_3502_ _0969_ _0802_ _0850_ VPWR VGND sg13g2_xnor2_1
X_3433_ net10 net605 _0903_ VPWR VGND sg13g2_nor2_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_44_1016 VPWR VGND sg13g2_decap_8
X_3364_ _0831_ _0832_ _0833_ _0834_ _0835_ VPWR VGND sg13g2_nor4_1
XFILLER_32_0 VPWR VGND sg13g2_fill_2
XFILLER_39_921 VPWR VGND sg13g2_decap_8
X_2315_ VPWR _1732_ _1731_ VGND sg13g2_inv_1
X_3295_ _0766_ _0748_ VPWR VGND net689 sg13g2_nand2b_2
X_2246_ _1663_ _1607_ net733 VPWR VGND sg13g2_nand2_1
XFILLER_39_998 VPWR VGND sg13g2_decap_8
X_2177_ net739 _1593_ _1594_ VPWR VGND sg13g2_nor2_1
XFILLER_38_475 VPWR VGND sg13g2_decap_8
XFILLER_41_607 VPWR VGND sg13g2_decap_8
XFILLER_15_59 VPWR VGND sg13g2_fill_1
XFILLER_21_331 VPWR VGND sg13g2_fill_1
XFILLER_22_865 VPWR VGND sg13g2_decap_8
Xoutput25 net25 uo_out[0] VPWR VGND sg13g2_buf_1
Xoutput14 net14 uio_oe[5] VPWR VGND sg13g2_buf_1
XFILLER_1_758 VPWR VGND sg13g2_decap_8
XFILLER_5_1010 VPWR VGND sg13g2_decap_8
XFILLER_17_604 VPWR VGND sg13g2_decap_8
XFILLER_45_946 VPWR VGND sg13g2_decap_8
XFILLER_44_456 VPWR VGND sg13g2_decap_8
XFILLER_25_681 VPWR VGND sg13g2_decap_8
XFILLER_13_865 VPWR VGND sg13g2_decap_8
XFILLER_40_695 VPWR VGND sg13g2_decap_8
XFILLER_9_858 VPWR VGND sg13g2_decap_8
XFILLER_4_585 VPWR VGND sg13g2_decap_8
X_3080_ VGND VPWR net775 _1528_ _0577_ _0546_ sg13g2_a21oi_1
XFILLER_0_791 VPWR VGND sg13g2_decap_8
X_2100_ VPWR _1518_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[1\]
+ VGND sg13g2_inv_1
XFILLER_48_773 VPWR VGND sg13g2_decap_8
XFILLER_36_946 VPWR VGND sg13g2_decap_8
XFILLER_35_434 VPWR VGND sg13g2_fill_1
X_3982_ _1358_ _1351_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[0\]
+ net796 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_16_681 VPWR VGND sg13g2_decap_8
X_2933_ VPWR VGND _0434_ net598 _0433_ _0227_ _0435_ net693 sg13g2_a221oi_1
X_2864_ VPWR VGND _0367_ _0365_ _0366_ _0342_ _0368_ _0356_ sg13g2_a221oi_1
XFILLER_31_684 VPWR VGND sg13g2_decap_8
X_2795_ VGND VPWR net726 _0308_ _0309_ _1725_ sg13g2_a21oi_1
Xfanout815 net816 net815 VPWR VGND sg13g2_buf_8
Xfanout804 net806 net804 VPWR VGND sg13g2_buf_8
X_3416_ _0886_ net675 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[1\]
+ net680 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[1\] VPWR VGND sg13g2_a22oi_1
Xfanout826 net836 net826 VPWR VGND sg13g2_buf_8
X_3347_ _0818_ net677 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[0\]
+ net684 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[0\] VPWR VGND sg13g2_a22oi_1
X_3278_ _0749_ _0652_ _0664_ VPWR VGND sg13g2_nand2_2
X_2229_ _1646_ _1574_ _1623_ VPWR VGND sg13g2_nand2_2
XFILLER_27_924 VPWR VGND sg13g2_decap_8
XFILLER_39_795 VPWR VGND sg13g2_decap_8
XFILLER_42_905 VPWR VGND sg13g2_decap_8
XFILLER_14_618 VPWR VGND sg13g2_decap_8
XFILLER_26_467 VPWR VGND sg13g2_decap_8
XFILLER_13_139 VPWR VGND sg13g2_fill_2
XFILLER_22_662 VPWR VGND sg13g2_decap_8
XFILLER_10_835 VPWR VGND sg13g2_decap_8
XFILLER_6_806 VPWR VGND sg13g2_decap_8
XFILLER_1_555 VPWR VGND sg13g2_decap_8
XFILLER_27_1022 VPWR VGND sg13g2_decap_8
XFILLER_49_559 VPWR VGND sg13g2_decap_8
XFILLER_18_935 VPWR VGND sg13g2_decap_8
XFILLER_45_743 VPWR VGND sg13g2_decap_8
XFILLER_17_478 VPWR VGND sg13g2_decap_8
XFILLER_41_971 VPWR VGND sg13g2_decap_8
XFILLER_13_662 VPWR VGND sg13g2_decap_8
XFILLER_34_1004 VPWR VGND sg13g2_decap_8
XFILLER_12_161 VPWR VGND sg13g2_fill_2
XFILLER_40_492 VPWR VGND sg13g2_decap_8
XFILLER_9_655 VPWR VGND sg13g2_decap_8
X_2580_ _1982_ _1990_ _1979_ net21 VPWR VGND sg13g2_nand3_1
X_4250_ net833 VGND VPWR _0107_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[1\]
+ clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3201_ _0672_ _1673_ net720 VPWR VGND sg13g2_nand2_1
X_4181_ net823 VGND VPWR _0038_ sap_3_inst.alu_inst.acc\[5\] clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3132_ _0617_ sap_3_inst.alu_inst.tmp\[2\] net700 VPWR VGND sg13g2_nand2_1
XFILLER_48_570 VPWR VGND sg13g2_decap_8
X_3063_ _0353_ _0551_ _0560_ _0561_ VPWR VGND sg13g2_nor3_1
XFILLER_35_220 VPWR VGND sg13g2_fill_2
XFILLER_36_743 VPWR VGND sg13g2_decap_8
XFILLER_24_927 VPWR VGND sg13g2_decap_8
X_3965_ _1341_ net801 VPWR VGND net802 sg13g2_nand2b_2
XFILLER_23_459 VPWR VGND sg13g2_decap_8
X_2916_ _0393_ _0417_ _0418_ VPWR VGND sg13g2_nor2b_1
X_3896_ _1095_ VPWR _1287_ VGND _0301_ _1285_ sg13g2_o21ai_1
X_2847_ _0344_ _0350_ _0351_ VPWR VGND sg13g2_nor2_1
X_2778_ _0301_ net577 VPWR VGND _0249_ sg13g2_nand2b_2
Xfanout612 _0745_ net612 VPWR VGND sg13g2_buf_8
Xfanout601 _1850_ net601 VPWR VGND sg13g2_buf_8
Xfanout623 _1853_ net623 VPWR VGND sg13g2_buf_8
Xfanout645 net646 net645 VPWR VGND sg13g2_buf_8
Xfanout634 _1233_ net634 VPWR VGND sg13g2_buf_8
Xfanout656 _0754_ net656 VPWR VGND sg13g2_buf_2
Xfanout667 _1809_ net667 VPWR VGND sg13g2_buf_8
Xfanout689 _0709_ net689 VPWR VGND sg13g2_buf_8
Xfanout678 net679 net678 VPWR VGND sg13g2_buf_8
XFILLER_2_1002 VPWR VGND sg13g2_decap_8
XFILLER_27_721 VPWR VGND sg13g2_decap_8
XFILLER_26_220 VPWR VGND sg13g2_fill_1
XFILLER_39_592 VPWR VGND sg13g2_decap_8
XFILLER_42_702 VPWR VGND sg13g2_decap_8
XFILLER_15_938 VPWR VGND sg13g2_decap_8
XFILLER_27_798 VPWR VGND sg13g2_decap_8
XFILLER_42_779 VPWR VGND sg13g2_decap_8
XFILLER_6_603 VPWR VGND sg13g2_decap_8
XFILLER_10_632 VPWR VGND sg13g2_decap_8
XFILLER_5_124 VPWR VGND sg13g2_fill_1
XFILLER_2_820 VPWR VGND sg13g2_decap_8
XFILLER_1_330 VPWR VGND sg13g2_fill_2
XFILLER_2_897 VPWR VGND sg13g2_decap_8
XFILLER_49_356 VPWR VGND sg13g2_decap_8
XFILLER_18_732 VPWR VGND sg13g2_decap_8
XFILLER_45_540 VPWR VGND sg13g2_decap_8
XFILLER_33_757 VPWR VGND sg13g2_decap_8
XFILLER_14_982 VPWR VGND sg13g2_decap_8
X_3750_ _1182_ _1183_ net678 _1186_ VPWR VGND _1185_ sg13g2_nand4_1
X_2701_ net788 net785 _0232_ VPWR VGND sg13g2_xor2_1
X_3681_ _0087_ _1125_ _1130_ net637 _1538_ VPWR VGND sg13g2_a22oi_1
X_2632_ _2041_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[1\] net630
+ VPWR VGND sg13g2_nand2_1
X_2563_ _1974_ net600 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[4\]
+ net624 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4302_ net833 VGND VPWR net74 regFile_serial_start clknet_3_4__leaf_clk sg13g2_dfrbpq_1
X_4233_ net828 VGND VPWR _0090_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[0\]
+ clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_2494_ _1911_ net622 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[7\]
+ net601 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4164_ net819 VGND VPWR _0025_ sap_3_inst.alu_flags\[0\] net36 sg13g2_dfrbpq_1
X_3115_ _2004_ _2006_ net761 _0603_ VPWR VGND sg13g2_nand3_1
X_4095_ _1452_ net699 _0444_ VPWR VGND sg13g2_nand2b_1
X_3046_ _0361_ VPWR _0544_ VGND net776 sap_3_inst.alu_inst.tmp\[6\] sg13g2_o21ai_1
XFILLER_36_540 VPWR VGND sg13g2_decap_8
XFILLER_24_724 VPWR VGND sg13g2_decap_8
XFILLER_12_919 VPWR VGND sg13g2_decap_8
XFILLER_17_1010 VPWR VGND sg13g2_decap_8
XFILLER_20_952 VPWR VGND sg13g2_decap_8
X_3948_ VGND VPWR net803 _1549_ _1325_ sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[1\]
+ sg13g2_a21oi_1
X_3879_ net654 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[0\] _1277_
+ _0138_ VPWR VGND sg13g2_a21o_1
XFILLER_2_149 VPWR VGND sg13g2_fill_2
XFILLER_24_1025 VPWR VGND sg13g2_decap_4
XFILLER_47_816 VPWR VGND sg13g2_decap_8
XFILLER_19_518 VPWR VGND sg13g2_decap_8
XFILLER_15_735 VPWR VGND sg13g2_decap_8
XFILLER_27_595 VPWR VGND sg13g2_decap_8
XFILLER_42_576 VPWR VGND sg13g2_decap_8
XFILLER_30_749 VPWR VGND sg13g2_decap_8
XFILLER_7_912 VPWR VGND sg13g2_decap_8
XFILLER_11_985 VPWR VGND sg13g2_decap_8
XFILLER_7_989 VPWR VGND sg13g2_decap_8
XFILLER_6_477 VPWR VGND sg13g2_decap_8
XFILLER_9_1019 VPWR VGND sg13g2_decap_8
XFILLER_2_694 VPWR VGND sg13g2_decap_8
XFILLER_46_860 VPWR VGND sg13g2_decap_8
XFILLER_33_554 VPWR VGND sg13g2_decap_8
XFILLER_21_727 VPWR VGND sg13g2_decap_8
X_3802_ _0115_ _1063_ _1223_ net657 _1515_ VPWR VGND sg13g2_a22oi_1
X_3733_ _1171_ _0302_ net602 VPWR VGND sg13g2_nand2_1
X_3664_ _1116_ _1114_ _1115_ net637 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[3\]
+ VPWR VGND sg13g2_a22oi_1
X_2615_ VGND VPWR _1916_ _2002_ _2024_ _2023_ sg13g2_a21oi_1
X_3595_ net591 net588 _1058_ VPWR VGND sg13g2_nor2_2
X_2546_ _1959_ net614 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[5\]
+ net618 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[5\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_0_609 VPWR VGND sg13g2_decap_8
X_2477_ net729 _1617_ _1894_ VPWR VGND sg13g2_nor2_1
Xclkbuf_5_29__f_sap_3_inst.alu_inst.clk_regs clknet_4_14_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
X_4216_ net809 VGND VPWR _0073_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[7\]
+ clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_1
XFILLER_29_838 VPWR VGND sg13g2_decap_8
X_4078_ _1438_ _0321_ _0322_ net723 _1592_ VPWR VGND sg13g2_a22oi_1
X_3029_ VPWR VGND _0348_ _0527_ _0524_ _0344_ _0528_ _0521_ sg13g2_a221oi_1
XFILLER_24_521 VPWR VGND sg13g2_decap_8
XFILLER_12_716 VPWR VGND sg13g2_decap_8
XFILLER_24_598 VPWR VGND sg13g2_decap_8
Xclkload2 VPWR clkload2/Y clknet_3_3__leaf_clk VGND sg13g2_inv_1
XFILLER_3_469 VPWR VGND sg13g2_decap_8
XFILLER_1_4 VPWR VGND sg13g2_decap_4
Xclkbuf_5_18__f_sap_3_inst.alu_inst.clk_regs clknet_4_9_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_47_613 VPWR VGND sg13g2_decap_8
XFILLER_46_189 VPWR VGND sg13g2_fill_2
XFILLER_15_532 VPWR VGND sg13g2_decap_8
XFILLER_43_885 VPWR VGND sg13g2_decap_8
XFILLER_30_546 VPWR VGND sg13g2_decap_8
XFILLER_11_782 VPWR VGND sg13g2_decap_8
XFILLER_7_786 VPWR VGND sg13g2_decap_8
X_2400_ net759 VPWR _1817_ VGND _1800_ _1815_ sg13g2_o21ai_1
X_3380_ _0802_ _0850_ _0793_ _0851_ VPWR VGND sg13g2_nand3_1
X_2331_ _1609_ _1630_ _1748_ VPWR VGND sg13g2_nor2_1
XFILLER_2_491 VPWR VGND sg13g2_decap_8
X_2262_ net745 net744 _1679_ VPWR VGND sg13g2_and2_1
X_4001_ _1375_ _1353_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[2\]
+ _1347_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2193_ net744 net745 _1610_ VPWR VGND sg13g2_nor2b_2
XFILLER_1_73 VPWR VGND sg13g2_fill_2
XFILLER_38_657 VPWR VGND sg13g2_decap_8
XFILLER_19_882 VPWR VGND sg13g2_decap_8
XFILLER_25_318 VPWR VGND sg13g2_decap_4
XFILLER_25_329 VPWR VGND sg13g2_fill_2
Xclkbuf_0_sap_3_inst.alu_inst.clk sap_3_inst.alu_inst.clk clknet_0_sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_34_885 VPWR VGND sg13g2_decap_8
XFILLER_21_524 VPWR VGND sg13g2_decap_8
XFILLER_14_1024 VPWR VGND sg13g2_decap_4
X_3716_ VGND VPWR _1147_ _1159_ _0093_ _1158_ sg13g2_a21oi_1
XFILLER_20_38 VPWR VGND sg13g2_fill_1
X_3647_ _0870_ _1101_ net639 _1102_ VPWR VGND sg13g2_nand3_1
X_3578_ _1042_ net664 _1041_ VPWR VGND sg13g2_nand2_1
X_2529_ VGND VPWR net710 net570 _0031_ _1942_ sg13g2_a21oi_1
Xhold14 sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[2\] VPWR VGND net61
+ sg13g2_dlygate4sd3_1
Xhold25 u_ser.shadow_reg\[6\] VPWR VGND net72 sg13g2_dlygate4sd3_1
XFILLER_29_635 VPWR VGND sg13g2_decap_8
XFILLER_21_1028 VPWR VGND sg13g2_fill_1
XFILLER_44_638 VPWR VGND sg13g2_decap_8
XFILLER_28_189 VPWR VGND sg13g2_fill_1
XFILLER_40_800 VPWR VGND sg13g2_decap_8
XFILLER_25_863 VPWR VGND sg13g2_decap_8
XFILLER_12_513 VPWR VGND sg13g2_decap_8
XFILLER_40_877 VPWR VGND sg13g2_decap_8
XFILLER_8_528 VPWR VGND sg13g2_decap_8
XFILLER_4_767 VPWR VGND sg13g2_decap_8
XFILLER_0_973 VPWR VGND sg13g2_decap_8
XFILLER_48_955 VPWR VGND sg13g2_decap_8
XFILLER_47_410 VPWR VGND sg13g2_decap_8
XFILLER_47_487 VPWR VGND sg13g2_decap_8
XFILLER_35_638 VPWR VGND sg13g2_decap_8
XFILLER_34_126 VPWR VGND sg13g2_fill_1
XFILLER_34_148 VPWR VGND sg13g2_fill_2
XFILLER_16_863 VPWR VGND sg13g2_decap_8
XFILLER_37_1013 VPWR VGND sg13g2_decap_8
XFILLER_43_682 VPWR VGND sg13g2_decap_8
X_2880_ sap_3_inst.alu_inst.tmp\[1\] _0363_ net790 _0383_ VPWR VGND sg13g2_nand3_1
XFILLER_31_866 VPWR VGND sg13g2_decap_8
XFILLER_7_583 VPWR VGND sg13g2_decap_8
X_3501_ net573 _0950_ _0968_ VPWR VGND sg13g2_xor2_1
X_3432_ VGND VPWR net664 _0900_ _0902_ net587 sg13g2_a21oi_1
X_3363_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[2\] net670 _0834_
+ VPWR VGND sg13g2_and2_1
XFILLER_39_900 VPWR VGND sg13g2_decap_8
X_2314_ _1581_ _1611_ _1731_ VPWR VGND sg13g2_nor2_2
X_3294_ net689 _0749_ _0765_ VPWR VGND sg13g2_nor2_1
X_2245_ VGND VPWR _1662_ _1641_ _1573_ sg13g2_or2_1
XFILLER_39_977 VPWR VGND sg13g2_decap_8
X_2176_ net730 _1592_ _1593_ VPWR VGND sg13g2_and2_1
XFILLER_25_126 VPWR VGND sg13g2_fill_2
XFILLER_25_148 VPWR VGND sg13g2_fill_1
XFILLER_26_649 VPWR VGND sg13g2_decap_8
XFILLER_22_844 VPWR VGND sg13g2_decap_8
XFILLER_34_682 VPWR VGND sg13g2_decap_8
Xoutput15 net15 uio_oe[6] VPWR VGND sg13g2_buf_1
Xoutput26 net26 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_737 VPWR VGND sg13g2_decap_8
XFILLER_45_925 VPWR VGND sg13g2_decap_8
XFILLER_44_435 VPWR VGND sg13g2_decap_8
XFILLER_25_660 VPWR VGND sg13g2_decap_8
XFILLER_13_844 VPWR VGND sg13g2_decap_8
XFILLER_40_674 VPWR VGND sg13g2_decap_8
XFILLER_9_837 VPWR VGND sg13g2_decap_8
XFILLER_21_70 VPWR VGND sg13g2_fill_1
XFILLER_4_564 VPWR VGND sg13g2_decap_8
XFILLER_39_207 VPWR VGND sg13g2_fill_1
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_48_752 VPWR VGND sg13g2_decap_8
XFILLER_36_925 VPWR VGND sg13g2_decap_8
XFILLER_16_660 VPWR VGND sg13g2_decap_8
X_3981_ _1357_ _1350_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[0\]
+ _1348_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2932_ net693 _0432_ _0434_ VPWR VGND sg13g2_nor2_1
XFILLER_31_663 VPWR VGND sg13g2_decap_8
X_2863_ _0367_ _0345_ _0349_ _0343_ _1487_ VPWR VGND sg13g2_a22oi_1
X_2794_ _1702_ _1711_ _0307_ _0308_ VPWR VGND sg13g2_nor3_1
XFILLER_8_892 VPWR VGND sg13g2_decap_8
XFILLER_11_1027 VPWR VGND sg13g2_fill_2
Xfanout805 net806 net805 VPWR VGND sg13g2_buf_8
X_3415_ _0885_ net683 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[1\]
+ net688 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[1\] VPWR VGND sg13g2_a22oi_1
Xfanout816 net836 net816 VPWR VGND sg13g2_buf_8
X_3346_ _0817_ net681 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[0\]
+ net687 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[0\] VPWR VGND sg13g2_a22oi_1
Xfanout827 net829 net827 VPWR VGND sg13g2_buf_8
X_3277_ _0653_ _0665_ _0748_ VPWR VGND sg13g2_nor2_2
XFILLER_27_903 VPWR VGND sg13g2_decap_8
X_2228_ _1574_ _1623_ _1645_ VPWR VGND sg13g2_and2_1
XFILLER_39_774 VPWR VGND sg13g2_decap_8
X_2159_ VGND VPWR _1576_ net770 net767 sg13g2_or2_1
XFILLER_26_446 VPWR VGND sg13g2_decap_8
XFILLER_22_641 VPWR VGND sg13g2_decap_8
XFILLER_10_814 VPWR VGND sg13g2_decap_8
XFILLER_5_328 VPWR VGND sg13g2_fill_2
XFILLER_1_534 VPWR VGND sg13g2_decap_8
XFILLER_27_1001 VPWR VGND sg13g2_decap_8
XFILLER_49_538 VPWR VGND sg13g2_decap_8
XFILLER_45_722 VPWR VGND sg13g2_decap_8
XFILLER_18_914 VPWR VGND sg13g2_decap_8
XFILLER_44_210 VPWR VGND sg13g2_fill_1
XFILLER_32_405 VPWR VGND sg13g2_fill_2
XFILLER_45_799 VPWR VGND sg13g2_decap_8
XFILLER_44_298 VPWR VGND sg13g2_fill_2
XFILLER_33_939 VPWR VGND sg13g2_decap_8
XFILLER_41_950 VPWR VGND sg13g2_decap_8
XFILLER_13_641 VPWR VGND sg13g2_decap_8
XFILLER_40_471 VPWR VGND sg13g2_decap_8
XFILLER_9_634 VPWR VGND sg13g2_decap_8
XFILLER_12_195 VPWR VGND sg13g2_fill_1
XFILLER_5_884 VPWR VGND sg13g2_decap_8
X_3200_ _0671_ _1587_ _1679_ VPWR VGND sg13g2_nand2_1
X_4180_ net823 VGND VPWR _0037_ sap_3_inst.alu_inst.acc\[4\] clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3131_ _0616_ VPWR _0051_ VGND _2051_ net701 sg13g2_o21ai_1
X_3062_ _0559_ VPWR _0560_ VGND _0349_ _0553_ sg13g2_o21ai_1
XFILLER_36_722 VPWR VGND sg13g2_decap_8
XFILLER_24_906 VPWR VGND sg13g2_decap_8
XFILLER_23_438 VPWR VGND sg13g2_decap_8
XFILLER_36_799 VPWR VGND sg13g2_decap_8
X_3964_ _1335_ _1339_ _1340_ VPWR VGND sg13g2_nor2_2
X_3895_ VPWR _1286_ _1285_ VGND sg13g2_inv_1
X_2915_ _0415_ _0416_ _0417_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_994 VPWR VGND sg13g2_decap_8
X_2846_ _0350_ _0346_ _0349_ VPWR VGND sg13g2_nand2_1
X_2777_ _0004_ _1682_ _0297_ _0300_ VPWR VGND sg13g2_and3_1
Xfanout613 _0745_ net613 VPWR VGND sg13g2_buf_1
Xfanout624 _1852_ net624 VPWR VGND sg13g2_buf_8
Xfanout602 net603 net602 VPWR VGND sg13g2_buf_8
Xfanout646 _0760_ net646 VPWR VGND sg13g2_buf_8
Xfanout635 _1233_ net635 VPWR VGND sg13g2_buf_8
Xfanout657 _0751_ net657 VPWR VGND sg13g2_buf_8
X_3329_ _0800_ net640 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[4\]
+ net641 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[4\] VPWR VGND sg13g2_a22oi_1
Xfanout679 _0753_ net679 VPWR VGND sg13g2_buf_8
Xfanout668 _0874_ net668 VPWR VGND sg13g2_buf_8
XFILLER_27_700 VPWR VGND sg13g2_decap_8
XFILLER_39_571 VPWR VGND sg13g2_decap_8
XFILLER_15_917 VPWR VGND sg13g2_decap_8
XFILLER_26_254 VPWR VGND sg13g2_decap_4
XFILLER_27_777 VPWR VGND sg13g2_decap_8
XFILLER_42_758 VPWR VGND sg13g2_decap_8
XFILLER_10_611 VPWR VGND sg13g2_decap_8
XFILLER_6_659 VPWR VGND sg13g2_decap_8
XFILLER_10_688 VPWR VGND sg13g2_decap_8
XFILLER_2_876 VPWR VGND sg13g2_decap_8
XFILLER_49_335 VPWR VGND sg13g2_decap_8
XFILLER_18_711 VPWR VGND sg13g2_decap_8
XFILLER_18_788 VPWR VGND sg13g2_decap_8
XFILLER_45_596 VPWR VGND sg13g2_decap_8
XFILLER_33_736 VPWR VGND sg13g2_decap_8
XFILLER_21_909 VPWR VGND sg13g2_decap_8
XFILLER_14_961 VPWR VGND sg13g2_decap_8
X_2700_ net793 net791 _0231_ VPWR VGND sg13g2_xor2_1
X_3680_ net636 _1128_ _1129_ _1130_ VPWR VGND sg13g2_nor3_1
X_2631_ net2 _1884_ _2040_ VPWR VGND sg13g2_and2_1
X_2562_ _1973_ net616 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[4\]
+ net628 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_681 VPWR VGND sg13g2_decap_8
X_4301_ net834 VGND VPWR _0158_ sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[2\]
+ clknet_3_6__leaf_clk sg13g2_dfrbpq_2
X_4232_ net809 VGND VPWR _0089_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[7\]
+ clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_2493_ _1910_ net616 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[7\]
+ net624 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_4_95 VPWR VGND sg13g2_fill_2
X_4163_ net818 VGND VPWR _0024_ u_ser.shadow_reg\[7\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
X_3114_ _0542_ _0573_ _0459_ _0602_ VPWR VGND _0601_ sg13g2_nand4_1
X_4148__6 VPWR net40 clknet_leaf_0_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
X_4094_ _1451_ VPWR _0179_ VGND net578 _1450_ sg13g2_o21ai_1
XFILLER_28_519 VPWR VGND sg13g2_decap_8
X_3045_ _0333_ _0542_ _2012_ _0543_ VPWR VGND sg13g2_nand3_1
XFILLER_24_703 VPWR VGND sg13g2_decap_8
XFILLER_36_596 VPWR VGND sg13g2_decap_8
X_3947_ net70 _0155_ _1324_ VPWR VGND sg13g2_nor2_1
XFILLER_20_931 VPWR VGND sg13g2_decap_8
XFILLER_32_791 VPWR VGND sg13g2_decap_8
X_3878_ net654 _1057_ _1058_ _1277_ VPWR VGND sg13g2_nor3_1
X_2829_ _2016_ _2018_ _0333_ VPWR VGND sg13g2_nor2_2
XFILLER_3_8 VPWR VGND sg13g2_fill_2
XFILLER_24_1004 VPWR VGND sg13g2_decap_8
XFILLER_46_349 VPWR VGND sg13g2_decap_8
XFILLER_15_714 VPWR VGND sg13g2_decap_8
XFILLER_27_574 VPWR VGND sg13g2_decap_8
XFILLER_42_555 VPWR VGND sg13g2_decap_8
XFILLER_14_279 VPWR VGND sg13g2_fill_1
XFILLER_30_728 VPWR VGND sg13g2_decap_8
XFILLER_11_964 VPWR VGND sg13g2_decap_8
XFILLER_7_968 VPWR VGND sg13g2_decap_8
XFILLER_10_485 VPWR VGND sg13g2_decap_8
XFILLER_6_456 VPWR VGND sg13g2_decap_8
XFILLER_2_673 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_fill_1
XFILLER_37_305 VPWR VGND sg13g2_fill_1
XFILLER_38_839 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_18_585 VPWR VGND sg13g2_decap_8
XFILLER_45_393 VPWR VGND sg13g2_decap_8
XFILLER_33_533 VPWR VGND sg13g2_decap_8
XFILLER_21_706 VPWR VGND sg13g2_decap_8
X_3801_ VGND VPWR net607 _0901_ _1223_ net657 sg13g2_a21oi_1
X_3732_ _1170_ net594 _0894_ VPWR VGND sg13g2_nand2b_1
Xclkload20 VPWR clkload20/Y clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs VGND sg13g2_inv_1
X_3663_ VPWR VGND net595 _0766_ _0951_ _0857_ _1115_ _0945_ sg13g2_a221oi_1
X_2614_ _2011_ _2022_ _2023_ VPWR VGND sg13g2_nor2b_1
X_3594_ net31 _1055_ _1056_ _1057_ VPWR VGND sg13g2_nor3_2
XFILLER_47_1026 VPWR VGND sg13g2_fill_2
X_2545_ net6 _1884_ _1958_ VPWR VGND sg13g2_and2_1
X_2476_ net729 _1616_ _1893_ VPWR VGND sg13g2_nor2_1
X_4215_ net810 VGND VPWR _0072_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[6\]
+ clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_1
XFILLER_29_817 VPWR VGND sg13g2_decap_8
X_4077_ _1436_ VPWR _0176_ VGND _1090_ _1437_ sg13g2_o21ai_1
X_3028_ _0527_ _0525_ _0526_ VPWR VGND sg13g2_nand2_1
XFILLER_24_500 VPWR VGND sg13g2_decap_8
XFILLER_37_894 VPWR VGND sg13g2_decap_8
XFILLER_24_577 VPWR VGND sg13g2_decap_8
XFILLER_34_59 VPWR VGND sg13g2_fill_2
Xclkload3 clknet_3_4__leaf_clk clkload3/X VPWR VGND sg13g2_buf_1
XFILLER_4_949 VPWR VGND sg13g2_decap_8
XFILLER_3_448 VPWR VGND sg13g2_decap_8
XFILLER_47_669 VPWR VGND sg13g2_decap_8
XFILLER_15_511 VPWR VGND sg13g2_decap_8
XFILLER_28_883 VPWR VGND sg13g2_decap_8
XFILLER_43_864 VPWR VGND sg13g2_decap_8
XFILLER_15_588 VPWR VGND sg13g2_decap_8
XFILLER_42_374 VPWR VGND sg13g2_fill_1
XFILLER_30_525 VPWR VGND sg13g2_decap_8
XFILLER_11_761 VPWR VGND sg13g2_decap_8
XFILLER_24_81 VPWR VGND sg13g2_fill_1
XFILLER_24_92 VPWR VGND sg13g2_fill_2
XFILLER_7_765 VPWR VGND sg13g2_decap_8
X_2330_ _1747_ net735 _1637_ VPWR VGND sg13g2_nand2b_1
X_2261_ net714 _1675_ _1677_ _1678_ VPWR VGND sg13g2_or3_1
XFILLER_2_470 VPWR VGND sg13g2_decap_8
XFILLER_27_4 VPWR VGND sg13g2_fill_2
X_4000_ _1374_ _1349_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[2\]
+ net796 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2192_ _1560_ net751 _1571_ _1609_ VPWR VGND sg13g2_or3_1
XFILLER_38_636 VPWR VGND sg13g2_decap_8
XFILLER_19_861 VPWR VGND sg13g2_decap_8
XFILLER_37_146 VPWR VGND sg13g2_fill_1
XFILLER_21_503 VPWR VGND sg13g2_decap_8
XFILLER_34_864 VPWR VGND sg13g2_decap_8
XFILLER_14_1003 VPWR VGND sg13g2_decap_8
X_3715_ _1069_ _1071_ _1159_ VPWR VGND sg13g2_nor2_2
X_3646_ _1099_ _1100_ _1095_ _1101_ VPWR VGND sg13g2_nand3_1
X_3577_ _1040_ _1025_ _1041_ VPWR VGND sg13g2_xor2_1
XFILLER_1_919 VPWR VGND sg13g2_decap_8
X_2528_ sap_3_inst.alu_flags\[6\] net710 _1942_ VPWR VGND sg13g2_nor2_1
X_2459_ _1876_ _1703_ _1731_ _1699_ _1684_ VPWR VGND sg13g2_a22oi_1
XFILLER_29_37 VPWR VGND sg13g2_fill_1
Xhold26 sap_3_inst.reg_file_inst.array_serializer_inst.state\[1\] VPWR VGND net73
+ sg13g2_dlygate4sd3_1
Xhold15 _1321_ VPWR VGND net62 sg13g2_dlygate4sd3_1
XFILLER_21_1007 VPWR VGND sg13g2_decap_8
XFILLER_28_102 VPWR VGND sg13g2_fill_2
XFILLER_29_614 VPWR VGND sg13g2_decap_8
X_4129_ net64 u_ser.state\[1\] net799 _0188_ VPWR VGND sg13g2_a21o_1
XFILLER_44_617 VPWR VGND sg13g2_decap_8
XFILLER_25_842 VPWR VGND sg13g2_decap_8
XFILLER_37_691 VPWR VGND sg13g2_decap_8
XFILLER_40_856 VPWR VGND sg13g2_decap_8
XFILLER_8_507 VPWR VGND sg13g2_decap_8
XFILLER_12_569 VPWR VGND sg13g2_decap_8
XFILLER_3_201 VPWR VGND sg13g2_fill_1
XFILLER_4_746 VPWR VGND sg13g2_decap_8
XFILLER_0_952 VPWR VGND sg13g2_decap_8
XFILLER_48_934 VPWR VGND sg13g2_decap_8
XFILLER_47_466 VPWR VGND sg13g2_decap_8
XFILLER_35_617 VPWR VGND sg13g2_decap_8
XFILLER_16_842 VPWR VGND sg13g2_decap_8
XFILLER_28_680 VPWR VGND sg13g2_decap_8
XFILLER_43_661 VPWR VGND sg13g2_decap_8
XFILLER_31_845 VPWR VGND sg13g2_decap_8
X_3500_ _0966_ VPWR _0967_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[4\]
+ net661 sg13g2_o21ai_1
XFILLER_7_562 VPWR VGND sg13g2_decap_8
X_3431_ VPWR _0901_ _0900_ VGND sg13g2_inv_1
X_3362_ _1505_ net690 _0749_ _0833_ VPWR VGND sg13g2_nor3_1
X_2313_ net764 _1660_ _1685_ _1730_ VPWR VGND sg13g2_nor3_2
X_3293_ _0764_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[0\] net670
+ VPWR VGND sg13g2_nand2_1
X_2244_ _1573_ _1641_ _1661_ VPWR VGND sg13g2_nor2_1
XFILLER_39_956 VPWR VGND sg13g2_decap_8
X_2175_ _1494_ _1560_ _1571_ _1592_ VGND VPWR _1576_ sg13g2_nor4_2
XFILLER_18_0 VPWR VGND sg13g2_fill_1
XFILLER_26_628 VPWR VGND sg13g2_decap_8
XFILLER_34_661 VPWR VGND sg13g2_decap_8
XFILLER_22_823 VPWR VGND sg13g2_decap_8
XFILLER_31_49 VPWR VGND sg13g2_fill_2
X_3629_ net584 _1084_ _1086_ VPWR VGND sg13g2_nor2_1
XFILLER_1_716 VPWR VGND sg13g2_decap_8
Xoutput27 net27 uo_out[2] VPWR VGND sg13g2_buf_1
Xoutput16 net16 uio_oe[7] VPWR VGND sg13g2_buf_1
XFILLER_45_904 VPWR VGND sg13g2_decap_8
XFILLER_44_414 VPWR VGND sg13g2_decap_8
Xclk_div_param_inst__2_ net808 VGND VPWR net35 clk_div_out clknet_3_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_29_488 VPWR VGND sg13g2_decap_8
XFILLER_17_639 VPWR VGND sg13g2_decap_8
XFILLER_32_609 VPWR VGND sg13g2_decap_8
XFILLER_13_823 VPWR VGND sg13g2_decap_8
XFILLER_40_653 VPWR VGND sg13g2_decap_8
XFILLER_9_816 VPWR VGND sg13g2_decap_8
XFILLER_4_543 VPWR VGND sg13g2_decap_8
Xclkbuf_4_0_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_0_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_48_731 VPWR VGND sg13g2_decap_8
XFILLER_36_904 VPWR VGND sg13g2_decap_8
XFILLER_47_252 VPWR VGND sg13g2_fill_1
XFILLER_46_90 VPWR VGND sg13g2_fill_2
X_3980_ _1356_ _1346_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[0\]
+ _1340_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_44_981 VPWR VGND sg13g2_decap_8
X_2931_ _0433_ sap_3_inst.alu_inst.act\[2\] net702 VPWR VGND sg13g2_nand2_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_642 VPWR VGND sg13g2_decap_8
X_2862_ _0366_ net748 _0342_ VPWR VGND sg13g2_nand2_1
X_2793_ _1651_ _1659_ _1674_ _0307_ VPWR VGND sg13g2_nor3_1
XFILLER_30_196 VPWR VGND sg13g2_fill_1
XFILLER_8_871 VPWR VGND sg13g2_decap_8
XFILLER_11_1006 VPWR VGND sg13g2_decap_8
X_3414_ _0884_ net660 _0883_ VPWR VGND sg13g2_nand2_1
Xfanout806 net807 net806 VPWR VGND sg13g2_buf_8
Xfanout817 net818 net817 VPWR VGND sg13g2_buf_8
X_3345_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[0\] net673 _0816_
+ VPWR VGND sg13g2_and2_1
Xfanout828 net832 net828 VPWR VGND sg13g2_buf_8
X_3276_ _0652_ _0664_ _0708_ _0747_ VPWR VGND sg13g2_nor3_1
X_2227_ _1575_ net749 _1641_ _1644_ VPWR VGND sg13g2_or3_1
XFILLER_39_753 VPWR VGND sg13g2_decap_8
XFILLER_38_263 VPWR VGND sg13g2_fill_2
X_2158_ VGND VPWR _1575_ net757 net760 sg13g2_or2_1
XFILLER_26_425 VPWR VGND sg13g2_decap_8
XFILLER_27_959 VPWR VGND sg13g2_decap_8
X_2089_ VPWR _1507_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[2\]
+ VGND sg13g2_inv_1
XFILLER_13_119 VPWR VGND sg13g2_fill_2
XFILLER_22_620 VPWR VGND sg13g2_decap_8
XFILLER_35_981 VPWR VGND sg13g2_decap_8
XFILLER_22_697 VPWR VGND sg13g2_decap_8
XFILLER_1_513 VPWR VGND sg13g2_decap_8
XFILLER_49_517 VPWR VGND sg13g2_decap_8
XFILLER_45_701 VPWR VGND sg13g2_decap_8
XFILLER_17_436 VPWR VGND sg13g2_fill_2
XFILLER_45_778 VPWR VGND sg13g2_decap_8
XFILLER_33_918 VPWR VGND sg13g2_decap_8
XFILLER_26_992 VPWR VGND sg13g2_decap_8
XFILLER_13_620 VPWR VGND sg13g2_decap_8
XFILLER_9_613 VPWR VGND sg13g2_decap_8
XFILLER_13_697 VPWR VGND sg13g2_decap_8
XFILLER_5_863 VPWR VGND sg13g2_decap_8
X_4155__13 VPWR net47 clknet_leaf_1_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
X_3130_ _0616_ sap_3_inst.alu_inst.tmp\[1\] net700 VPWR VGND sg13g2_nand2_1
X_3061_ _0559_ _0557_ _0558_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_701 VPWR VGND sg13g2_decap_8
XFILLER_36_778 VPWR VGND sg13g2_decap_8
X_3963_ _1339_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[1\] VPWR
+ VGND sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[0\] sg13g2_nand2b_2
X_2914_ _0375_ _0405_ _0373_ _0416_ VPWR VGND sg13g2_nand3_1
X_3894_ _1285_ _0719_ net648 VPWR VGND sg13g2_nand2_2
XFILLER_32_973 VPWR VGND sg13g2_decap_8
X_2845_ VGND VPWR _0349_ _2054_ _2010_ sg13g2_or2_1
X_2776_ _0300_ _1681_ net744 VPWR VGND sg13g2_nand2b_1
Xfanout603 _1164_ net603 VPWR VGND sg13g2_buf_8
Xfanout614 net615 net614 VPWR VGND sg13g2_buf_8
X_3328_ _0795_ _0796_ _0797_ _0798_ _0799_ VPWR VGND sg13g2_and4_1
Xfanout647 net648 net647 VPWR VGND sg13g2_buf_8
Xfanout658 _0751_ net658 VPWR VGND sg13g2_buf_2
Xfanout625 _1852_ net625 VPWR VGND sg13g2_buf_8
Xfanout636 net637 net636 VPWR VGND sg13g2_buf_8
Xfanout669 net670 net669 VPWR VGND sg13g2_buf_8
X_3259_ _0728_ _0729_ _0730_ VPWR VGND sg13g2_and2_1
XFILLER_39_550 VPWR VGND sg13g2_decap_8
XFILLER_27_756 VPWR VGND sg13g2_decap_8
XFILLER_42_737 VPWR VGND sg13g2_decap_8
XFILLER_14_439 VPWR VGND sg13g2_fill_2
XFILLER_41_269 VPWR VGND sg13g2_fill_2
XFILLER_23_984 VPWR VGND sg13g2_decap_8
XFILLER_22_494 VPWR VGND sg13g2_decap_8
XFILLER_10_667 VPWR VGND sg13g2_decap_8
XFILLER_6_638 VPWR VGND sg13g2_decap_8
XFILLER_2_855 VPWR VGND sg13g2_decap_8
XFILLER_1_332 VPWR VGND sg13g2_fill_1
XFILLER_49_314 VPWR VGND sg13g2_decap_8
XFILLER_40_1010 VPWR VGND sg13g2_decap_8
XFILLER_37_509 VPWR VGND sg13g2_decap_8
XFILLER_18_767 VPWR VGND sg13g2_decap_8
XFILLER_45_575 VPWR VGND sg13g2_decap_8
XFILLER_33_715 VPWR VGND sg13g2_decap_8
XFILLER_14_940 VPWR VGND sg13g2_decap_8
XFILLER_13_494 VPWR VGND sg13g2_decap_8
X_2630_ VGND VPWR net695 _2038_ _2039_ _2037_ sg13g2_a21oi_1
XFILLER_9_487 VPWR VGND sg13g2_decap_8
X_2561_ _1972_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[4\] net601
+ VPWR VGND sg13g2_nand2_1
XFILLER_5_660 VPWR VGND sg13g2_decap_8
X_2492_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[7\] net620
+ net600 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[7\] _1909_ net711
+ sg13g2_a221oi_1
X_4300_ net834 VGND VPWR net55 sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[1\]
+ clknet_3_6__leaf_clk sg13g2_dfrbpq_2
X_4231_ net812 VGND VPWR _0088_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[6\]
+ clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4162_ net821 VGND VPWR _0023_ u_ser.shadow_reg\[6\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
X_3113_ _0475_ _0508_ _0601_ VPWR VGND sg13g2_and2_1
X_4093_ _1451_ sap_3_inst.alu_inst.act\[2\] net578 VPWR VGND sg13g2_nand2_1
XFILLER_49_881 VPWR VGND sg13g2_decap_8
X_3044_ sap_3_inst.alu_inst.tmp\[6\] net775 _0542_ VPWR VGND sg13g2_xor2_1
XFILLER_36_575 VPWR VGND sg13g2_decap_8
XFILLER_23_236 VPWR VGND sg13g2_fill_1
XFILLER_24_759 VPWR VGND sg13g2_decap_8
XFILLER_20_910 VPWR VGND sg13g2_decap_8
X_3946_ regFile_serial_start net73 _0154_ _0159_ VPWR VGND sg13g2_a21o_1
XFILLER_32_770 VPWR VGND sg13g2_decap_8
X_3877_ _1272_ VPWR _0137_ VGND _1275_ _1276_ sg13g2_o21ai_1
X_2828_ _0332_ _2002_ _0331_ VPWR VGND sg13g2_nand2_1
XFILLER_20_987 VPWR VGND sg13g2_decap_8
X_2759_ _1707_ _0281_ _0284_ _0285_ _0286_ VPWR VGND sg13g2_nor4_1
XFILLER_2_129 VPWR VGND sg13g2_fill_1
Xclkbuf_5_31__f_sap_3_inst.alu_inst.clk_regs clknet_4_15_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_48_36 VPWR VGND sg13g2_fill_1
XFILLER_27_553 VPWR VGND sg13g2_decap_8
XFILLER_42_534 VPWR VGND sg13g2_decap_8
XFILLER_30_707 VPWR VGND sg13g2_decap_8
XFILLER_11_943 VPWR VGND sg13g2_decap_8
XFILLER_23_781 VPWR VGND sg13g2_decap_8
XFILLER_10_431 VPWR VGND sg13g2_fill_1
XFILLER_7_947 VPWR VGND sg13g2_decap_8
Xclkbuf_5_20__f_sap_3_inst.alu_inst.clk_regs clknet_4_10_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_2_652 VPWR VGND sg13g2_decap_8
XFILLER_29_8 VPWR VGND sg13g2_fill_1
XFILLER_38_818 VPWR VGND sg13g2_decap_8
XFILLER_46_895 VPWR VGND sg13g2_decap_8
XFILLER_45_372 VPWR VGND sg13g2_decap_8
XFILLER_18_564 VPWR VGND sg13g2_decap_8
XFILLER_33_512 VPWR VGND sg13g2_decap_8
X_3800_ net587 _0900_ _1222_ VPWR VGND sg13g2_nor2_1
XFILLER_33_589 VPWR VGND sg13g2_decap_8
X_3731_ _1169_ VPWR _0098_ VGND _1521_ net677 sg13g2_o21ai_1
Xclkload10 VPWR clkload10/Y clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs VGND sg13g2_inv_1
X_3662_ _1113_ VPWR _1114_ VGND _0303_ net668 sg13g2_o21ai_1
X_2613_ VGND VPWR _2008_ _2020_ _2022_ _2021_ sg13g2_a21oi_1
X_4150__8 VPWR net42 clknet_leaf_2_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
X_3593_ VGND VPWR _0720_ net589 _1056_ net659 sg13g2_a21oi_1
X_2544_ VGND VPWR net695 _1956_ _1957_ _1955_ sg13g2_a21oi_1
XFILLER_47_1005 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_2475_ _1891_ VPWR _1892_ VGND _1601_ _1886_ sg13g2_o21ai_1
X_4214_ net809 VGND VPWR _0071_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[5\]
+ clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4076_ _1437_ net651 _1091_ VPWR VGND sg13g2_nand2_1
X_3027_ _0526_ _0359_ net775 net692 net781 VPWR VGND sg13g2_a22oi_1
XFILLER_37_873 VPWR VGND sg13g2_decap_8
XFILLER_24_556 VPWR VGND sg13g2_decap_8
XFILLER_11_239 VPWR VGND sg13g2_fill_2
X_3929_ _0153_ _1145_ _1312_ net643 _1546_ VPWR VGND sg13g2_a22oi_1
Xclkload4 VPWR clkload4/Y clknet_3_5__leaf_clk VGND sg13g2_inv_1
XFILLER_20_784 VPWR VGND sg13g2_decap_8
XFILLER_4_928 VPWR VGND sg13g2_decap_8
Xclkbuf_5_9__f_sap_3_inst.alu_inst.clk_regs clknet_4_4_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_47_648 VPWR VGND sg13g2_decap_8
XFILLER_46_103 VPWR VGND sg13g2_fill_2
XFILLER_28_862 VPWR VGND sg13g2_decap_8
XFILLER_43_843 VPWR VGND sg13g2_decap_8
XFILLER_15_567 VPWR VGND sg13g2_decap_8
XFILLER_30_504 VPWR VGND sg13g2_decap_8
XFILLER_11_740 VPWR VGND sg13g2_decap_8
XFILLER_7_744 VPWR VGND sg13g2_decap_8
XFILLER_3_994 VPWR VGND sg13g2_decap_8
X_2260_ VGND VPWR net724 _1673_ _1677_ _1644_ sg13g2_a21oi_1
X_2191_ _1560_ _1607_ _1608_ VPWR VGND sg13g2_nor2_1
XFILLER_38_615 VPWR VGND sg13g2_decap_8
XFILLER_19_840 VPWR VGND sg13g2_decap_8
XFILLER_46_692 VPWR VGND sg13g2_decap_8
XFILLER_34_843 VPWR VGND sg13g2_decap_8
XFILLER_21_559 VPWR VGND sg13g2_decap_8
X_3714_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[3\] _1147_ _1158_
+ VPWR VGND sg13g2_nor2_1
X_3645_ _1100_ net637 _1055_ VPWR VGND sg13g2_nand2_1
X_3576_ _1040_ _1037_ _1039_ net664 _1545_ VPWR VGND sg13g2_a22oi_1
X_2527_ net23 net570 VPWR VGND sg13g2_inv_2
X_2458_ _1554_ net751 _1571_ _1875_ VGND VPWR _1611_ sg13g2_nor4_2
Xhold16 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[4\] VPWR VGND net63
+ sg13g2_dlygate4sd3_1
Xhold27 _0159_ VPWR VGND net74 sg13g2_dlygate4sd3_1
X_2389_ _1806_ _1804_ _1805_ net714 _1637_ VPWR VGND sg13g2_a22oi_1
X_4128_ VPWR _0187_ _1478_ VGND sg13g2_inv_1
XFILLER_28_136 VPWR VGND sg13g2_fill_2
X_4059_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[7\] _1427_
+ _1350_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[7\] _1428_ net796
+ sg13g2_a221oi_1
XFILLER_37_670 VPWR VGND sg13g2_decap_8
XFILLER_24_320 VPWR VGND sg13g2_fill_1
XFILLER_25_821 VPWR VGND sg13g2_decap_8
XFILLER_40_835 VPWR VGND sg13g2_decap_8
XFILLER_25_898 VPWR VGND sg13g2_decap_8
XFILLER_12_548 VPWR VGND sg13g2_decap_8
XFILLER_20_581 VPWR VGND sg13g2_decap_8
XFILLER_4_725 VPWR VGND sg13g2_decap_8
XFILLER_10_84 VPWR VGND sg13g2_fill_1
XFILLER_0_931 VPWR VGND sg13g2_decap_8
XFILLER_48_913 VPWR VGND sg13g2_decap_8
XFILLER_47_445 VPWR VGND sg13g2_decap_8
XFILLER_16_821 VPWR VGND sg13g2_decap_8
XFILLER_43_640 VPWR VGND sg13g2_decap_8
XFILLER_16_898 VPWR VGND sg13g2_decap_8
XFILLER_30_301 VPWR VGND sg13g2_fill_2
XFILLER_31_824 VPWR VGND sg13g2_decap_8
XFILLER_7_541 VPWR VGND sg13g2_decap_8
X_3430_ VGND VPWR _0900_ _0899_ _0898_ sg13g2_or2_1
X_3361_ _1506_ net690 _0746_ _0832_ VPWR VGND sg13g2_nor3_1
X_2312_ net722 VPWR _1729_ VGND net734 _1703_ sg13g2_o21ai_1
XFILLER_3_791 VPWR VGND sg13g2_decap_8
XFILLER_2_290 VPWR VGND sg13g2_fill_2
X_3292_ _0688_ _0689_ _0708_ _0710_ _0763_ VPWR VGND sg13g2_and4_1
XFILLER_39_935 VPWR VGND sg13g2_decap_8
X_2243_ _1572_ _1655_ _1561_ _1660_ VPWR VGND sg13g2_nand3_1
X_2174_ VPWR _1591_ _1590_ VGND sg13g2_inv_1
XFILLER_26_607 VPWR VGND sg13g2_decap_8
XFILLER_38_489 VPWR VGND sg13g2_decap_8
XFILLER_25_128 VPWR VGND sg13g2_fill_1
XFILLER_22_802 VPWR VGND sg13g2_decap_8
XFILLER_34_640 VPWR VGND sg13g2_decap_8
XFILLER_22_879 VPWR VGND sg13g2_decap_8
X_3628_ _1085_ net609 _1022_ VPWR VGND sg13g2_nand2_1
Xoutput17 net31 uio_out[0] VPWR VGND sg13g2_buf_1
Xoutput28 net28 uo_out[3] VPWR VGND sg13g2_buf_1
X_3559_ VGND VPWR net663 _1021_ _1024_ _1023_ sg13g2_a21oi_1
XFILLER_5_1024 VPWR VGND sg13g2_decap_4
XFILLER_17_618 VPWR VGND sg13g2_decap_8
XFILLER_16_128 VPWR VGND sg13g2_fill_1
XFILLER_13_802 VPWR VGND sg13g2_decap_8
XFILLER_25_695 VPWR VGND sg13g2_decap_8
XFILLER_40_632 VPWR VGND sg13g2_decap_8
XFILLER_13_879 VPWR VGND sg13g2_decap_8
XFILLER_4_522 VPWR VGND sg13g2_decap_8
XFILLER_21_50 VPWR VGND sg13g2_fill_2
XFILLER_4_599 VPWR VGND sg13g2_decap_8
XFILLER_48_710 VPWR VGND sg13g2_decap_8
XFILLER_48_787 VPWR VGND sg13g2_decap_8
XFILLER_47_297 VPWR VGND sg13g2_decap_4
XFILLER_44_960 VPWR VGND sg13g2_decap_8
X_2930_ net702 _0430_ _0431_ _0432_ VPWR VGND sg13g2_nor3_1
XFILLER_16_695 VPWR VGND sg13g2_decap_8
XFILLER_31_621 VPWR VGND sg13g2_decap_8
X_2861_ _0362_ _0364_ _0360_ _0365_ VPWR VGND sg13g2_nand3_1
XFILLER_8_850 VPWR VGND sg13g2_decap_8
X_2792_ net741 net731 _1559_ _0000_ VPWR VGND sg13g2_nand3_1
XFILLER_31_698 VPWR VGND sg13g2_decap_8
X_3413_ _0883_ _0848_ _0882_ VPWR VGND sg13g2_nand2_2
Xfanout807 net808 net807 VPWR VGND sg13g2_buf_2
Xfanout818 net826 net818 VPWR VGND sg13g2_buf_8
XFILLER_30_0 VPWR VGND sg13g2_fill_2
X_3344_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[0\] net649 _0815_
+ VPWR VGND sg13g2_and2_1
Xfanout829 net832 net829 VPWR VGND sg13g2_buf_2
X_3275_ _0746_ _0653_ _0665_ VPWR VGND sg13g2_nand2_2
X_2226_ _1575_ net749 _1641_ _1643_ VPWR VGND sg13g2_nor3_1
XFILLER_39_732 VPWR VGND sg13g2_decap_8
X_2157_ net763 net765 net753 _1574_ VGND VPWR net755 sg13g2_nor4_2
XFILLER_27_938 VPWR VGND sg13g2_decap_8
XFILLER_42_919 VPWR VGND sg13g2_decap_8
X_2088_ VPWR _1506_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[2\]
+ VGND sg13g2_inv_1
XFILLER_35_960 VPWR VGND sg13g2_decap_8
XFILLER_22_676 VPWR VGND sg13g2_decap_8
XFILLER_10_849 VPWR VGND sg13g2_decap_8
XFILLER_1_569 VPWR VGND sg13g2_decap_8
XFILLER_18_949 VPWR VGND sg13g2_decap_8
XFILLER_29_286 VPWR VGND sg13g2_fill_1
XFILLER_45_757 VPWR VGND sg13g2_decap_8
XFILLER_26_971 VPWR VGND sg13g2_decap_8
XFILLER_12_120 VPWR VGND sg13g2_fill_1
XFILLER_25_492 VPWR VGND sg13g2_decap_8
XFILLER_41_985 VPWR VGND sg13g2_decap_8
XFILLER_12_142 VPWR VGND sg13g2_fill_1
XFILLER_13_676 VPWR VGND sg13g2_decap_8
XFILLER_34_1018 VPWR VGND sg13g2_decap_8
XFILLER_9_669 VPWR VGND sg13g2_decap_8
XFILLER_32_60 VPWR VGND sg13g2_fill_1
XFILLER_5_842 VPWR VGND sg13g2_decap_8
X_3060_ _0344_ VPWR _0558_ VGND _0520_ _0555_ sg13g2_o21ai_1
XFILLER_48_584 VPWR VGND sg13g2_decap_8
XFILLER_36_757 VPWR VGND sg13g2_decap_8
XFILLER_17_982 VPWR VGND sg13g2_decap_8
X_3962_ net801 net802 _1336_ _1338_ VPWR VGND sg13g2_nor3_1
XFILLER_16_492 VPWR VGND sg13g2_decap_8
XFILLER_32_952 VPWR VGND sg13g2_decap_8
X_3893_ net652 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[7\] _1284_
+ _0145_ VPWR VGND sg13g2_a21o_1
X_2913_ VGND VPWR _0373_ _0375_ _0415_ _0405_ sg13g2_a21oi_1
X_2844_ _2010_ _2054_ _0348_ VPWR VGND sg13g2_nor2_2
XFILLER_31_495 VPWR VGND sg13g2_decap_8
X_2775_ _0299_ _1681_ _0003_ VPWR VGND sg13g2_nor2b_1
Xfanout615 _1864_ net615 VPWR VGND sg13g2_buf_8
Xfanout604 _1096_ net604 VPWR VGND sg13g2_buf_8
X_3327_ _0798_ net678 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[4\]
+ net686 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[4\] VPWR VGND sg13g2_a22oi_1
Xfanout648 net651 net648 VPWR VGND sg13g2_buf_8
Xfanout637 _0766_ net637 VPWR VGND sg13g2_buf_8
Xfanout626 net627 net626 VPWR VGND sg13g2_buf_8
Xfanout659 _0730_ net659 VPWR VGND sg13g2_buf_8
X_3258_ _0729_ _0644_ _1493_ _1586_ _1551_ VPWR VGND sg13g2_a22oi_1
X_2209_ net762 _1625_ _1626_ VPWR VGND sg13g2_nor2_1
XFILLER_2_1027 VPWR VGND sg13g2_fill_2
XFILLER_2_1016 VPWR VGND sg13g2_decap_8
X_3189_ _1659_ VPWR _0660_ VGND net722 _0659_ sg13g2_o21ai_1
XFILLER_27_735 VPWR VGND sg13g2_decap_8
XFILLER_42_716 VPWR VGND sg13g2_decap_8
XFILLER_23_963 VPWR VGND sg13g2_decap_8
XFILLER_22_473 VPWR VGND sg13g2_decap_8
XFILLER_6_617 VPWR VGND sg13g2_decap_8
XFILLER_10_646 VPWR VGND sg13g2_decap_8
XFILLER_2_834 VPWR VGND sg13g2_decap_8
XFILLER_1_300 VPWR VGND sg13g2_fill_2
XFILLER_45_554 VPWR VGND sg13g2_decap_8
XFILLER_18_746 VPWR VGND sg13g2_decap_8
XFILLER_41_782 VPWR VGND sg13g2_decap_8
XFILLER_13_473 VPWR VGND sg13g2_decap_8
XFILLER_14_996 VPWR VGND sg13g2_decap_8
X_2560_ _1971_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[4\] net621
+ VPWR VGND sg13g2_nand2_1
X_2491_ _1908_ _1906_ _1907_ VPWR VGND sg13g2_nand2_1
XFILLER_4_42 VPWR VGND sg13g2_decap_4
X_4230_ net810 VGND VPWR _0087_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[5\]
+ clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4161_ net822 VGND VPWR _0022_ u_ser.shadow_reg\[5\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_4_97 VPWR VGND sg13g2_fill_1
XFILLER_49_860 VPWR VGND sg13g2_decap_8
X_3112_ _0598_ _0577_ _0599_ _0600_ VPWR VGND sg13g2_a21o_1
X_4092_ _1449_ VPWR _1450_ VGND net787 net699 sg13g2_o21ai_1
X_3043_ _0541_ _0363_ _0540_ VPWR VGND sg13g2_nand2_1
XFILLER_48_381 VPWR VGND sg13g2_decap_8
XFILLER_36_554 VPWR VGND sg13g2_decap_8
XFILLER_24_738 VPWR VGND sg13g2_decap_8
XFILLER_17_1024 VPWR VGND sg13g2_decap_4
X_3945_ _0158_ net62 _1322_ VPWR VGND sg13g2_nand2_1
XFILLER_20_966 VPWR VGND sg13g2_decap_8
X_3876_ net671 VPWR _1276_ VGND net587 _1045_ sg13g2_o21ai_1
X_2827_ net703 net694 _0331_ VPWR VGND sg13g2_nor2_1
X_2758_ _1835_ VPWR _0285_ VGND net735 _1682_ sg13g2_o21ai_1
XFILLER_3_609 VPWR VGND sg13g2_decap_8
X_2689_ _0221_ net600 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[2\]
+ net619 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[2\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_27_532 VPWR VGND sg13g2_decap_8
XFILLER_42_513 VPWR VGND sg13g2_decap_8
XFILLER_14_237 VPWR VGND sg13g2_fill_2
XFILLER_15_749 VPWR VGND sg13g2_decap_8
XFILLER_23_760 VPWR VGND sg13g2_decap_8
XFILLER_11_922 VPWR VGND sg13g2_decap_8
XFILLER_7_926 VPWR VGND sg13g2_decap_8
XFILLER_11_999 VPWR VGND sg13g2_decap_8
XFILLER_2_631 VPWR VGND sg13g2_decap_8
XFILLER_18_543 VPWR VGND sg13g2_decap_8
XFILLER_46_874 VPWR VGND sg13g2_decap_8
XFILLER_45_351 VPWR VGND sg13g2_decap_8
XFILLER_33_568 VPWR VGND sg13g2_decap_8
XFILLER_14_793 VPWR VGND sg13g2_decap_8
X_3730_ _0870_ _1168_ net677 _1169_ VPWR VGND sg13g2_nand3_1
X_3661_ VGND VPWR net32 _1097_ _1113_ _0732_ sg13g2_a21oi_1
X_2612_ _2019_ VPWR _2021_ VGND net760 _2013_ sg13g2_o21ai_1
Xclkload11 VPWR clkload11/Y clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs VGND sg13g2_inv_1
X_3592_ net595 net589 _1055_ VPWR VGND sg13g2_and2_1
XFILLER_6_981 VPWR VGND sg13g2_decap_8
X_2543_ _1956_ sap_3_inst.alu_flags\[5\] _1902_ VPWR VGND sg13g2_nand2_1
XFILLER_47_1028 VPWR VGND sg13g2_fill_1
X_2474_ _1887_ _1888_ net716 _1891_ VPWR VGND _1889_ sg13g2_nand4_1
X_4213_ net810 VGND VPWR _0070_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[4\]
+ clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4144_ _0195_ _1490_ _1486_ _1489_ net68 VPWR VGND sg13g2_a22oi_1
XFILLER_18_29 VPWR VGND sg13g2_fill_1
X_4075_ _1436_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[7\] net644
+ VPWR VGND sg13g2_nand2_1
XFILLER_37_852 VPWR VGND sg13g2_decap_8
X_3026_ sap_3_inst.alu_inst.tmp\[5\] _0363_ net778 _0525_ VPWR VGND sg13g2_nand3_1
XFILLER_24_535 VPWR VGND sg13g2_decap_8
X_3928_ net16 net643 _1142_ _1312_ VPWR VGND sg13g2_nor3_1
Xclkload5 VPWR clkload5/Y clknet_3_6__leaf_clk VGND sg13g2_inv_1
X_3859_ net13 _1073_ _1261_ _1262_ VPWR VGND sg13g2_nor3_1
XFILLER_20_763 VPWR VGND sg13g2_decap_8
XFILLER_4_907 VPWR VGND sg13g2_decap_8
XFILLER_3_406 VPWR VGND sg13g2_fill_1
XFILLER_8_1011 VPWR VGND sg13g2_decap_8
XFILLER_47_627 VPWR VGND sg13g2_decap_8
XFILLER_28_841 VPWR VGND sg13g2_decap_8
XFILLER_43_822 VPWR VGND sg13g2_decap_8
XFILLER_15_546 VPWR VGND sg13g2_decap_8
XFILLER_43_899 VPWR VGND sg13g2_decap_8
XFILLER_7_723 VPWR VGND sg13g2_decap_8
XFILLER_11_796 VPWR VGND sg13g2_decap_8
XFILLER_3_973 VPWR VGND sg13g2_decap_8
X_2190_ _1607_ _1570_ VPWR VGND net751 sg13g2_nand2b_2
XFILLER_46_671 VPWR VGND sg13g2_decap_8
XFILLER_37_159 VPWR VGND sg13g2_fill_2
XFILLER_19_896 VPWR VGND sg13g2_decap_8
XFILLER_34_822 VPWR VGND sg13g2_decap_8
XFILLER_21_538 VPWR VGND sg13g2_decap_8
XFILLER_34_899 VPWR VGND sg13g2_decap_8
XFILLER_14_590 VPWR VGND sg13g2_decap_8
X_3713_ VPWR _0092_ _1157_ VGND sg13g2_inv_1
X_3644_ _1098_ VPWR _1099_ VGND net31 net604 sg13g2_o21ai_1
X_3575_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[7\] _1038_
+ net638 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[7\] _1039_ net641
+ sg13g2_a221oi_1
Xclkbuf_4_1_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_1_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2526_ _1941_ _1929_ _1932_ _1940_ VPWR VGND sg13g2_and3_2
X_2457_ _1605_ _1723_ _1874_ VPWR VGND sg13g2_nor2_1
Xhold28 sap_3_outputReg_serial VPWR VGND net75 sg13g2_dlygate4sd3_1
Xhold17 sap_3_outputReg_start_sync VPWR VGND net64 sg13g2_dlygate4sd3_1
X_2388_ net714 _1795_ _1802_ _1803_ _1805_ VPWR VGND sg13g2_nor4_1
X_4127_ _1477_ VPWR _1478_ VGND net75 _0186_ sg13g2_o21ai_1
XFILLER_29_649 VPWR VGND sg13g2_decap_8
XFILLER_25_800 VPWR VGND sg13g2_decap_8
X_4058_ _1424_ _1425_ _1423_ _1427_ VPWR VGND _1426_ sg13g2_nand4_1
XFILLER_43_129 VPWR VGND sg13g2_fill_1
X_3009_ _0506_ _0507_ _0508_ VPWR VGND sg13g2_nor2b_2
XFILLER_24_354 VPWR VGND sg13g2_fill_1
XFILLER_25_877 VPWR VGND sg13g2_decap_8
XFILLER_40_814 VPWR VGND sg13g2_decap_8
XFILLER_12_527 VPWR VGND sg13g2_decap_8
XFILLER_20_560 VPWR VGND sg13g2_decap_8
XFILLER_4_704 VPWR VGND sg13g2_decap_8
XFILLER_10_63 VPWR VGND sg13g2_fill_2
XFILLER_0_910 VPWR VGND sg13g2_decap_8
XFILLER_0_987 VPWR VGND sg13g2_decap_8
XFILLER_48_969 VPWR VGND sg13g2_decap_8
XFILLER_47_424 VPWR VGND sg13g2_decap_8
XFILLER_16_800 VPWR VGND sg13g2_decap_8
XFILLER_16_877 VPWR VGND sg13g2_decap_8
XFILLER_31_803 VPWR VGND sg13g2_decap_8
XFILLER_43_696 VPWR VGND sg13g2_decap_8
XFILLER_30_313 VPWR VGND sg13g2_fill_1
XFILLER_37_1027 VPWR VGND sg13g2_fill_2
XFILLER_7_520 VPWR VGND sg13g2_decap_8
XFILLER_11_593 VPWR VGND sg13g2_decap_8
XFILLER_7_597 VPWR VGND sg13g2_decap_8
X_3360_ _1507_ _0667_ net690 _0831_ VPWR VGND sg13g2_nor3_1
XFILLER_44_1009 VPWR VGND sg13g2_decap_8
XFILLER_3_770 VPWR VGND sg13g2_decap_8
X_2311_ VPWR _1728_ _1727_ VGND sg13g2_inv_1
X_3291_ net689 _0746_ _0762_ VPWR VGND sg13g2_nor2_2
XFILLER_39_914 VPWR VGND sg13g2_decap_8
X_2242_ _1562_ _1573_ _1656_ _1659_ VPWR VGND sg13g2_nor3_2
X_2173_ _1590_ net739 net727 VPWR VGND sg13g2_nand2_1
XFILLER_47_991 VPWR VGND sg13g2_decap_8
XFILLER_19_693 VPWR VGND sg13g2_decap_8
XFILLER_34_696 VPWR VGND sg13g2_decap_8
XFILLER_22_858 VPWR VGND sg13g2_decap_8
X_3627_ _1084_ net570 _1083_ VPWR VGND sg13g2_nand2_1
X_3558_ net609 VPWR _1023_ VGND net663 _1022_ sg13g2_o21ai_1
Xoutput18 net18 uio_out[1] VPWR VGND sg13g2_buf_1
Xoutput29 net29 uo_out[4] VPWR VGND sg13g2_buf_1
X_2509_ _1924_ net616 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[6\]
+ net622 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[6\] VPWR VGND sg13g2_a22oi_1
X_3489_ VGND VPWR _0813_ _0860_ _0957_ _0881_ sg13g2_a21oi_1
XFILLER_5_1003 VPWR VGND sg13g2_decap_8
XFILLER_45_939 VPWR VGND sg13g2_decap_8
XFILLER_44_449 VPWR VGND sg13g2_decap_8
XFILLER_40_611 VPWR VGND sg13g2_decap_8
XFILLER_25_674 VPWR VGND sg13g2_decap_8
XFILLER_13_858 VPWR VGND sg13g2_decap_8
XFILLER_40_688 VPWR VGND sg13g2_decap_8
XFILLER_4_501 VPWR VGND sg13g2_decap_8
XFILLER_4_578 VPWR VGND sg13g2_decap_8
XFILLER_0_784 VPWR VGND sg13g2_decap_8
XFILLER_48_766 VPWR VGND sg13g2_decap_8
XFILLER_36_939 VPWR VGND sg13g2_decap_8
XFILLER_16_674 VPWR VGND sg13g2_decap_8
XFILLER_31_600 VPWR VGND sg13g2_decap_8
XFILLER_43_493 VPWR VGND sg13g2_decap_8
X_2860_ _0364_ _0363_ _0341_ VPWR VGND sg13g2_nand2b_1
XFILLER_15_195 VPWR VGND sg13g2_fill_1
XFILLER_31_677 VPWR VGND sg13g2_decap_8
XFILLER_12_891 VPWR VGND sg13g2_decap_8
X_2791_ net16 _0306_ VPWR VGND sg13g2_inv_2
X_3412_ VGND VPWR _0882_ _0847_ net589 sg13g2_or2_1
Xfanout808 net836 net808 VPWR VGND sg13g2_buf_8
Xfanout819 net826 net819 VPWR VGND sg13g2_buf_8
X_3343_ _0808_ _0809_ _0810_ _0812_ _0814_ VPWR VGND sg13g2_or4_1
XFILLER_23_0 VPWR VGND sg13g2_fill_2
X_3274_ _0745_ _0720_ net659 VPWR VGND sg13g2_nand2_1
XFILLER_39_711 VPWR VGND sg13g2_decap_8
X_2225_ _1575_ _1641_ _1642_ VPWR VGND sg13g2_nor2_1
XFILLER_27_917 VPWR VGND sg13g2_decap_8
XFILLER_39_788 VPWR VGND sg13g2_decap_8
X_2156_ net766 net754 net755 _1573_ VPWR VGND sg13g2_or3_1
XFILLER_19_490 VPWR VGND sg13g2_decap_8
X_2087_ VPWR _1505_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[2\]
+ VGND sg13g2_inv_1
XFILLER_21_110 VPWR VGND sg13g2_fill_1
XFILLER_34_493 VPWR VGND sg13g2_decap_8
XFILLER_22_655 VPWR VGND sg13g2_decap_8
XFILLER_10_828 VPWR VGND sg13g2_decap_8
X_2989_ VGND VPWR _0438_ _0457_ _0489_ _0437_ sg13g2_a21oi_1
XFILLER_1_548 VPWR VGND sg13g2_decap_8
XFILLER_27_1015 VPWR VGND sg13g2_decap_8
XFILLER_45_736 VPWR VGND sg13g2_decap_8
XFILLER_18_928 VPWR VGND sg13g2_decap_8
XFILLER_26_950 VPWR VGND sg13g2_decap_8
XFILLER_29_298 VPWR VGND sg13g2_fill_1
XFILLER_25_471 VPWR VGND sg13g2_decap_8
XFILLER_41_964 VPWR VGND sg13g2_decap_8
XFILLER_13_655 VPWR VGND sg13g2_decap_8
XFILLER_40_485 VPWR VGND sg13g2_decap_8
XFILLER_9_648 VPWR VGND sg13g2_decap_8
XFILLER_12_176 VPWR VGND sg13g2_fill_2
XFILLER_5_821 VPWR VGND sg13g2_decap_8
XFILLER_5_898 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_48_563 VPWR VGND sg13g2_decap_8
XFILLER_36_736 VPWR VGND sg13g2_decap_8
XFILLER_17_961 VPWR VGND sg13g2_decap_8
X_3961_ _1335_ _1336_ _1337_ VPWR VGND sg13g2_nor2_1
X_2912_ _0414_ _0348_ _0413_ VPWR VGND sg13g2_nand2_1
XFILLER_32_931 VPWR VGND sg13g2_decap_8
X_3892_ net652 _1090_ _1092_ _1284_ VPWR VGND sg13g2_nor3_1
X_2843_ VPWR _0347_ _0346_ VGND sg13g2_inv_1
X_2774_ _0297_ VPWR _0299_ VGND net745 _1580_ sg13g2_o21ai_1
Xfanout605 net606 net605 VPWR VGND sg13g2_buf_8
Xfanout649 net651 net649 VPWR VGND sg13g2_buf_8
X_3326_ _0797_ net680 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[4\]
+ net684 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[4\] VPWR VGND sg13g2_a22oi_1
Xfanout627 _1849_ net627 VPWR VGND sg13g2_buf_8
Xfanout616 net617 net616 VPWR VGND sg13g2_buf_8
Xfanout638 net640 net638 VPWR VGND sg13g2_buf_8
X_3257_ _0288_ VPWR _0728_ VGND _0721_ _0727_ sg13g2_o21ai_1
X_2208_ net754 net756 _1625_ VPWR VGND net766 sg13g2_nand3b_1
X_3188_ _1491_ net746 _1493_ _1680_ _0659_ VPWR VGND sg13g2_nor4_1
XFILLER_27_714 VPWR VGND sg13g2_decap_8
XFILLER_39_585 VPWR VGND sg13g2_decap_8
X_2139_ _1552_ _1554_ _1556_ VPWR VGND sg13g2_nor2_2
XFILLER_23_942 VPWR VGND sg13g2_decap_8
XFILLER_22_452 VPWR VGND sg13g2_decap_8
XFILLER_10_625 VPWR VGND sg13g2_decap_8
XFILLER_2_813 VPWR VGND sg13g2_decap_8
XFILLER_49_349 VPWR VGND sg13g2_decap_8
XFILLER_18_725 VPWR VGND sg13g2_decap_8
XFILLER_45_533 VPWR VGND sg13g2_decap_8
XFILLER_32_216 VPWR VGND sg13g2_fill_1
XFILLER_41_761 VPWR VGND sg13g2_decap_8
XFILLER_14_975 VPWR VGND sg13g2_decap_8
Xclkbuf_0_sap_3_inst.alu_inst.clk_regs sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
X_2490_ _1907_ net628 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[7\]
+ net631 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_695 VPWR VGND sg13g2_decap_8
X_4160_ net822 VGND VPWR _0021_ u_ser.shadow_reg\[4\] clknet_3_3__leaf_clk sg13g2_dfrbpq_1
X_3111_ _0587_ VPWR _0599_ VGND net773 _1529_ sg13g2_o21ai_1
X_4091_ _1449_ net698 _0412_ VPWR VGND sg13g2_nand2b_1
XFILLER_48_360 VPWR VGND sg13g2_decap_8
X_3042_ net775 sap_3_inst.alu_inst.tmp\[6\] _0540_ VPWR VGND sg13g2_and2_1
XFILLER_36_533 VPWR VGND sg13g2_decap_8
XFILLER_24_717 VPWR VGND sg13g2_decap_8
XFILLER_17_1003 VPWR VGND sg13g2_decap_8
X_3944_ _1320_ _1323_ _0157_ VPWR VGND sg13g2_nor2_1
X_3875_ net16 net607 _1087_ _1274_ _1275_ VPWR VGND sg13g2_nor4_1
X_2826_ _0329_ VPWR _0330_ VGND net742 _0327_ sg13g2_o21ai_1
XFILLER_20_945 VPWR VGND sg13g2_decap_8
X_2757_ _0283_ VPWR _0284_ VGND _1647_ _1673_ sg13g2_o21ai_1
X_2688_ _0220_ net601 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[2\]
+ net629 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_24_1018 VPWR VGND sg13g2_decap_8
XFILLER_47_809 VPWR VGND sg13g2_decap_8
X_4289_ net828 VGND VPWR _0146_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[0\]
+ clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3309_ _0773_ _0778_ _0772_ _0780_ VPWR VGND sg13g2_nand3_1
XFILLER_27_511 VPWR VGND sg13g2_decap_8
XFILLER_15_728 VPWR VGND sg13g2_decap_8
XFILLER_27_588 VPWR VGND sg13g2_decap_8
XFILLER_42_569 VPWR VGND sg13g2_decap_8
XFILLER_11_901 VPWR VGND sg13g2_decap_8
XFILLER_14_249 VPWR VGND sg13g2_fill_2
Xfanout31 net17 net31 VPWR VGND sg13g2_buf_2
XFILLER_7_905 VPWR VGND sg13g2_decap_8
XFILLER_11_978 VPWR VGND sg13g2_decap_8
XFILLER_6_448 VPWR VGND sg13g2_fill_1
XFILLER_10_499 VPWR VGND sg13g2_decap_8
XFILLER_2_610 VPWR VGND sg13g2_decap_8
XFILLER_2_687 VPWR VGND sg13g2_decap_8
XFILLER_38_60 VPWR VGND sg13g2_fill_2
XFILLER_46_853 VPWR VGND sg13g2_decap_8
XFILLER_18_522 VPWR VGND sg13g2_decap_8
XFILLER_18_599 VPWR VGND sg13g2_decap_8
XFILLER_33_547 VPWR VGND sg13g2_decap_8
XFILLER_14_772 VPWR VGND sg13g2_decap_8
X_3660_ _1112_ VPWR _0084_ VGND _1506_ net639 sg13g2_o21ai_1
X_2611_ _2020_ _1655_ _1996_ VPWR VGND sg13g2_nand2_1
Xclkload12 clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs clkload12/X VPWR VGND sg13g2_buf_1
X_3591_ _1054_ net606 VPWR VGND net642 sg13g2_nand2b_2
XFILLER_6_960 VPWR VGND sg13g2_decap_8
X_2542_ net780 net695 _1955_ VPWR VGND sg13g2_nor2_1
Xclkbuf_5_0__f_sap_3_inst.alu_inst.clk_regs clknet_4_0_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_5_492 VPWR VGND sg13g2_decap_8
X_2473_ VGND VPWR net734 _1684_ _1890_ _1602_ sg13g2_a21oi_1
X_4212_ net828 VGND VPWR _0069_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[3\]
+ clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4143_ net800 _1465_ u_ser.bit_pos\[1\] _1486_ VPWR VGND sg13g2_nand3_1
X_4074_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[6\] _1162_ net647
+ _0175_ VPWR VGND sg13g2_mux2_1
X_3025_ _0524_ _0523_ _0522_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_831 VPWR VGND sg13g2_decap_8
XFILLER_24_514 VPWR VGND sg13g2_decap_8
XFILLER_12_709 VPWR VGND sg13g2_decap_8
X_3927_ VGND VPWR _1540_ net644 _0152_ _1311_ sg13g2_a21oi_1
XFILLER_20_742 VPWR VGND sg13g2_decap_8
X_3858_ net585 _0977_ _1260_ _1261_ VPWR VGND sg13g2_nor3_1
Xclkload6 VPWR clkload6/Y clknet_3_7__leaf_clk VGND sg13g2_inv_1
X_2809_ net56 sap_3_inst.out\[2\] net799 _0019_ VPWR VGND sg13g2_mux2_1
XFILLER_30_1022 VPWR VGND sg13g2_decap_8
X_3789_ _1216_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[3\] net580
+ _0109_ VPWR VGND sg13g2_mux2_1
XFILLER_1_8 VPWR VGND sg13g2_fill_2
XFILLER_47_606 VPWR VGND sg13g2_decap_8
XFILLER_46_116 VPWR VGND sg13g2_fill_2
XFILLER_28_820 VPWR VGND sg13g2_decap_8
XFILLER_43_801 VPWR VGND sg13g2_decap_8
XFILLER_15_525 VPWR VGND sg13g2_decap_8
XFILLER_28_897 VPWR VGND sg13g2_decap_8
XFILLER_43_878 VPWR VGND sg13g2_decap_8
XFILLER_30_539 VPWR VGND sg13g2_decap_8
XFILLER_7_702 VPWR VGND sg13g2_decap_8
XFILLER_11_775 VPWR VGND sg13g2_decap_8
XFILLER_7_779 VPWR VGND sg13g2_decap_8
XFILLER_3_952 VPWR VGND sg13g2_decap_8
XFILLER_2_484 VPWR VGND sg13g2_decap_8
XFILLER_37_127 VPWR VGND sg13g2_fill_2
XFILLER_46_650 VPWR VGND sg13g2_decap_8
XFILLER_1_99 VPWR VGND sg13g2_fill_2
XFILLER_1_66 VPWR VGND sg13g2_decap_8
XFILLER_19_875 VPWR VGND sg13g2_decap_8
XFILLER_34_801 VPWR VGND sg13g2_decap_8
XFILLER_34_878 VPWR VGND sg13g2_decap_8
XFILLER_21_517 VPWR VGND sg13g2_decap_8
XFILLER_14_1017 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
X_3712_ _1157_ _1154_ _1156_ net582 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[2\]
+ VPWR VGND sg13g2_a22oi_1
X_3643_ _1098_ _0301_ _1096_ VPWR VGND sg13g2_nand2_1
X_3574_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[7\] net669 _1038_
+ VPWR VGND sg13g2_and2_1
X_2525_ net576 VPWR _1940_ VGND _1935_ _1939_ sg13g2_o21ai_1
X_2456_ net716 VPWR _1873_ VGND _1660_ _1872_ sg13g2_o21ai_1
Xhold29 u_ser.shadow_reg\[5\] VPWR VGND net76 sg13g2_dlygate4sd3_1
Xhold18 _0188_ VPWR VGND net65 sg13g2_dlygate4sd3_1
X_2387_ _1799_ _1798_ _1804_ VPWR VGND sg13g2_nor2b_1
X_4126_ _1473_ _1475_ _0186_ _1477_ VPWR VGND _1476_ sg13g2_nand4_1
XFILLER_29_628 VPWR VGND sg13g2_decap_8
X_4057_ _1426_ _1352_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[7\]
+ _1346_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3008_ _0507_ net778 sap_3_inst.alu_inst.tmp\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_25_856 VPWR VGND sg13g2_decap_8
XFILLER_12_506 VPWR VGND sg13g2_decap_8
XFILLER_0_966 VPWR VGND sg13g2_decap_8
XFILLER_47_403 VPWR VGND sg13g2_decap_8
XFILLER_48_948 VPWR VGND sg13g2_decap_8
XFILLER_28_694 VPWR VGND sg13g2_decap_8
XFILLER_16_856 VPWR VGND sg13g2_decap_8
XFILLER_37_1006 VPWR VGND sg13g2_decap_8
XFILLER_43_675 VPWR VGND sg13g2_decap_8
XFILLER_31_859 VPWR VGND sg13g2_decap_8
XFILLER_11_572 VPWR VGND sg13g2_decap_8
XFILLER_7_576 VPWR VGND sg13g2_decap_8
X_2310_ _1727_ _1726_ _1694_ VPWR VGND sg13g2_nand2b_1
X_3290_ _0761_ net649 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[0\]
+ net673 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_2_292 VPWR VGND sg13g2_fill_1
X_2241_ VGND VPWR _1656_ _1657_ _1658_ _1654_ sg13g2_a21oi_1
XFILLER_25_4 VPWR VGND sg13g2_fill_2
X_2172_ _1589_ _1578_ _1588_ VPWR VGND sg13g2_nand2_1
XFILLER_47_970 VPWR VGND sg13g2_decap_8
XFILLER_19_672 VPWR VGND sg13g2_decap_8
XFILLER_34_675 VPWR VGND sg13g2_decap_8
XFILLER_22_837 VPWR VGND sg13g2_decap_8
X_3626_ _1083_ net593 _1028_ VPWR VGND sg13g2_nand2_1
Xoutput19 net19 uio_out[2] VPWR VGND sg13g2_buf_1
X_3557_ _1022_ _0786_ _0867_ VPWR VGND sg13g2_xnor2_1
X_2508_ _1923_ net614 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[6\]
+ net618 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[6\] VPWR VGND
+ sg13g2_a22oi_1
X_3488_ VGND VPWR _0303_ _0875_ _0956_ _0955_ sg13g2_a21oi_1
X_2439_ _1807_ _1828_ _1830_ _1843_ _1856_ VPWR VGND sg13g2_and4_1
XFILLER_45_918 VPWR VGND sg13g2_decap_8
X_4109_ _1462_ VPWR _0183_ VGND net578 _1461_ sg13g2_o21ai_1
XFILLER_44_428 VPWR VGND sg13g2_decap_8
XFILLER_25_653 VPWR VGND sg13g2_decap_8
XFILLER_13_837 VPWR VGND sg13g2_decap_8
XFILLER_40_667 VPWR VGND sg13g2_decap_8
XFILLER_21_881 VPWR VGND sg13g2_decap_8
XFILLER_4_557 VPWR VGND sg13g2_decap_8
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_48_745 VPWR VGND sg13g2_decap_8
XFILLER_36_918 VPWR VGND sg13g2_decap_8
XFILLER_29_992 VPWR VGND sg13g2_decap_8
XFILLER_35_406 VPWR VGND sg13g2_fill_1
XFILLER_28_491 VPWR VGND sg13g2_decap_8
XFILLER_44_995 VPWR VGND sg13g2_decap_8
XFILLER_16_653 VPWR VGND sg13g2_decap_8
XFILLER_43_472 VPWR VGND sg13g2_decap_8
XFILLER_30_111 VPWR VGND sg13g2_fill_1
XFILLER_30_133 VPWR VGND sg13g2_fill_1
XFILLER_31_656 VPWR VGND sg13g2_decap_8
XFILLER_12_870 VPWR VGND sg13g2_decap_8
X_2790_ _0306_ net576 VPWR VGND _1867_ sg13g2_nand2b_2
XFILLER_8_885 VPWR VGND sg13g2_decap_8
X_3411_ _0743_ VPWR _0066_ VGND _0856_ _0880_ sg13g2_o21ai_1
X_3342_ _0808_ _0809_ _0810_ _0813_ VGND VPWR _0812_ sg13g2_nor4_2
Xfanout809 net813 net809 VPWR VGND sg13g2_buf_8
X_3273_ _0719_ _0731_ _0744_ VPWR VGND sg13g2_nor2_1
X_2224_ net770 net762 _1641_ VPWR VGND net767 sg13g2_nand3b_1
X_2155_ net766 net754 net755 _1572_ VPWR VGND sg13g2_nor3_1
XFILLER_39_767 VPWR VGND sg13g2_decap_8
X_2086_ VPWR _1504_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[2\]
+ VGND sg13g2_inv_1
XFILLER_26_439 VPWR VGND sg13g2_decap_8
XFILLER_22_634 VPWR VGND sg13g2_decap_8
XFILLER_35_995 VPWR VGND sg13g2_decap_8
XFILLER_10_807 VPWR VGND sg13g2_decap_8
X_2988_ _0487_ VPWR _0488_ VGND net781 _0334_ sg13g2_o21ai_1
XFILLER_21_188 VPWR VGND sg13g2_fill_1
X_3609_ VGND VPWR _1069_ _1068_ net32 sg13g2_or2_1
XFILLER_1_527 VPWR VGND sg13g2_decap_8
XFILLER_18_907 VPWR VGND sg13g2_decap_8
XFILLER_45_715 VPWR VGND sg13g2_decap_8
XFILLER_25_450 VPWR VGND sg13g2_decap_8
XFILLER_41_943 VPWR VGND sg13g2_decap_8
XFILLER_12_100 VPWR VGND sg13g2_fill_2
XFILLER_13_634 VPWR VGND sg13g2_decap_8
XFILLER_40_464 VPWR VGND sg13g2_decap_8
XFILLER_9_627 VPWR VGND sg13g2_decap_8
XFILLER_5_800 VPWR VGND sg13g2_decap_8
XFILLER_4_321 VPWR VGND sg13g2_fill_2
XFILLER_5_877 VPWR VGND sg13g2_decap_8
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_48_542 VPWR VGND sg13g2_decap_8
XFILLER_36_715 VPWR VGND sg13g2_decap_8
XFILLER_17_940 VPWR VGND sg13g2_decap_8
XFILLER_32_910 VPWR VGND sg13g2_decap_8
X_3960_ _1336_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[0\] sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[1\]
+ VPWR VGND sg13g2_nand2_2
XFILLER_44_792 VPWR VGND sg13g2_decap_8
X_2911_ _0380_ _0405_ _0413_ VPWR VGND sg13g2_and2_1
X_3891_ VGND VPWR _1541_ net653 _0144_ _1283_ sg13g2_a21oi_1
X_2842_ _2016_ _2018_ _2011_ _0346_ VPWR VGND sg13g2_nand3_1
XFILLER_32_987 VPWR VGND sg13g2_decap_8
X_2773_ _1587_ _0298_ _0002_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_682 VPWR VGND sg13g2_decap_8
Xfanout606 _0876_ net606 VPWR VGND sg13g2_buf_8
X_3325_ _0690_ _0748_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[4\]
+ _0796_ VPWR VGND sg13g2_nand3_1
Xfanout639 net640 net639 VPWR VGND sg13g2_buf_8
Xfanout628 net629 net628 VPWR VGND sg13g2_buf_8
Xfanout617 _1860_ net617 VPWR VGND sg13g2_buf_8
X_3256_ _0725_ _0726_ _0715_ _0727_ VPWR VGND sg13g2_nand3_1
X_2207_ _1624_ net770 net767 VPWR VGND sg13g2_nand2b_1
X_3187_ VPWR VGND net764 _0657_ _1886_ _1629_ _0658_ net734 sg13g2_a221oi_1
XFILLER_39_564 VPWR VGND sg13g2_decap_8
X_2138_ _1555_ net743 VPWR VGND sap_3_inst.controller_inst.stage\[1\] sg13g2_nand2b_2
X_2069_ _1487_ net748 VPWR VGND sg13g2_inv_2
XFILLER_23_921 VPWR VGND sg13g2_decap_8
XFILLER_35_792 VPWR VGND sg13g2_decap_8
XFILLER_10_604 VPWR VGND sg13g2_decap_8
XFILLER_23_998 VPWR VGND sg13g2_decap_8
XFILLER_2_869 VPWR VGND sg13g2_decap_8
XFILLER_49_328 VPWR VGND sg13g2_decap_8
XFILLER_45_512 VPWR VGND sg13g2_decap_8
XFILLER_40_1024 VPWR VGND sg13g2_decap_4
XFILLER_18_704 VPWR VGND sg13g2_decap_8
XFILLER_17_247 VPWR VGND sg13g2_fill_2
XFILLER_33_729 VPWR VGND sg13g2_decap_8
XFILLER_45_589 VPWR VGND sg13g2_decap_8
XFILLER_41_740 VPWR VGND sg13g2_decap_8
XFILLER_14_954 VPWR VGND sg13g2_decap_8
XFILLER_9_446 VPWR VGND sg13g2_fill_2
XFILLER_5_674 VPWR VGND sg13g2_decap_8
XFILLER_4_33 VPWR VGND sg13g2_fill_2
X_3110_ _0598_ net772 _1529_ VPWR VGND sg13g2_nand2_1
XFILLER_4_88 VPWR VGND sg13g2_decap_8
XFILLER_1_891 VPWR VGND sg13g2_decap_8
X_4090_ _1448_ VPWR _0178_ VGND net579 _1447_ sg13g2_o21ai_1
XFILLER_49_895 VPWR VGND sg13g2_decap_8
X_3041_ _0537_ _0538_ net704 _0539_ VPWR VGND sg13g2_nand3_1
XFILLER_36_512 VPWR VGND sg13g2_decap_8
XFILLER_36_589 VPWR VGND sg13g2_decap_8
X_3943_ _1314_ VPWR _1323_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[2\]
+ _1322_ sg13g2_o21ai_1
XFILLER_20_924 VPWR VGND sg13g2_decap_8
XFILLER_32_784 VPWR VGND sg13g2_decap_8
X_3874_ net659 _1273_ _1274_ VPWR VGND sg13g2_nor2_1
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
X_2825_ net723 _1761_ net742 _0329_ VPWR VGND sg13g2_nand3_1
X_2756_ _1620_ _1876_ _0279_ _0282_ _0283_ VPWR VGND sg13g2_and4_1
XFILLER_9_991 VPWR VGND sg13g2_decap_8
X_2687_ net3 _1884_ _0219_ VPWR VGND sg13g2_and2_1
X_4288_ net814 VGND VPWR _0145_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[7\]
+ clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3308_ _0779_ _0772_ _0773_ _0778_ VPWR VGND sg13g2_and3_2
X_3239_ VPWR VGND _0663_ _0650_ _0662_ net740 _0710_ _0647_ sg13g2_a221oi_1
XFILLER_15_707 VPWR VGND sg13g2_decap_8
XFILLER_27_567 VPWR VGND sg13g2_decap_8
XFILLER_42_548 VPWR VGND sg13g2_decap_8
Xfanout32 net20 net32 VPWR VGND sg13g2_buf_2
XFILLER_11_957 VPWR VGND sg13g2_decap_8
XFILLER_23_795 VPWR VGND sg13g2_decap_8
XFILLER_10_478 VPWR VGND sg13g2_decap_8
Xclkbuf_4_2_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_2_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_2_666 VPWR VGND sg13g2_decap_8
XFILLER_18_501 VPWR VGND sg13g2_decap_8
XFILLER_46_832 VPWR VGND sg13g2_decap_8
XFILLER_18_578 VPWR VGND sg13g2_decap_8
XFILLER_45_386 VPWR VGND sg13g2_decap_8
XFILLER_33_526 VPWR VGND sg13g2_decap_8
XFILLER_14_751 VPWR VGND sg13g2_decap_8
X_3590_ net641 _0875_ _1053_ VPWR VGND sg13g2_nor2_1
Xclkload13 VPWR clkload13/Y clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs VGND sg13g2_inv_1
X_2610_ _2019_ _2016_ _2018_ VPWR VGND sg13g2_nand2_1
X_2541_ _1768_ _1953_ _1954_ VPWR VGND sg13g2_nor2_1
XFILLER_47_1019 VPWR VGND sg13g2_decap_8
XFILLER_5_471 VPWR VGND sg13g2_decap_8
X_2472_ net734 VPWR _1889_ VGND _1629_ _1684_ sg13g2_o21ai_1
X_4211_ net813 VGND VPWR _0068_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[2\]
+ clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4142_ VGND VPWR _1467_ _0186_ _0194_ _1485_ sg13g2_a21oi_1
X_4073_ VGND VPWR net650 _1081_ _0174_ _1435_ sg13g2_a21oi_1
XFILLER_37_810 VPWR VGND sg13g2_decap_8
XFILLER_49_692 VPWR VGND sg13g2_decap_8
X_3024_ _0515_ VPWR _0523_ VGND _0479_ _0481_ sg13g2_o21ai_1
XFILLER_37_887 VPWR VGND sg13g2_decap_8
X_3926_ _1139_ _1307_ _1309_ _1310_ _1311_ VPWR VGND sg13g2_nor4_1
XFILLER_20_721 VPWR VGND sg13g2_decap_8
XFILLER_32_581 VPWR VGND sg13g2_decap_8
Xclkload7 clknet_1_1__leaf_clk_div_out clkload7/X VPWR VGND sg13g2_buf_1
XFILLER_30_1001 VPWR VGND sg13g2_decap_8
X_3857_ net572 net574 _1260_ VPWR VGND sg13g2_and2_1
X_2808_ net60 sap_3_inst.out\[1\] net799 _0018_ VPWR VGND sg13g2_mux2_1
XFILLER_20_798 VPWR VGND sg13g2_decap_8
X_3788_ _1216_ _1070_ _1071_ VPWR VGND sg13g2_nand2b_1
X_2739_ _0268_ _0266_ _0267_ VPWR VGND sg13g2_nand2_1
Xclkbuf_5_24__f_sap_3_inst.alu_inst.clk_regs clknet_4_12_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_28_876 VPWR VGND sg13g2_decap_8
XFILLER_15_504 VPWR VGND sg13g2_decap_8
XFILLER_43_857 VPWR VGND sg13g2_decap_8
XFILLER_23_592 VPWR VGND sg13g2_decap_8
XFILLER_11_754 VPWR VGND sg13g2_decap_8
XFILLER_7_758 VPWR VGND sg13g2_decap_8
XFILLER_3_931 VPWR VGND sg13g2_decap_8
XFILLER_2_463 VPWR VGND sg13g2_decap_8
Xclkbuf_5_13__f_sap_3_inst.alu_inst.clk_regs clknet_4_6_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_38_629 VPWR VGND sg13g2_decap_8
XFILLER_19_854 VPWR VGND sg13g2_decap_8
XFILLER_34_857 VPWR VGND sg13g2_decap_8
X_3711_ net582 _1155_ _1156_ VPWR VGND sg13g2_nor2_1
X_3642_ _1097_ net604 VPWR VGND sg13g2_inv_2
X_3573_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[7\] _1036_
+ net648 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[7\] _1037_ net671
+ sg13g2_a221oi_1
XFILLER_46_0 VPWR VGND sg13g2_decap_4
X_2524_ _1937_ _1938_ _1936_ _1939_ VPWR VGND sg13g2_nand3_1
X_2455_ VGND VPWR net764 _1686_ _1872_ _1633_ sg13g2_a21oi_1
X_2386_ _1803_ _1801_ _1697_ VPWR VGND sg13g2_nand2b_1
Xhold19 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[1\] VPWR VGND net66
+ sg13g2_dlygate4sd3_1
X_4125_ u_ser.shadow_reg\[0\] VPWR _1476_ VGND u_ser.state\[0\] _1489_ sg13g2_o21ai_1
XFILLER_29_607 VPWR VGND sg13g2_decap_8
X_4056_ _1425_ _1349_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[7\]
+ _1347_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3007_ net778 sap_3_inst.alu_inst.tmp\[5\] _0506_ VPWR VGND sg13g2_nor2_1
XFILLER_25_835 VPWR VGND sg13g2_decap_8
XFILLER_37_684 VPWR VGND sg13g2_decap_8
XFILLER_40_849 VPWR VGND sg13g2_decap_8
XFILLER_33_890 VPWR VGND sg13g2_decap_8
X_3909_ _1295_ _1296_ _0149_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_595 VPWR VGND sg13g2_decap_8
XFILLER_4_739 VPWR VGND sg13g2_decap_8
XFILLER_10_65 VPWR VGND sg13g2_fill_1
XFILLER_0_945 VPWR VGND sg13g2_decap_8
XFILLER_48_927 VPWR VGND sg13g2_decap_8
XFILLER_47_459 VPWR VGND sg13g2_decap_8
XFILLER_16_835 VPWR VGND sg13g2_decap_8
XFILLER_28_673 VPWR VGND sg13g2_decap_8
XFILLER_43_654 VPWR VGND sg13g2_decap_8
XFILLER_31_838 VPWR VGND sg13g2_decap_8
XFILLER_11_551 VPWR VGND sg13g2_decap_8
XFILLER_7_555 VPWR VGND sg13g2_decap_8
X_2240_ _1562_ _1573_ _1657_ VPWR VGND sg13g2_nor2_2
XFILLER_39_949 VPWR VGND sg13g2_decap_8
X_2171_ VPWR VGND net743 net718 net737 net741 _1588_ net727 sg13g2_a221oi_1
XFILLER_19_651 VPWR VGND sg13g2_decap_8
XFILLER_20_1022 VPWR VGND sg13g2_decap_8
XFILLER_18_172 VPWR VGND sg13g2_fill_1
XFILLER_22_816 VPWR VGND sg13g2_decap_8
XFILLER_34_654 VPWR VGND sg13g2_decap_8
XFILLER_30_882 VPWR VGND sg13g2_decap_8
X_3625_ VGND VPWR _1054_ _1081_ _0079_ _1082_ sg13g2_a21oi_1
XFILLER_1_709 VPWR VGND sg13g2_decap_8
X_3556_ _1017_ _1005_ _1020_ _1021_ VPWR VGND sg13g2_a21o_2
X_2507_ net697 net626 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[6\]
+ _1922_ VPWR VGND sg13g2_nand3_1
X_3487_ net32 _0875_ _0955_ VPWR VGND sg13g2_nor2_1
X_2438_ _1851_ _1854_ _1848_ _1855_ VPWR VGND sg13g2_nand3_1
X_2369_ VGND VPWR net725 _1630_ _1786_ _1609_ sg13g2_a21oi_1
X_4108_ _1462_ sap_3_inst.alu_inst.act\[6\] net578 VPWR VGND sg13g2_nand2_1
XFILLER_44_407 VPWR VGND sg13g2_decap_8
X_4039_ _0154_ VPWR _1410_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[5\]
+ _1344_ sg13g2_o21ai_1
XFILLER_38_993 VPWR VGND sg13g2_decap_8
XFILLER_25_632 VPWR VGND sg13g2_decap_8
XFILLER_13_816 VPWR VGND sg13g2_decap_8
XFILLER_9_809 VPWR VGND sg13g2_decap_8
XFILLER_40_646 VPWR VGND sg13g2_decap_8
XFILLER_8_319 VPWR VGND sg13g2_fill_1
XFILLER_21_860 VPWR VGND sg13g2_decap_8
XFILLER_4_536 VPWR VGND sg13g2_decap_8
XFILLER_43_1011 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_48_724 VPWR VGND sg13g2_decap_8
XFILLER_47_267 VPWR VGND sg13g2_fill_2
Xclkbuf_4_10_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs
+ clknet_4_10_0_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_29_971 VPWR VGND sg13g2_decap_8
XFILLER_16_632 VPWR VGND sg13g2_decap_8
XFILLER_28_470 VPWR VGND sg13g2_decap_8
XFILLER_44_974 VPWR VGND sg13g2_decap_8
XFILLER_43_451 VPWR VGND sg13g2_decap_8
XFILLER_31_635 VPWR VGND sg13g2_decap_8
XFILLER_8_864 VPWR VGND sg13g2_decap_8
XFILLER_7_55 VPWR VGND sg13g2_fill_2
XFILLER_7_66 VPWR VGND sg13g2_fill_2
X_3410_ _0881_ _0720_ _0731_ VPWR VGND sg13g2_nand2_2
X_3341_ net642 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[3\] _0811_
+ _0812_ VPWR VGND sg13g2_a21o_1
X_3272_ _0743_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[0\] net596
+ VPWR VGND sg13g2_nand2_1
X_2223_ net763 _1575_ _1616_ net749 _1640_ VPWR VGND sg13g2_or4_1
X_2154_ VGND VPWR _1571_ net755 net753 sg13g2_or2_1
XFILLER_39_746 VPWR VGND sg13g2_decap_8
XFILLER_38_278 VPWR VGND sg13g2_fill_2
X_2085_ VPWR _1503_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[2\]
+ VGND sg13g2_inv_1
XFILLER_35_974 VPWR VGND sg13g2_decap_8
XFILLER_22_613 VPWR VGND sg13g2_decap_8
X_2987_ _0487_ net691 net778 net692 net783 VPWR VGND sg13g2_a22oi_1
X_3608_ net613 _0952_ _1068_ VPWR VGND sg13g2_nor2_1
XFILLER_1_506 VPWR VGND sg13g2_decap_8
X_3539_ net590 net571 net573 _0990_ _1005_ VPWR VGND sg13g2_or4_1
XFILLER_38_790 VPWR VGND sg13g2_decap_8
XFILLER_26_985 VPWR VGND sg13g2_decap_8
XFILLER_41_922 VPWR VGND sg13g2_decap_8
XFILLER_13_613 VPWR VGND sg13g2_decap_8
XFILLER_9_606 VPWR VGND sg13g2_decap_8
XFILLER_41_999 VPWR VGND sg13g2_decap_8
XFILLER_5_856 VPWR VGND sg13g2_decap_8
XFILLER_10_1010 VPWR VGND sg13g2_decap_8
XFILLER_4_388 VPWR VGND sg13g2_fill_1
XFILLER_48_521 VPWR VGND sg13g2_decap_8
XFILLER_48_598 VPWR VGND sg13g2_decap_8
XFILLER_44_771 VPWR VGND sg13g2_decap_8
X_2910_ _0411_ _0405_ _0412_ VPWR VGND sg13g2_xor2_1
XFILLER_17_996 VPWR VGND sg13g2_decap_8
X_3890_ net653 _1139_ _1162_ _1283_ VPWR VGND sg13g2_nor3_1
XFILLER_32_966 VPWR VGND sg13g2_decap_8
X_2841_ _0345_ _2011_ _0333_ VPWR VGND sg13g2_nand2_1
X_2772_ _1491_ _0298_ _0001_ VPWR VGND sg13g2_and2_1
XFILLER_8_661 VPWR VGND sg13g2_decap_8
X_3324_ _0795_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[4\] net672
+ VPWR VGND sg13g2_nand2_1
Xfanout607 net608 net607 VPWR VGND sg13g2_buf_8
Xfanout629 _1847_ net629 VPWR VGND sg13g2_buf_8
Xfanout618 net619 net618 VPWR VGND sg13g2_buf_8
X_3255_ _1753_ VPWR _0726_ VGND _1651_ _0692_ sg13g2_o21ai_1
X_2206_ net767 net770 _1623_ VPWR VGND sg13g2_nor2b_2
XFILLER_39_543 VPWR VGND sg13g2_decap_8
X_3186_ net750 net727 _1837_ _0657_ VPWR VGND sg13g2_nor3_1
X_2137_ VGND VPWR _1554_ net746 net747 sg13g2_or2_1
XFILLER_27_749 VPWR VGND sg13g2_decap_8
XFILLER_23_900 VPWR VGND sg13g2_decap_8
XFILLER_35_771 VPWR VGND sg13g2_decap_8
XFILLER_23_977 VPWR VGND sg13g2_decap_8
XFILLER_22_487 VPWR VGND sg13g2_decap_8
XFILLER_2_848 VPWR VGND sg13g2_decap_8
XFILLER_49_307 VPWR VGND sg13g2_decap_8
XFILLER_40_1003 VPWR VGND sg13g2_decap_8
XFILLER_45_568 VPWR VGND sg13g2_decap_8
XFILLER_33_708 VPWR VGND sg13g2_decap_8
XFILLER_14_933 VPWR VGND sg13g2_decap_8
XFILLER_26_782 VPWR VGND sg13g2_decap_8
XFILLER_25_292 VPWR VGND sg13g2_decap_4
XFILLER_41_796 VPWR VGND sg13g2_decap_8
XFILLER_13_487 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_sap_3_inst.alu_inst.clk clknet_0_sap_3_inst.alu_inst.clk clknet_1_1__leaf_sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_5_653 VPWR VGND sg13g2_decap_8
XFILLER_4_141 VPWR VGND sg13g2_fill_2
XFILLER_4_67 VPWR VGND sg13g2_fill_2
XFILLER_1_870 VPWR VGND sg13g2_decap_8
XFILLER_49_874 VPWR VGND sg13g2_decap_8
X_3040_ _0535_ _0536_ _0502_ _0538_ VPWR VGND sg13g2_nand3_1
XFILLER_48_395 VPWR VGND sg13g2_decap_8
XFILLER_36_568 VPWR VGND sg13g2_decap_8
XFILLER_17_793 VPWR VGND sg13g2_decap_8
X_3942_ _1322_ _1315_ _1316_ VPWR VGND sg13g2_nand2_1
XFILLER_20_903 VPWR VGND sg13g2_decap_8
XFILLER_32_763 VPWR VGND sg13g2_decap_8
X_3873_ _1273_ _1018_ _1040_ VPWR VGND sg13g2_xnor2_1
X_2824_ net740 _1762_ _0328_ VPWR VGND sg13g2_nor2_1
XFILLER_9_970 VPWR VGND sg13g2_decap_8
X_2755_ _0282_ _1639_ _1692_ VPWR VGND sg13g2_nand2_1
X_2686_ VGND VPWR _1500_ _1900_ _0218_ _0217_ sg13g2_a21oi_1
X_3307_ _0774_ _0775_ _0776_ _0777_ _0778_ VPWR VGND sg13g2_and4_1
X_4287_ net811 VGND VPWR _0144_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[6\]
+ clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3238_ _0689_ _0708_ _0688_ _0709_ VPWR VGND sg13g2_nand3_1
X_3169_ _1889_ _0638_ _1816_ _0640_ VPWR VGND _0639_ sg13g2_nand4_1
XFILLER_27_546 VPWR VGND sg13g2_decap_8
XFILLER_42_527 VPWR VGND sg13g2_decap_8
XFILLER_23_774 VPWR VGND sg13g2_decap_8
XFILLER_11_936 VPWR VGND sg13g2_decap_8
XFILLER_2_645 VPWR VGND sg13g2_decap_8
XFILLER_1_122 VPWR VGND sg13g2_fill_2
XFILLER_46_811 VPWR VGND sg13g2_decap_8
XFILLER_18_557 VPWR VGND sg13g2_decap_8
XFILLER_46_888 VPWR VGND sg13g2_decap_8
XFILLER_45_365 VPWR VGND sg13g2_decap_8
XFILLER_33_505 VPWR VGND sg13g2_decap_8
XFILLER_14_730 VPWR VGND sg13g2_decap_8
XFILLER_41_593 VPWR VGND sg13g2_decap_8
Xclkload14 clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs clkload14/X VPWR VGND sg13g2_buf_1
X_2540_ _1943_ VPWR _1953_ VGND _1949_ _1952_ sg13g2_o21ai_1
XFILLER_5_450 VPWR VGND sg13g2_decap_8
X_2471_ _1612_ _1635_ _1557_ _1888_ VPWR VGND sg13g2_nand3_1
XFILLER_6_995 VPWR VGND sg13g2_decap_8
X_4210_ net805 VGND VPWR _0067_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_1
X_4141_ VGND VPWR net800 _0186_ _1485_ net71 sg13g2_a21oi_1
X_4072_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[5\] net650 _1435_
+ VPWR VGND sg13g2_nor2_1
XFILLER_49_671 VPWR VGND sg13g2_decap_8
X_3023_ _0475_ _0481_ _0508_ _0522_ VPWR VGND sg13g2_nor3_2
XFILLER_37_866 VPWR VGND sg13g2_decap_8
XFILLER_17_590 VPWR VGND sg13g2_decap_8
XFILLER_24_549 VPWR VGND sg13g2_decap_8
X_3925_ net647 VPWR _1310_ VGND net586 _1021_ sg13g2_o21ai_1
XFILLER_20_700 VPWR VGND sg13g2_decap_8
XFILLER_32_560 VPWR VGND sg13g2_decap_8
X_3856_ net652 _1119_ _1259_ VPWR VGND sg13g2_nor2_1
Xclkload8 clknet_1_1__leaf_sap_3_inst.alu_inst.clk clkload8/X VPWR VGND sg13g2_buf_8
XFILLER_20_777 VPWR VGND sg13g2_decap_8
X_2807_ net58 sap_3_inst.out\[0\] net799 _0017_ VPWR VGND sg13g2_mux2_1
X_3787_ VPWR _0108_ _1215_ VGND sg13g2_inv_1
X_2738_ sap_3_inst.alu_inst.act\[1\] sap_3_inst.alu_inst.act\[0\] sap_3_inst.alu_inst.act\[3\]
+ sap_3_inst.alu_inst.act\[2\] _0267_ VPWR VGND sg13g2_nor4_1
X_2669_ _0201_ _0202_ _0200_ _0203_ VPWR VGND sg13g2_nand3_1
XFILLER_8_1025 VPWR VGND sg13g2_decap_4
XFILLER_28_855 VPWR VGND sg13g2_decap_8
XFILLER_43_836 VPWR VGND sg13g2_decap_8
XFILLER_11_733 VPWR VGND sg13g2_decap_8
XFILLER_23_571 VPWR VGND sg13g2_decap_8
XFILLER_24_53 VPWR VGND sg13g2_fill_2
XFILLER_10_243 VPWR VGND sg13g2_fill_2
XFILLER_24_86 VPWR VGND sg13g2_fill_1
XFILLER_7_737 VPWR VGND sg13g2_decap_8
XFILLER_3_910 VPWR VGND sg13g2_decap_8
XFILLER_3_987 VPWR VGND sg13g2_decap_8
XFILLER_38_608 VPWR VGND sg13g2_decap_8
Xfanout790 net791 net790 VPWR VGND sg13g2_buf_1
XFILLER_19_833 VPWR VGND sg13g2_decap_8
XFILLER_46_685 VPWR VGND sg13g2_decap_8
XFILLER_34_836 VPWR VGND sg13g2_decap_8
XFILLER_42_891 VPWR VGND sg13g2_decap_8
X_3710_ net611 _0931_ _1155_ VPWR VGND sg13g2_and2_1
X_3641_ net636 net668 _1096_ VPWR VGND sg13g2_nor2_1
X_3572_ _1034_ _1035_ net660 _1036_ VPWR VGND sg13g2_nand3_1
X_2523_ _1938_ net616 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[6\]
+ net618 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[6\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_6_792 VPWR VGND sg13g2_decap_8
X_2454_ _1627_ _1648_ _1654_ _1699_ _1871_ VPWR VGND sg13g2_nor4_1
X_2385_ VGND VPWR _1640_ _1647_ _1802_ _1631_ sg13g2_a21oi_1
XFILLER_39_0 VPWR VGND sg13g2_fill_2
X_4124_ _1465_ _1474_ _1490_ _1475_ VPWR VGND sg13g2_nand3_1
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
X_4055_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[7\] _1351_
+ _1424_ net794 sg13g2_a21oi_1
X_3006_ VGND VPWR _0501_ _0503_ _0505_ _0504_ sg13g2_a21oi_1
XFILLER_25_814 VPWR VGND sg13g2_decap_8
XFILLER_37_663 VPWR VGND sg13g2_decap_8
XFILLER_40_828 VPWR VGND sg13g2_decap_8
XFILLER_24_379 VPWR VGND sg13g2_fill_1
X_3908_ net649 _1182_ _0303_ _1296_ VPWR VGND _1183_ sg13g2_nand4_1
XFILLER_20_574 VPWR VGND sg13g2_decap_8
X_3839_ _0865_ net585 _1246_ VPWR VGND sg13g2_nor2_1
XFILLER_4_718 VPWR VGND sg13g2_decap_8
XFILLER_0_924 VPWR VGND sg13g2_decap_8
XFILLER_48_906 VPWR VGND sg13g2_decap_8
XFILLER_47_438 VPWR VGND sg13g2_decap_8
XFILLER_19_42 VPWR VGND sg13g2_fill_1
XFILLER_28_652 VPWR VGND sg13g2_decap_8
XFILLER_16_814 VPWR VGND sg13g2_decap_8
XFILLER_43_633 VPWR VGND sg13g2_decap_8
XFILLER_15_368 VPWR VGND sg13g2_fill_2
XFILLER_31_817 VPWR VGND sg13g2_decap_8
XFILLER_30_327 VPWR VGND sg13g2_fill_1
XFILLER_11_530 VPWR VGND sg13g2_decap_8
XFILLER_30_338 VPWR VGND sg13g2_fill_2
XFILLER_7_534 VPWR VGND sg13g2_decap_8
XFILLER_3_784 VPWR VGND sg13g2_decap_8
XFILLER_39_928 VPWR VGND sg13g2_decap_8
X_2170_ _1587_ net747 net746 VPWR VGND sg13g2_xnor2_1
XFILLER_19_630 VPWR VGND sg13g2_decap_8
XFILLER_20_1001 VPWR VGND sg13g2_decap_8
XFILLER_46_482 VPWR VGND sg13g2_decap_8
XFILLER_34_633 VPWR VGND sg13g2_decap_8
XFILLER_14_390 VPWR VGND sg13g2_fill_2
XFILLER_30_861 VPWR VGND sg13g2_decap_8
X_3624_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[5\] _1054_ _1082_
+ VPWR VGND sg13g2_nor2_1
X_3555_ net590 net571 net573 _1019_ _1020_ VPWR VGND sg13g2_nor4_1
X_2506_ _1921_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[6\] net628
+ VPWR VGND sg13g2_nand2_1
X_3486_ VGND VPWR net665 _0951_ _0954_ _0953_ sg13g2_a21oi_1
X_2437_ _1854_ net623 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[7\]
+ net624 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_1017 VPWR VGND sg13g2_decap_8
X_2368_ _1785_ net730 _1602_ _1775_ VPWR VGND sg13g2_and3_1
X_2299_ _1665_ VPWR _1716_ VGND _1678_ _1715_ sg13g2_o21ai_1
X_4107_ _1460_ VPWR _1461_ VGND _0547_ _1439_ sg13g2_o21ai_1
XFILLER_38_972 VPWR VGND sg13g2_decap_8
X_4038_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[5\] _1408_
+ _1352_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[5\] _1409_ _1347_
+ sg13g2_a221oi_1
XFILLER_25_611 VPWR VGND sg13g2_decap_8
XFILLER_24_143 VPWR VGND sg13g2_fill_2
XFILLER_40_625 VPWR VGND sg13g2_decap_8
XFILLER_25_688 VPWR VGND sg13g2_decap_8
XFILLER_4_515 VPWR VGND sg13g2_decap_8
XFILLER_0_721 VPWR VGND sg13g2_decap_8
XFILLER_48_703 VPWR VGND sg13g2_decap_8
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_29_950 VPWR VGND sg13g2_decap_8
XFILLER_16_611 VPWR VGND sg13g2_decap_8
XFILLER_44_953 VPWR VGND sg13g2_decap_8
XFILLER_16_688 VPWR VGND sg13g2_decap_8
XFILLER_31_614 VPWR VGND sg13g2_decap_8
XFILLER_8_843 VPWR VGND sg13g2_decap_8
XFILLER_7_89 VPWR VGND sg13g2_decap_8
X_3340_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[3\] _0763_ _0811_
+ VPWR VGND sg13g2_and2_1
XFILLER_3_581 VPWR VGND sg13g2_decap_8
X_3271_ _0742_ net596 VPWR VGND sg13g2_inv_2
X_2222_ net762 _1575_ _1616_ _1639_ VGND VPWR _1625_ sg13g2_nor4_2
XFILLER_39_725 VPWR VGND sg13g2_decap_8
X_2153_ net753 net755 _1570_ VPWR VGND sg13g2_nor2_1
XFILLER_26_419 VPWR VGND sg13g2_fill_2
X_2084_ VPWR _1502_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[2\]
+ VGND sg13g2_inv_1
XFILLER_35_953 VPWR VGND sg13g2_decap_8
XFILLER_22_669 VPWR VGND sg13g2_decap_8
X_2986_ _0485_ VPWR _0486_ VGND _0346_ _0480_ sg13g2_o21ai_1
X_3607_ _0076_ _1065_ _1067_ net583 _1507_ VPWR VGND sg13g2_a22oi_1
X_3538_ net571 net574 _0990_ _1004_ VPWR VGND sg13g2_nor3_1
X_3469_ _0937_ net639 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[3\]
+ net642 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_41_901 VPWR VGND sg13g2_decap_8
XFILLER_26_964 VPWR VGND sg13g2_decap_8
XFILLER_12_102 VPWR VGND sg13g2_fill_1
XFILLER_25_485 VPWR VGND sg13g2_decap_8
XFILLER_41_978 VPWR VGND sg13g2_decap_8
XFILLER_13_669 VPWR VGND sg13g2_decap_8
XFILLER_40_499 VPWR VGND sg13g2_decap_8
XFILLER_32_86 VPWR VGND sg13g2_fill_2
XFILLER_5_835 VPWR VGND sg13g2_decap_8
XFILLER_4_323 VPWR VGND sg13g2_fill_1
XFILLER_48_500 VPWR VGND sg13g2_decap_8
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_48_577 VPWR VGND sg13g2_decap_8
XFILLER_44_750 VPWR VGND sg13g2_decap_8
XFILLER_17_975 VPWR VGND sg13g2_decap_8
XFILLER_16_485 VPWR VGND sg13g2_decap_8
X_2840_ _2011_ _0333_ _0344_ VPWR VGND sg13g2_and2_1
XFILLER_32_945 VPWR VGND sg13g2_decap_8
XFILLER_8_640 VPWR VGND sg13g2_decap_8
X_2771_ _1581_ net743 _0297_ _0298_ VPWR VGND sg13g2_a21o_1
Xclkbuf_4_3_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_3_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
Xfanout608 net611 net608 VPWR VGND sg13g2_buf_2
Xfanout619 _1859_ net619 VPWR VGND sg13g2_buf_8
X_3323_ _0791_ _0792_ _0789_ _0794_ VPWR VGND sg13g2_nand3_1
X_3254_ _0668_ _0722_ _0723_ _0724_ _0725_ VPWR VGND sg13g2_nor4_1
X_2205_ _1621_ _1615_ _1602_ _1622_ VPWR VGND sg13g2_a21o_1
XFILLER_39_522 VPWR VGND sg13g2_decap_8
XFILLER_2_1009 VPWR VGND sg13g2_decap_8
X_3185_ _0656_ _1731_ _1782_ VPWR VGND sg13g2_nand2_1
X_2136_ net747 net746 _1553_ VPWR VGND sg13g2_nor2_2
XFILLER_27_728 VPWR VGND sg13g2_decap_8
XFILLER_39_599 VPWR VGND sg13g2_decap_8
XFILLER_42_709 VPWR VGND sg13g2_decap_8
XFILLER_35_750 VPWR VGND sg13g2_decap_8
XFILLER_41_219 VPWR VGND sg13g2_fill_1
XFILLER_23_956 VPWR VGND sg13g2_decap_8
XFILLER_22_466 VPWR VGND sg13g2_decap_8
X_2969_ _0453_ VPWR _0469_ VGND net783 net708 sg13g2_o21ai_1
XFILLER_10_639 VPWR VGND sg13g2_decap_8
XFILLER_2_827 VPWR VGND sg13g2_decap_8
XFILLER_18_739 VPWR VGND sg13g2_decap_8
XFILLER_45_547 VPWR VGND sg13g2_decap_8
XFILLER_14_912 VPWR VGND sg13g2_decap_8
XFILLER_26_761 VPWR VGND sg13g2_decap_8
XFILLER_41_775 VPWR VGND sg13g2_decap_8
XFILLER_40_230 VPWR VGND sg13g2_fill_2
XFILLER_14_989 VPWR VGND sg13g2_decap_8
XFILLER_40_274 VPWR VGND sg13g2_fill_2
XFILLER_9_437 VPWR VGND sg13g2_fill_2
XFILLER_9_448 VPWR VGND sg13g2_fill_1
XFILLER_5_632 VPWR VGND sg13g2_decap_8
XFILLER_4_197 VPWR VGND sg13g2_fill_2
XFILLER_4_46 VPWR VGND sg13g2_fill_2
XFILLER_4_35 VPWR VGND sg13g2_fill_1
XFILLER_4_79 VPWR VGND sg13g2_decap_4
XFILLER_49_853 VPWR VGND sg13g2_decap_8
XFILLER_48_374 VPWR VGND sg13g2_decap_8
XFILLER_36_547 VPWR VGND sg13g2_decap_8
XFILLER_17_772 VPWR VGND sg13g2_decap_8
XFILLER_32_742 VPWR VGND sg13g2_decap_8
X_3941_ _1321_ net61 _1314_ VPWR VGND sg13g2_nand2_1
X_3872_ _1272_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[7\] net652
+ VPWR VGND sg13g2_nand2_1
XFILLER_17_1017 VPWR VGND sg13g2_decap_8
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
XFILLER_31_252 VPWR VGND sg13g2_fill_2
X_2823_ VPWR VGND _0325_ _0326_ _0321_ _1592_ _0327_ net723 sg13g2_a221oi_1
XFILLER_20_959 VPWR VGND sg13g2_decap_8
X_2754_ VGND VPWR net705 _0280_ _0281_ _1651_ sg13g2_a21oi_1
X_2685_ VGND VPWR sap_3_inst.alu_flags\[2\] _1902_ _0217_ _1900_ sg13g2_a21oi_1
X_3306_ _0777_ net638 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[7\]
+ net671 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4286_ net830 VGND VPWR _0143_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[5\]
+ clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3237_ _0708_ _1869_ VPWR VGND _0706_ sg13g2_nand2b_2
X_3168_ _0639_ _1822_ _1875_ _1699_ _1633_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_525 VPWR VGND sg13g2_decap_8
X_2119_ VPWR _1537_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[5\]
+ VGND sg13g2_inv_1
XFILLER_42_506 VPWR VGND sg13g2_decap_8
X_3099_ net599 net773 _0595_ _0040_ VPWR VGND sg13g2_a21o_1
XFILLER_11_915 VPWR VGND sg13g2_decap_8
XFILLER_23_753 VPWR VGND sg13g2_decap_8
XFILLER_10_403 VPWR VGND sg13g2_fill_2
XFILLER_7_919 VPWR VGND sg13g2_decap_8
XFILLER_2_624 VPWR VGND sg13g2_decap_8
XFILLER_1_101 VPWR VGND sg13g2_fill_1
XFILLER_38_85 VPWR VGND sg13g2_fill_2
XFILLER_46_867 VPWR VGND sg13g2_decap_8
XFILLER_18_536 VPWR VGND sg13g2_decap_8
XFILLER_41_572 VPWR VGND sg13g2_decap_8
XFILLER_14_786 VPWR VGND sg13g2_decap_8
Xclkload15 VPWR clkload15/Y clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs VGND sg13g2_inv_1
XFILLER_6_974 VPWR VGND sg13g2_decap_8
X_2470_ VGND VPWR _1887_ _1876_ net764 sg13g2_or2_1
X_4140_ VGND VPWR net800 _0186_ _0193_ _1484_ sg13g2_a21oi_1
XFILLER_49_650 VPWR VGND sg13g2_decap_8
X_4071_ _0173_ _1075_ _1434_ net646 _1530_ VPWR VGND sg13g2_a22oi_1
X_3022_ _0519_ _0491_ _0521_ VPWR VGND sg13g2_xor2_1
XFILLER_37_845 VPWR VGND sg13g2_decap_8
XFILLER_24_528 VPWR VGND sg13g2_decap_8
X_3924_ VGND VPWR net570 net644 _1309_ _1308_ sg13g2_a21oi_1
XFILLER_20_756 VPWR VGND sg13g2_decap_8
Xclkload9 VPWR clkload9/Y clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs VGND sg13g2_inv_1
X_3855_ _0133_ _1183_ _1258_ net654 _1498_ VPWR VGND sg13g2_a22oi_1
X_2806_ u_ser.state\[0\] u_ser.state\[1\] _0185_ VPWR VGND sg13g2_nor2_2
X_3786_ _1215_ _1214_ _1154_ net580 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[2\]
+ VPWR VGND sg13g2_a22oi_1
X_2737_ sap_3_inst.alu_inst.act\[5\] sap_3_inst.alu_inst.act\[4\] sap_3_inst.alu_inst.act\[7\]
+ sap_3_inst.alu_inst.act\[6\] _0266_ VPWR VGND sg13g2_nor4_1
X_2668_ _0202_ net618 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[3\]
+ net632 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_8_1004 VPWR VGND sg13g2_decap_8
X_2599_ net731 _1618_ _2008_ VPWR VGND sg13g2_and2_1
X_4338_ net818 VGND VPWR net69 u_ser.bit_pos\[2\] clknet_3_0__leaf_clk sg13g2_dfrbpq_1
X_4269_ net815 VGND VPWR _0126_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[4\]
+ clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_28_834 VPWR VGND sg13g2_decap_8
XFILLER_43_815 VPWR VGND sg13g2_decap_8
XFILLER_42_303 VPWR VGND sg13g2_fill_1
XFILLER_15_539 VPWR VGND sg13g2_decap_8
XFILLER_23_550 VPWR VGND sg13g2_decap_8
XFILLER_11_712 VPWR VGND sg13g2_decap_8
XFILLER_7_716 VPWR VGND sg13g2_decap_8
XFILLER_11_789 VPWR VGND sg13g2_decap_8
XFILLER_46_1021 VPWR VGND sg13g2_decap_8
XFILLER_3_966 VPWR VGND sg13g2_decap_8
XFILLER_2_498 VPWR VGND sg13g2_decap_8
Xfanout791 sap_3_inst.alu_inst.acc\[1\] net791 VPWR VGND sg13g2_buf_8
Xfanout780 sap_3_inst.alu_inst.acc\[5\] net780 VPWR VGND sg13g2_buf_8
XFILLER_19_812 VPWR VGND sg13g2_decap_8
Xclkbuf_5_4__f_sap_3_inst.alu_inst.clk_regs clknet_4_2_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_46_664 VPWR VGND sg13g2_decap_8
XFILLER_19_889 VPWR VGND sg13g2_decap_8
XFILLER_33_303 VPWR VGND sg13g2_fill_2
XFILLER_34_815 VPWR VGND sg13g2_decap_8
XFILLER_42_870 VPWR VGND sg13g2_decap_8
XFILLER_14_583 VPWR VGND sg13g2_decap_8
X_3640_ VGND VPWR net595 _0855_ _1095_ _1056_ sg13g2_a21oi_1
X_3571_ _1035_ net680 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[7\]
+ net686 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2522_ _1937_ net622 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[6\]
+ net628 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_771 VPWR VGND sg13g2_decap_8
X_2453_ _1578_ VPWR _1870_ VGND net740 net722 sg13g2_o21ai_1
X_2384_ _1801_ _1800_ _1557_ _1686_ _1654_ VPWR VGND sg13g2_a22oi_1
X_4123_ u_ser.bit_pos\[0\] u_ser.shadow_reg\[1\] u_ser.shadow_reg\[2\] u_ser.shadow_reg\[3\]
+ u_ser.shadow_reg\[4\] u_ser.bit_pos\[1\] _1474_ VPWR VGND sg13g2_mux4_1
Xclkbuf_4_11_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs
+ clknet_4_11_0_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
X_4054_ _1423_ _1340_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[7\]
+ net797 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3005_ net704 VPWR _0504_ VGND _0501_ _0503_ sg13g2_o21ai_1
XFILLER_37_642 VPWR VGND sg13g2_decap_8
XFILLER_40_807 VPWR VGND sg13g2_decap_8
X_3907_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[3\] net650 _1295_
+ VPWR VGND sg13g2_nor2_1
XFILLER_20_553 VPWR VGND sg13g2_decap_8
X_3838_ _0771_ VPWR _1245_ VGND _0779_ _0864_ sg13g2_o21ai_1
X_3769_ _1140_ _1200_ _1201_ _1202_ VPWR VGND sg13g2_nor3_1
XFILLER_10_56 VPWR VGND sg13g2_fill_1
XFILLER_0_903 VPWR VGND sg13g2_decap_8
XFILLER_47_417 VPWR VGND sg13g2_decap_8
XFILLER_28_631 VPWR VGND sg13g2_decap_8
XFILLER_43_612 VPWR VGND sg13g2_decap_8
XFILLER_35_75 VPWR VGND sg13g2_fill_1
XFILLER_43_689 VPWR VGND sg13g2_decap_8
XFILLER_42_166 VPWR VGND sg13g2_fill_2
XFILLER_24_892 VPWR VGND sg13g2_decap_8
XFILLER_7_513 VPWR VGND sg13g2_decap_8
XFILLER_11_586 VPWR VGND sg13g2_decap_8
XFILLER_3_763 VPWR VGND sg13g2_decap_8
XFILLER_39_907 VPWR VGND sg13g2_decap_8
XFILLER_47_984 VPWR VGND sg13g2_decap_8
XFILLER_46_461 VPWR VGND sg13g2_decap_8
XFILLER_19_686 VPWR VGND sg13g2_decap_8
XFILLER_33_100 VPWR VGND sg13g2_fill_1
XFILLER_34_612 VPWR VGND sg13g2_decap_8
XFILLER_34_689 VPWR VGND sg13g2_decap_8
XFILLER_30_840 VPWR VGND sg13g2_decap_8
X_3623_ _1081_ _1079_ _1080_ VPWR VGND sg13g2_nand2_2
X_3554_ VGND VPWR _1019_ _1017_ _0990_ sg13g2_or2_1
X_2505_ _1920_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[6\] net711
+ VPWR VGND sg13g2_nand2_1
X_3485_ _0952_ _0713_ net613 _0953_ VPWR VGND sg13g2_a21o_1
X_2436_ net667 net666 net707 _1844_ _1853_ VPWR VGND sg13g2_and4_1
X_2367_ VGND VPWR _1672_ _1699_ _1784_ _1710_ sg13g2_a21oi_1
X_2298_ _1695_ _1713_ _1689_ _1715_ VPWR VGND _1714_ sg13g2_nand4_1
X_4106_ VGND VPWR _1460_ net699 net776 sg13g2_or2_1
XFILLER_38_951 VPWR VGND sg13g2_decap_8
X_4037_ _1405_ _1406_ _1403_ _1408_ VPWR VGND _1407_ sg13g2_nand4_1
XFILLER_25_667 VPWR VGND sg13g2_decap_8
XFILLER_40_604 VPWR VGND sg13g2_decap_8
XFILLER_21_895 VPWR VGND sg13g2_decap_8
XFILLER_0_700 VPWR VGND sg13g2_decap_8
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_48_759 VPWR VGND sg13g2_decap_8
XFILLER_46_63 VPWR VGND sg13g2_fill_1
XFILLER_44_932 VPWR VGND sg13g2_decap_8
XFILLER_15_122 VPWR VGND sg13g2_fill_1
XFILLER_16_667 VPWR VGND sg13g2_decap_8
XFILLER_43_486 VPWR VGND sg13g2_decap_8
XFILLER_8_822 VPWR VGND sg13g2_decap_8
XFILLER_12_884 VPWR VGND sg13g2_decap_8
XFILLER_8_899 VPWR VGND sg13g2_decap_8
XFILLER_7_343 VPWR VGND sg13g2_fill_2
XFILLER_7_68 VPWR VGND sg13g2_fill_1
XFILLER_3_560 VPWR VGND sg13g2_decap_8
X_3270_ net664 VPWR _0741_ VGND _0732_ _0740_ sg13g2_o21ai_1
X_2221_ net770 net749 _1638_ VPWR VGND sg13g2_nor2_1
XFILLER_39_704 VPWR VGND sg13g2_decap_8
X_2152_ _1569_ _1559_ _1564_ VPWR VGND sg13g2_nand2_2
X_2083_ _1501_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[2\] VPWR
+ VGND sg13g2_inv_2
XFILLER_47_781 VPWR VGND sg13g2_decap_8
XFILLER_19_483 VPWR VGND sg13g2_decap_8
XFILLER_35_932 VPWR VGND sg13g2_decap_8
XFILLER_22_648 VPWR VGND sg13g2_decap_8
X_2985_ _0485_ _0363_ _0473_ VPWR VGND sg13g2_nand2_1
XFILLER_21_169 VPWR VGND sg13g2_fill_1
X_3606_ net583 _1066_ _1067_ VPWR VGND sg13g2_nor2_1
X_3537_ _0997_ _0999_ _1002_ _1003_ VPWR VGND sg13g2_nor3_1
XFILLER_27_1008 VPWR VGND sg13g2_decap_8
X_3468_ _0936_ net650 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[3\]
+ net673 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2419_ net764 _1835_ _1836_ VPWR VGND sg13g2_nor2_1
X_3399_ _0870_ net608 _0869_ VPWR VGND sg13g2_nand2_2
XFILLER_45_729 VPWR VGND sg13g2_decap_8
XFILLER_26_943 VPWR VGND sg13g2_decap_8
XFILLER_25_464 VPWR VGND sg13g2_decap_8
XFILLER_41_957 VPWR VGND sg13g2_decap_8
XFILLER_13_648 VPWR VGND sg13g2_decap_8
XFILLER_40_478 VPWR VGND sg13g2_decap_8
XFILLER_21_692 VPWR VGND sg13g2_decap_8
XFILLER_5_814 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_48_556 VPWR VGND sg13g2_decap_8
XFILLER_36_729 VPWR VGND sg13g2_decap_8
XFILLER_17_954 VPWR VGND sg13g2_decap_8
XFILLER_32_924 VPWR VGND sg13g2_decap_8
XFILLER_12_681 VPWR VGND sg13g2_decap_8
X_2770_ _0296_ VPWR _0297_ VGND net751 _1569_ sg13g2_o21ai_1
XFILLER_8_696 VPWR VGND sg13g2_decap_8
XFILLER_7_195 VPWR VGND sg13g2_fill_2
Xfanout609 net610 net609 VPWR VGND sg13g2_buf_8
X_3322_ _0793_ _0789_ _0791_ _0792_ VPWR VGND sg13g2_and3_2
X_3253_ _1620_ VPWR _0724_ VGND _1613_ _1776_ sg13g2_o21ai_1
XFILLER_39_501 VPWR VGND sg13g2_decap_8
X_2204_ VPWR _1621_ _1620_ VGND sg13g2_inv_1
X_3184_ VGND VPWR _1658_ _0654_ _0655_ net721 sg13g2_a21oi_1
X_2135_ VGND VPWR _1552_ net744 net745 sg13g2_or2_1
XFILLER_27_707 VPWR VGND sg13g2_decap_8
XFILLER_39_578 VPWR VGND sg13g2_decap_8
XFILLER_23_935 VPWR VGND sg13g2_decap_8
XFILLER_34_283 VPWR VGND sg13g2_fill_2
XFILLER_10_618 VPWR VGND sg13g2_decap_8
XFILLER_22_445 VPWR VGND sg13g2_decap_8
X_2968_ _0468_ net781 net708 VPWR VGND sg13g2_xnor2_1
XFILLER_33_1023 VPWR VGND sg13g2_decap_4
X_2899_ VGND VPWR _2051_ net694 _0402_ net599 sg13g2_a21oi_1
XFILLER_2_806 VPWR VGND sg13g2_decap_8
XFILLER_18_718 VPWR VGND sg13g2_decap_8
XFILLER_45_526 VPWR VGND sg13g2_decap_8
XFILLER_26_740 VPWR VGND sg13g2_decap_8
XFILLER_41_754 VPWR VGND sg13g2_decap_8
XFILLER_14_968 VPWR VGND sg13g2_decap_8
XFILLER_5_611 VPWR VGND sg13g2_decap_8
XFILLER_5_688 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_fill_2
XFILLER_4_58 VPWR VGND sg13g2_decap_4
XFILLER_4_69 VPWR VGND sg13g2_fill_1
XFILLER_49_832 VPWR VGND sg13g2_decap_8
XFILLER_48_353 VPWR VGND sg13g2_decap_8
XFILLER_36_526 VPWR VGND sg13g2_decap_8
XFILLER_1_1010 VPWR VGND sg13g2_decap_8
XFILLER_17_751 VPWR VGND sg13g2_decap_8
X_3940_ VGND VPWR net803 _0155_ _1320_ net54 sg13g2_a21oi_1
XFILLER_32_721 VPWR VGND sg13g2_decap_8
X_3871_ _1271_ VPWR _0136_ VGND _1542_ net674 sg13g2_o21ai_1
X_2822_ _1565_ net728 _1762_ _0326_ VPWR VGND sg13g2_nor3_1
XFILLER_20_938 VPWR VGND sg13g2_decap_8
XFILLER_32_798 VPWR VGND sg13g2_decap_8
X_2753_ _1692_ VPWR _0280_ VGND _1627_ _1635_ sg13g2_o21ai_1
XFILLER_8_493 VPWR VGND sg13g2_decap_8
X_2684_ VPWR VGND _0215_ _1768_ _0211_ _1501_ _0216_ net633 sg13g2_a221oi_1
X_3305_ _0776_ net675 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[7\]
+ net665 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4285_ net815 VGND VPWR _0142_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[4\]
+ clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3236_ _1870_ _0706_ _0707_ VPWR VGND sg13g2_nor2_2
X_3167_ _1659_ VPWR _0638_ VGND _1633_ _1705_ sg13g2_o21ai_1
XFILLER_27_504 VPWR VGND sg13g2_decap_8
XFILLER_39_375 VPWR VGND sg13g2_fill_2
X_2118_ VPWR _1536_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[5\]
+ VGND sg13g2_inv_1
X_3098_ VPWR VGND _0594_ net599 _0593_ _1914_ _0595_ net694 sg13g2_a221oi_1
XFILLER_23_732 VPWR VGND sg13g2_decap_8
XFILLER_10_459 VPWR VGND sg13g2_fill_1
XFILLER_2_603 VPWR VGND sg13g2_decap_8
XFILLER_49_128 VPWR VGND sg13g2_fill_1
XFILLER_38_31 VPWR VGND sg13g2_fill_2
XFILLER_18_515 VPWR VGND sg13g2_decap_8
XFILLER_46_846 VPWR VGND sg13g2_decap_8
XFILLER_41_551 VPWR VGND sg13g2_decap_8
XFILLER_14_765 VPWR VGND sg13g2_decap_8
XFILLER_9_213 VPWR VGND sg13g2_fill_1
Xclkload16 VPWR clkload16/Y clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs VGND sg13g2_inv_1
XFILLER_10_982 VPWR VGND sg13g2_decap_8
XFILLER_6_953 VPWR VGND sg13g2_decap_8
XFILLER_5_485 VPWR VGND sg13g2_decap_8
X_4070_ net644 _1074_ _1434_ VPWR VGND sg13g2_nor2_1
X_3021_ _0491_ _0519_ _0520_ VPWR VGND sg13g2_nor2_1
XFILLER_37_824 VPWR VGND sg13g2_decap_8
XFILLER_24_507 VPWR VGND sg13g2_decap_8
XFILLER_45_890 VPWR VGND sg13g2_decap_8
X_3923_ net15 net644 _1308_ VPWR VGND sg13g2_nor2_1
X_3854_ VGND VPWR net572 _1256_ _1258_ _1257_ sg13g2_a21oi_1
X_2805_ VGND VPWR mem_mar_we _0318_ _1556_ sg13g2_or2_1
XFILLER_20_735 VPWR VGND sg13g2_decap_8
XFILLER_32_595 VPWR VGND sg13g2_decap_8
X_3785_ _1155_ net580 _1214_ VPWR VGND sg13g2_nor2_1
XFILLER_30_1015 VPWR VGND sg13g2_decap_8
X_2736_ _0263_ _0264_ _2056_ _0265_ VPWR VGND sg13g2_nand3_1
X_2667_ _0201_ net600 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[3\]
+ net629 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2598_ _1570_ _1893_ net765 _2007_ VPWR VGND sg13g2_nand3_1
X_4337_ net818 VGND VPWR _0194_ u_ser.bit_pos\[1\] clknet_3_1__leaf_clk sg13g2_dfrbpq_2
X_4268_ net831 VGND VPWR _0125_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[3\]
+ clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3219_ _0690_ _0688_ _0689_ VPWR VGND sg13g2_nand2_2
XFILLER_28_813 VPWR VGND sg13g2_decap_8
X_4199_ net824 VGND VPWR _0056_ sap_3_inst.alu_inst.tmp\[6\] clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_27_312 VPWR VGND sg13g2_fill_2
XFILLER_15_518 VPWR VGND sg13g2_decap_8
XFILLER_36_890 VPWR VGND sg13g2_decap_8
XFILLER_24_33 VPWR VGND sg13g2_fill_2
XFILLER_10_245 VPWR VGND sg13g2_fill_1
XFILLER_11_768 VPWR VGND sg13g2_decap_8
XFILLER_46_1000 VPWR VGND sg13g2_decap_8
XFILLER_3_945 VPWR VGND sg13g2_decap_8
XFILLER_2_477 VPWR VGND sg13g2_decap_8
Xfanout781 net782 net781 VPWR VGND sg13g2_buf_8
Xfanout792 net793 net792 VPWR VGND sg13g2_buf_8
Xfanout770 net771 net770 VPWR VGND sg13g2_buf_8
XFILLER_46_643 VPWR VGND sg13g2_decap_8
XFILLER_18_334 VPWR VGND sg13g2_fill_2
XFILLER_19_868 VPWR VGND sg13g2_decap_8
XFILLER_14_562 VPWR VGND sg13g2_decap_8
X_3570_ _1034_ net675 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[7\]
+ net683 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[7\] VPWR VGND sg13g2_a22oi_1
X_2521_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[6\] net621
+ net601 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[6\] _1936_ net711
+ sg13g2_a221oi_1
XFILLER_6_750 VPWR VGND sg13g2_decap_8
XFILLER_5_282 VPWR VGND sg13g2_fill_1
X_2452_ VGND VPWR net741 net721 _1869_ _1579_ sg13g2_a21oi_1
X_2383_ VGND VPWR net733 _1800_ net721 _1693_ sg13g2_a21oi_2
XFILLER_39_2 VPWR VGND sg13g2_fill_1
X_4122_ _1465_ _1472_ u_ser.bit_pos\[2\] _1473_ VPWR VGND sg13g2_nand3_1
X_4053_ _1422_ _1353_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[7\]
+ _1348_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3004_ net709 net778 _0503_ VPWR VGND sg13g2_xor2_1
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_37_621 VPWR VGND sg13g2_decap_8
XFILLER_25_849 VPWR VGND sg13g2_decap_8
XFILLER_37_698 VPWR VGND sg13g2_decap_8
X_3906_ VGND VPWR _1502_ net645 _0148_ _1294_ sg13g2_a21oi_1
XFILLER_20_532 VPWR VGND sg13g2_decap_8
Xclkbuf_5_28__f_sap_3_inst.alu_inst.clk_regs clknet_4_14_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
X_3837_ _1244_ net673 _0870_ VPWR VGND sg13g2_nand2_1
X_3768_ net23 net15 net602 _1201_ VPWR VGND sg13g2_mux2_1
X_2719_ _0239_ VPWR _0249_ VGND _0243_ _0248_ sg13g2_o21ai_1
X_3699_ net670 net604 _1146_ VPWR VGND sg13g2_nor2_2
XFILLER_0_959 VPWR VGND sg13g2_decap_8
XFILLER_19_77 VPWR VGND sg13g2_fill_2
XFILLER_28_610 VPWR VGND sg13g2_decap_8
XFILLER_27_142 VPWR VGND sg13g2_fill_1
XFILLER_15_304 VPWR VGND sg13g2_fill_2
XFILLER_16_849 VPWR VGND sg13g2_decap_8
XFILLER_28_687 VPWR VGND sg13g2_decap_8
XFILLER_43_668 VPWR VGND sg13g2_decap_8
XFILLER_27_197 VPWR VGND sg13g2_fill_1
XFILLER_24_871 VPWR VGND sg13g2_decap_8
Xclkbuf_5_17__f_sap_3_inst.alu_inst.clk_regs clknet_4_8_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_11_565 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_1_sap_3_inst.alu_inst.clk clknet_1_1__leaf_sap_3_inst.alu_inst.clk clknet_leaf_1_sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_7_569 VPWR VGND sg13g2_decap_8
XFILLER_3_742 VPWR VGND sg13g2_decap_8
XFILLER_38_407 VPWR VGND sg13g2_fill_1
XFILLER_47_963 VPWR VGND sg13g2_decap_8
XFILLER_46_440 VPWR VGND sg13g2_decap_8
XFILLER_19_665 VPWR VGND sg13g2_decap_8
XFILLER_34_668 VPWR VGND sg13g2_decap_8
XFILLER_15_882 VPWR VGND sg13g2_decap_8
X_3622_ _1080_ net611 _1009_ VPWR VGND sg13g2_nand2_1
XFILLER_30_896 VPWR VGND sg13g2_decap_8
X_3553_ net571 net573 _0990_ _1017_ _1018_ VPWR VGND sg13g2_nor4_1
XFILLER_44_0 VPWR VGND sg13g2_fill_1
X_2504_ net667 net626 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[6\]
+ _1919_ VPWR VGND sg13g2_nand3_1
X_3484_ _0952_ _0813_ _0849_ VPWR VGND sg13g2_xnor2_1
X_2435_ VPWR VGND _1842_ _1793_ _1832_ net666 _1852_ net707 sg13g2_a221oi_1
X_2366_ _1783_ _1782_ _1672_ _1777_ _1692_ VPWR VGND sg13g2_a22oi_1
X_4105_ _1459_ VPWR _0182_ VGND _1442_ _1458_ sg13g2_o21ai_1
X_2297_ _1697_ _1701_ _1704_ _1707_ _1714_ VPWR VGND sg13g2_nor4_1
XFILLER_38_930 VPWR VGND sg13g2_decap_8
X_4036_ _1407_ _1349_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[5\]
+ net797 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_25_646 VPWR VGND sg13g2_decap_8
XFILLER_37_495 VPWR VGND sg13g2_decap_8
XFILLER_24_145 VPWR VGND sg13g2_fill_1
XFILLER_21_874 VPWR VGND sg13g2_decap_8
Xclkbuf_4_4_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_4_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_43_1025 VPWR VGND sg13g2_decap_4
XFILLER_48_738 VPWR VGND sg13g2_decap_8
XFILLER_44_911 VPWR VGND sg13g2_decap_8
XFILLER_43_410 VPWR VGND sg13g2_fill_2
XFILLER_28_484 VPWR VGND sg13g2_decap_8
XFILLER_29_985 VPWR VGND sg13g2_decap_8
XFILLER_16_646 VPWR VGND sg13g2_decap_8
XFILLER_44_988 VPWR VGND sg13g2_decap_8
XFILLER_43_465 VPWR VGND sg13g2_decap_8
XFILLER_31_649 VPWR VGND sg13g2_decap_8
XFILLER_8_801 VPWR VGND sg13g2_decap_8
XFILLER_12_863 VPWR VGND sg13g2_decap_8
XFILLER_8_878 VPWR VGND sg13g2_decap_8
X_2220_ VGND VPWR _1632_ _1637_ _1635_ _1633_ sg13g2_a21oi_2
X_2151_ _1560_ net750 _1568_ VPWR VGND sg13g2_nor2_1
XFILLER_16_4 VPWR VGND sg13g2_fill_2
XFILLER_47_760 VPWR VGND sg13g2_decap_8
X_2082_ VPWR _1500_ net788 VGND sg13g2_inv_1
XFILLER_35_911 VPWR VGND sg13g2_decap_8
XFILLER_35_988 VPWR VGND sg13g2_decap_8
X_2984_ _0483_ VPWR _0484_ VGND _0349_ _0482_ sg13g2_o21ai_1
XFILLER_22_627 VPWR VGND sg13g2_decap_8
XFILLER_30_693 VPWR VGND sg13g2_decap_8
X_3605_ net588 _0931_ _1066_ VPWR VGND sg13g2_nor2_1
X_3536_ _1002_ net588 _1001_ VPWR VGND sg13g2_nand2_2
X_3467_ _0935_ net662 _0933_ _0934_ VPWR VGND sg13g2_and3_1
X_2418_ _1659_ _1679_ net738 _1835_ VPWR VGND sg13g2_nand3_1
X_3398_ _0869_ _0770_ _0868_ VPWR VGND sg13g2_xnor2_1
X_2349_ net739 _1593_ _1764_ _1765_ _1766_ VPWR VGND sg13g2_nor4_1
XFILLER_45_708 VPWR VGND sg13g2_decap_8
XFILLER_29_259 VPWR VGND sg13g2_fill_2
X_4019_ _0154_ VPWR _1392_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[3\]
+ _1344_ sg13g2_o21ai_1
XFILLER_26_922 VPWR VGND sg13g2_decap_8
XFILLER_25_443 VPWR VGND sg13g2_decap_8
XFILLER_26_999 VPWR VGND sg13g2_decap_8
XFILLER_41_936 VPWR VGND sg13g2_decap_8
XFILLER_13_627 VPWR VGND sg13g2_decap_8
XFILLER_21_671 VPWR VGND sg13g2_decap_8
XFILLER_32_66 VPWR VGND sg13g2_fill_2
XFILLER_10_1024 VPWR VGND sg13g2_decap_4
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_535 VPWR VGND sg13g2_decap_8
XFILLER_36_708 VPWR VGND sg13g2_decap_8
XFILLER_29_782 VPWR VGND sg13g2_decap_8
XFILLER_17_933 VPWR VGND sg13g2_decap_8
XFILLER_44_785 VPWR VGND sg13g2_decap_8
XFILLER_32_903 VPWR VGND sg13g2_decap_8
XFILLER_12_660 VPWR VGND sg13g2_decap_8
XFILLER_8_675 VPWR VGND sg13g2_decap_8
X_3321_ _0792_ net639 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[5\]
+ net649 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[5\] VPWR VGND
+ sg13g2_a22oi_1
X_3252_ VGND VPWR net725 _1733_ _0723_ _1660_ sg13g2_a21oi_1
XFILLER_26_1020 VPWR VGND sg13g2_decap_8
X_3183_ VGND VPWR net752 _1627_ _0654_ _1777_ sg13g2_a21oi_1
X_2203_ _1618_ _1619_ _1620_ VPWR VGND sg13g2_nor2_2
X_2134_ net745 net744 _1551_ VPWR VGND sg13g2_nor2_2
XFILLER_39_557 VPWR VGND sg13g2_decap_8
XFILLER_26_218 VPWR VGND sg13g2_fill_2
XFILLER_23_914 VPWR VGND sg13g2_decap_8
XFILLER_35_785 VPWR VGND sg13g2_decap_8
XFILLER_33_1002 VPWR VGND sg13g2_decap_8
X_2967_ net598 net783 _0467_ _0036_ VPWR VGND sg13g2_a21o_1
X_2898_ _0400_ _0372_ net694 _0401_ VPWR VGND sg13g2_a21o_1
XFILLER_30_490 VPWR VGND sg13g2_decap_8
X_3519_ _0983_ _0984_ net662 _0985_ VPWR VGND sg13g2_nand3_1
XFILLER_40_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_1017 VPWR VGND sg13g2_decap_8
XFILLER_45_505 VPWR VGND sg13g2_decap_8
XFILLER_27_22 VPWR VGND sg13g2_fill_1
XFILLER_41_733 VPWR VGND sg13g2_decap_8
XFILLER_14_947 VPWR VGND sg13g2_decap_8
XFILLER_26_796 VPWR VGND sg13g2_decap_8
XFILLER_43_65 VPWR VGND sg13g2_fill_1
XFILLER_40_232 VPWR VGND sg13g2_fill_1
XFILLER_40_221 VPWR VGND sg13g2_decap_4
XFILLER_43_76 VPWR VGND sg13g2_fill_1
XFILLER_40_276 VPWR VGND sg13g2_fill_1
XFILLER_9_439 VPWR VGND sg13g2_fill_1
XFILLER_22_991 VPWR VGND sg13g2_decap_8
XFILLER_5_667 VPWR VGND sg13g2_decap_8
XFILLER_4_199 VPWR VGND sg13g2_fill_1
XFILLER_49_811 VPWR VGND sg13g2_decap_8
XFILLER_1_884 VPWR VGND sg13g2_decap_8
XFILLER_48_332 VPWR VGND sg13g2_decap_8
XFILLER_49_888 VPWR VGND sg13g2_decap_8
XFILLER_36_505 VPWR VGND sg13g2_decap_8
XFILLER_17_730 VPWR VGND sg13g2_decap_8
XFILLER_32_700 VPWR VGND sg13g2_decap_8
XFILLER_44_582 VPWR VGND sg13g2_decap_8
X_3870_ _1270_ VPWR _1271_ VGND _1268_ _1269_ sg13g2_o21ai_1
XFILLER_20_917 VPWR VGND sg13g2_decap_8
X_2821_ _0325_ _0324_ _1877_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_254 VPWR VGND sg13g2_fill_1
XFILLER_32_777 VPWR VGND sg13g2_decap_8
X_2752_ _0279_ _1612_ _1607_ VPWR VGND sg13g2_nand2b_1
XFILLER_13_991 VPWR VGND sg13g2_decap_8
XFILLER_8_472 VPWR VGND sg13g2_decap_8
XFILLER_9_984 VPWR VGND sg13g2_decap_8
X_2683_ _0215_ _0212_ _0213_ _0214_ VPWR VGND sg13g2_and3_1
X_3304_ _0775_ net669 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[7\]
+ net686 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[7\] VPWR VGND sg13g2_a22oi_1
X_4284_ net831 VGND VPWR _0141_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[3\]
+ clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3235_ VPWR VGND _1759_ _0705_ _0699_ net741 _0706_ _1775_ sg13g2_a221oi_1
X_3166_ _0637_ _0636_ _1634_ _1776_ _1646_ VPWR VGND sg13g2_a22oi_1
X_2117_ VPWR _1535_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[4\]
+ VGND sg13g2_inv_1
X_3097_ VGND VPWR sap_3_inst.alu_inst.act\[7\] net703 _0594_ net694 sg13g2_a21oi_1
XFILLER_23_711 VPWR VGND sg13g2_decap_8
XFILLER_35_582 VPWR VGND sg13g2_decap_8
XFILLER_23_788 VPWR VGND sg13g2_decap_8
X_3999_ _1373_ _1348_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[2\]
+ net797 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_2_659 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_fill_1
XFILLER_1_169 VPWR VGND sg13g2_fill_1
Xclkbuf_4_12_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs
+ clknet_4_12_0_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_46_825 VPWR VGND sg13g2_decap_8
XFILLER_45_379 VPWR VGND sg13g2_decap_8
XFILLER_33_519 VPWR VGND sg13g2_decap_8
XFILLER_41_530 VPWR VGND sg13g2_decap_8
XFILLER_14_744 VPWR VGND sg13g2_decap_8
XFILLER_26_593 VPWR VGND sg13g2_decap_8
XFILLER_10_961 VPWR VGND sg13g2_decap_8
Xclkload17 VPWR clkload17/Y clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs VGND sg13g2_inv_1
XFILLER_6_932 VPWR VGND sg13g2_decap_8
XFILLER_5_464 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_fill_2
XFILLER_1_681 VPWR VGND sg13g2_decap_8
XFILLER_23_1012 VPWR VGND sg13g2_decap_8
XFILLER_49_685 VPWR VGND sg13g2_decap_8
X_3020_ _0518_ _0508_ _0519_ VPWR VGND sg13g2_xor2_1
XFILLER_37_803 VPWR VGND sg13g2_decap_8
X_3922_ _1027_ _1306_ _1307_ VPWR VGND sg13g2_nor2_1
XFILLER_20_714 VPWR VGND sg13g2_decap_8
XFILLER_32_574 VPWR VGND sg13g2_decap_8
X_3853_ _1257_ _0303_ net673 VPWR VGND sg13g2_nand2_1
X_2804_ VGND VPWR net740 _0317_ _0318_ _1589_ sg13g2_a21oi_1
XFILLER_9_781 VPWR VGND sg13g2_decap_8
X_3784_ _0107_ _1213_ _1063_ net580 _1516_ VPWR VGND sg13g2_a22oi_1
X_2735_ net785 net788 net791 net793 _0264_ VPWR VGND sg13g2_nor4_1
X_2666_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[3\] net620
+ net601 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[3\] _0200_ net712
+ sg13g2_a221oi_1
XFILLER_5_80 VPWR VGND sg13g2_fill_1
X_4336_ net818 VGND VPWR _0193_ u_ser.bit_pos\[0\] clknet_3_1__leaf_clk sg13g2_dfrbpq_1
X_2597_ _1494_ _1571_ net728 _1616_ _2006_ VPWR VGND sg13g2_nor4_1
X_4267_ net819 VGND VPWR _0124_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[2\]
+ clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4198_ net821 VGND VPWR _0055_ sap_3_inst.alu_inst.tmp\[5\] clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
X_3218_ _0689_ _0644_ _1557_ net737 net743 VPWR VGND sg13g2_a22oi_1
X_3149_ _0624_ VPWR _0061_ VGND _1493_ net717 sg13g2_o21ai_1
XFILLER_28_869 VPWR VGND sg13g2_decap_8
XFILLER_11_747 VPWR VGND sg13g2_decap_8
XFILLER_23_585 VPWR VGND sg13g2_decap_8
XFILLER_10_268 VPWR VGND sg13g2_fill_2
XFILLER_3_924 VPWR VGND sg13g2_decap_8
XFILLER_2_456 VPWR VGND sg13g2_decap_8
Xfanout760 net761 net760 VPWR VGND sg13g2_buf_8
Xfanout793 sap_3_inst.alu_inst.acc\[0\] net793 VPWR VGND sg13g2_buf_8
XFILLER_1_38 VPWR VGND sg13g2_fill_2
Xfanout771 sap_3_inst.controller_inst.opcode\[0\] net771 VPWR VGND sg13g2_buf_2
Xfanout782 sap_3_inst.alu_inst.acc\[4\] net782 VPWR VGND sg13g2_buf_8
XFILLER_46_622 VPWR VGND sg13g2_decap_8
XFILLER_19_847 VPWR VGND sg13g2_decap_8
XFILLER_46_699 VPWR VGND sg13g2_decap_8
XFILLER_14_541 VPWR VGND sg13g2_decap_8
X_2520_ _1935_ _1933_ _1934_ VPWR VGND sg13g2_nand2_1
X_2451_ VGND VPWR _1868_ _1867_ _1768_ sg13g2_or2_1
X_2382_ net724 _1725_ _1799_ VPWR VGND sg13g2_nor2_1
X_4121_ _1469_ VPWR _1472_ VGND u_ser.bit_pos\[1\] _1471_ sg13g2_o21ai_1
X_4052_ _1421_ VPWR _0167_ VGND _1550_ _0154_ sg13g2_o21ai_1
XFILLER_37_600 VPWR VGND sg13g2_decap_8
XFILLER_49_482 VPWR VGND sg13g2_decap_8
X_3003_ _0502_ net778 net709 VPWR VGND sg13g2_nand2_1
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
XFILLER_37_677 VPWR VGND sg13g2_decap_8
XFILLER_25_828 VPWR VGND sg13g2_decap_8
X_3905_ VPWR VGND _1293_ _1292_ _0928_ net595 _1294_ _0917_ sg13g2_a221oi_1
XFILLER_33_883 VPWR VGND sg13g2_decap_8
XFILLER_20_511 VPWR VGND sg13g2_decap_8
X_3836_ _1243_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[0\] net654
+ VPWR VGND sg13g2_nand2_1
X_3767_ _1027_ _1199_ _1200_ VPWR VGND sg13g2_nor2_1
XFILLER_20_588 VPWR VGND sg13g2_decap_8
XFILLER_3_209 VPWR VGND sg13g2_fill_1
X_2718_ _0245_ _0246_ _0244_ _0248_ VPWR VGND _0247_ sg13g2_nand4_1
X_3698_ _0089_ _1144_ _1145_ net636 _1548_ VPWR VGND sg13g2_a22oi_1
X_2649_ _2056_ _2010_ _2055_ VPWR VGND sg13g2_nand2_2
XFILLER_0_938 VPWR VGND sg13g2_decap_8
X_4319_ net816 VGND VPWR _0176_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[7\]
+ clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_28_666 VPWR VGND sg13g2_decap_8
XFILLER_16_828 VPWR VGND sg13g2_decap_8
XFILLER_43_647 VPWR VGND sg13g2_decap_8
XFILLER_24_850 VPWR VGND sg13g2_decap_8
XFILLER_11_544 VPWR VGND sg13g2_decap_8
XFILLER_7_548 VPWR VGND sg13g2_decap_8
XFILLER_3_721 VPWR VGND sg13g2_decap_8
XFILLER_3_798 VPWR VGND sg13g2_decap_8
XFILLER_47_942 VPWR VGND sg13g2_decap_8
Xfanout590 net591 net590 VPWR VGND sg13g2_buf_1
XFILLER_19_644 VPWR VGND sg13g2_decap_8
XFILLER_20_1015 VPWR VGND sg13g2_decap_8
XFILLER_46_496 VPWR VGND sg13g2_decap_8
XFILLER_22_809 VPWR VGND sg13g2_decap_8
XFILLER_34_647 VPWR VGND sg13g2_decap_8
XFILLER_15_861 VPWR VGND sg13g2_decap_8
XFILLER_30_875 VPWR VGND sg13g2_decap_8
X_3621_ _1079_ _1078_ _1002_ VPWR VGND sg13g2_nand2b_1
X_3552_ _1016_ VPWR _1017_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[6\]
+ net661 sg13g2_o21ai_1
X_2503_ _1918_ _1539_ net631 VPWR VGND sg13g2_nand2_1
X_3483_ _0951_ _0916_ _0940_ VPWR VGND sg13g2_xnor2_1
X_2434_ net696 net626 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[7\]
+ _1851_ VPWR VGND sg13g2_nand3_1
X_2365_ _1782_ _1644_ _1666_ VPWR VGND sg13g2_nand2_1
X_4104_ _1459_ sap_3_inst.alu_inst.act\[5\] net579 VPWR VGND sg13g2_nand2_1
X_2296_ _1698_ _1702_ _1711_ _1712_ _1713_ VPWR VGND sg13g2_nor4_1
X_4035_ _1406_ _1353_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[5\]
+ _1346_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_25_625 VPWR VGND sg13g2_decap_8
XFILLER_38_986 VPWR VGND sg13g2_decap_8
XFILLER_13_809 VPWR VGND sg13g2_decap_8
XFILLER_40_639 VPWR VGND sg13g2_decap_8
XFILLER_33_680 VPWR VGND sg13g2_decap_8
XFILLER_21_853 VPWR VGND sg13g2_decap_8
X_3819_ _1057_ _1058_ net634 _1234_ VPWR VGND sg13g2_nor3_1
XFILLER_4_529 VPWR VGND sg13g2_decap_8
XFILLER_43_1004 VPWR VGND sg13g2_decap_8
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_48_717 VPWR VGND sg13g2_decap_8
XFILLER_29_964 VPWR VGND sg13g2_decap_8
XFILLER_16_625 VPWR VGND sg13g2_decap_8
XFILLER_28_463 VPWR VGND sg13g2_decap_8
XFILLER_44_967 VPWR VGND sg13g2_decap_8
XFILLER_43_444 VPWR VGND sg13g2_decap_8
XFILLER_43_433 VPWR VGND sg13g2_fill_2
XFILLER_43_422 VPWR VGND sg13g2_decap_8
XFILLER_15_157 VPWR VGND sg13g2_fill_1
XFILLER_30_127 VPWR VGND sg13g2_fill_1
XFILLER_31_628 VPWR VGND sg13g2_decap_8
XFILLER_12_842 VPWR VGND sg13g2_decap_8
XFILLER_30_149 VPWR VGND sg13g2_fill_1
XFILLER_8_857 VPWR VGND sg13g2_decap_8
XFILLER_3_595 VPWR VGND sg13g2_decap_8
X_2150_ VGND VPWR _1567_ net750 net751 sg13g2_or2_1
XFILLER_39_739 VPWR VGND sg13g2_decap_8
X_2081_ VPWR _1499_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[3\]
+ VGND sg13g2_inv_1
XFILLER_38_249 VPWR VGND sg13g2_fill_1
XFILLER_35_967 VPWR VGND sg13g2_decap_8
XFILLER_22_606 VPWR VGND sg13g2_decap_8
X_2983_ _0361_ VPWR _0483_ VGND net782 sap_3_inst.alu_inst.tmp\[4\] sg13g2_o21ai_1
XFILLER_30_672 VPWR VGND sg13g2_decap_8
X_3604_ net19 _1064_ _1065_ VPWR VGND sg13g2_nor2_2
X_3535_ _1001_ _0863_ _1000_ VPWR VGND sg13g2_nand2_1
X_3466_ _0934_ net678 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[3\]
+ net682 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2417_ VGND VPWR net750 _1620_ _1834_ _1749_ sg13g2_a21oi_1
X_3397_ _0779_ net589 _0864_ _0868_ VPWR VGND sg13g2_nor3_2
X_2348_ net750 _1749_ _1765_ VPWR VGND sg13g2_nor2_1
X_2279_ VGND VPWR net724 _1693_ _1696_ _1646_ sg13g2_a21oi_1
XFILLER_26_901 VPWR VGND sg13g2_decap_8
X_4018_ _1386_ _1390_ _1391_ VPWR VGND sg13g2_nor2_1
XFILLER_38_783 VPWR VGND sg13g2_decap_8
XFILLER_25_422 VPWR VGND sg13g2_decap_8
XFILLER_41_915 VPWR VGND sg13g2_decap_8
XFILLER_13_606 VPWR VGND sg13g2_decap_8
XFILLER_16_46 VPWR VGND sg13g2_fill_2
XFILLER_26_978 VPWR VGND sg13g2_decap_8
XFILLER_25_499 VPWR VGND sg13g2_decap_8
XFILLER_21_650 VPWR VGND sg13g2_decap_8
XFILLER_4_304 VPWR VGND sg13g2_fill_2
XFILLER_10_1003 VPWR VGND sg13g2_decap_8
XFILLER_5_849 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_514 VPWR VGND sg13g2_decap_8
XFILLER_17_912 VPWR VGND sg13g2_decap_8
XFILLER_29_761 VPWR VGND sg13g2_decap_8
XFILLER_44_764 VPWR VGND sg13g2_decap_8
XFILLER_17_989 VPWR VGND sg13g2_decap_8
XFILLER_16_499 VPWR VGND sg13g2_decap_8
XFILLER_32_959 VPWR VGND sg13g2_decap_8
XFILLER_8_654 VPWR VGND sg13g2_decap_8
X_3320_ _0791_ _0787_ _0788_ _0790_ VPWR VGND sg13g2_and3_1
XFILLER_4_893 VPWR VGND sg13g2_decap_8
X_3251_ _0722_ _0279_ _0684_ VPWR VGND sg13g2_nand2_1
X_2202_ _1605_ _1609_ _1596_ _1619_ VPWR VGND sg13g2_nand3_1
X_3182_ _0647_ _1567_ _0650_ _0653_ VPWR VGND sg13g2_a21o_2
XFILLER_39_536 VPWR VGND sg13g2_decap_8
XFILLER_35_764 VPWR VGND sg13g2_decap_8
XFILLER_22_425 VPWR VGND sg13g2_fill_2
X_2966_ net598 _0436_ _0466_ _0467_ VPWR VGND sg13g2_nor3_1
X_2897_ _0391_ _0392_ _0383_ _0400_ VPWR VGND _0399_ sg13g2_nand4_1
XFILLER_31_992 VPWR VGND sg13g2_decap_8
X_3518_ _0984_ net678 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[5\]
+ net687 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[5\] VPWR VGND sg13g2_a22oi_1
X_3449_ net660 _0917_ _0918_ VPWR VGND sg13g2_nor2_1
XFILLER_38_580 VPWR VGND sg13g2_decap_8
XFILLER_26_775 VPWR VGND sg13g2_decap_8
XFILLER_41_712 VPWR VGND sg13g2_decap_8
XFILLER_13_414 VPWR VGND sg13g2_fill_2
XFILLER_14_926 VPWR VGND sg13g2_decap_8
XFILLER_41_789 VPWR VGND sg13g2_decap_8
XFILLER_22_970 VPWR VGND sg13g2_decap_8
XFILLER_5_646 VPWR VGND sg13g2_decap_8
XFILLER_4_123 VPWR VGND sg13g2_fill_2
XFILLER_49_1021 VPWR VGND sg13g2_decap_8
XFILLER_4_27 VPWR VGND sg13g2_fill_1
XFILLER_1_863 VPWR VGND sg13g2_decap_8
XFILLER_48_311 VPWR VGND sg13g2_decap_8
XFILLER_49_867 VPWR VGND sg13g2_decap_8
XFILLER_48_388 VPWR VGND sg13g2_decap_8
XFILLER_44_561 VPWR VGND sg13g2_decap_8
XFILLER_17_786 VPWR VGND sg13g2_decap_8
XFILLER_32_756 VPWR VGND sg13g2_decap_8
X_2820_ VPWR VGND _1731_ _0322_ _0323_ _1761_ _0324_ _1875_ sg13g2_a221oi_1
XFILLER_13_970 VPWR VGND sg13g2_decap_8
X_2751_ _1670_ VPWR _0278_ VGND _0275_ _0277_ sg13g2_o21ai_1
XFILLER_9_963 VPWR VGND sg13g2_decap_8
X_2682_ _0214_ net617 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[2\]
+ net601 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_4_690 VPWR VGND sg13g2_decap_8
X_4283_ net827 VGND VPWR _0140_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[2\]
+ clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3303_ _0774_ net680 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[7\]
+ net683 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[7\] VPWR VGND sg13g2_a22oi_1
X_3234_ VGND VPWR _0703_ _0704_ _0705_ _1656_ sg13g2_a21oi_1
X_3165_ _1645_ _1692_ net761 _0636_ VPWR VGND sg13g2_nand3_1
X_2116_ VPWR _1534_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[4\]
+ VGND sg13g2_inv_1
X_3096_ _0592_ VPWR _0593_ VGND net575 _0575_ sg13g2_o21ai_1
XFILLER_27_539 VPWR VGND sg13g2_decap_8
XFILLER_35_561 VPWR VGND sg13g2_decap_8
XFILLER_23_767 VPWR VGND sg13g2_decap_8
XFILLER_11_929 VPWR VGND sg13g2_decap_8
X_3998_ net798 net66 _1372_ _0162_ VPWR VGND sg13g2_a21o_1
X_2949_ _0450_ _0448_ _0449_ VPWR VGND sg13g2_nand2_1
XFILLER_2_638 VPWR VGND sg13g2_decap_8
XFILLER_46_804 VPWR VGND sg13g2_decap_8
XFILLER_45_358 VPWR VGND sg13g2_decap_8
XFILLER_14_723 VPWR VGND sg13g2_decap_8
XFILLER_26_572 VPWR VGND sg13g2_decap_8
XFILLER_41_586 VPWR VGND sg13g2_decap_8
XFILLER_9_226 VPWR VGND sg13g2_fill_2
XFILLER_6_911 VPWR VGND sg13g2_decap_8
XFILLER_10_940 VPWR VGND sg13g2_decap_8
Xclkload18 clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs clkload18/X VPWR VGND sg13g2_buf_1
XFILLER_6_988 VPWR VGND sg13g2_decap_8
XFILLER_1_660 VPWR VGND sg13g2_decap_8
XFILLER_49_664 VPWR VGND sg13g2_decap_8
XFILLER_37_859 VPWR VGND sg13g2_decap_8
XFILLER_17_583 VPWR VGND sg13g2_decap_8
X_3921_ net592 VPWR _1306_ VGND net647 _1028_ sg13g2_o21ai_1
XFILLER_32_553 VPWR VGND sg13g2_decap_8
X_3852_ VGND VPWR _0927_ _0940_ _1256_ _0881_ sg13g2_a21oi_1
X_2803_ _1590_ VPWR _0317_ VGND _1599_ _0316_ sg13g2_o21ai_1
XFILLER_9_760 VPWR VGND sg13g2_decap_8
X_3783_ _1060_ net580 _1213_ VPWR VGND sg13g2_nor2_1
X_2734_ net774 net780 net782 net777 _0263_ VPWR VGND sg13g2_nor4_1
X_2665_ _0199_ _0197_ _0198_ VPWR VGND sg13g2_nand2_1
X_2596_ _2005_ net757 _1996_ VPWR VGND sg13g2_nand2_2
X_4335_ net831 VGND VPWR _0192_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[3\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_2
XFILLER_8_1018 VPWR VGND sg13g2_decap_8
X_4266_ net820 VGND VPWR _0123_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[1\]
+ clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3217_ _0288_ VPWR _0688_ VGND _1621_ _0687_ sg13g2_o21ai_1
X_4197_ net823 VGND VPWR _0054_ sap_3_inst.alu_inst.tmp\[4\] clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
X_3148_ _0624_ net717 net32 VPWR VGND sg13g2_nand2_1
XFILLER_28_848 VPWR VGND sg13g2_decap_8
XFILLER_43_829 VPWR VGND sg13g2_decap_8
X_3079_ _0576_ _0557_ _0575_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_564 VPWR VGND sg13g2_decap_8
XFILLER_11_726 VPWR VGND sg13g2_decap_8
Xclkbuf_5_30__f_sap_3_inst.alu_inst.clk_regs clknet_4_15_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_3_903 VPWR VGND sg13g2_decap_8
XFILLER_49_98 VPWR VGND sg13g2_fill_2
Xfanout750 _1565_ net750 VPWR VGND sg13g2_buf_8
XFILLER_46_601 VPWR VGND sg13g2_decap_8
Xfanout794 _1343_ net794 VPWR VGND sg13g2_buf_8
Xfanout772 net773 net772 VPWR VGND sg13g2_buf_8
Xfanout783 net785 net783 VPWR VGND sg13g2_buf_8
Xfanout761 sap_3_inst.controller_inst.opcode\[4\] net761 VPWR VGND sg13g2_buf_8
XFILLER_19_826 VPWR VGND sg13g2_decap_8
XFILLER_46_678 VPWR VGND sg13g2_decap_8
XFILLER_45_166 VPWR VGND sg13g2_fill_1
XFILLER_34_829 VPWR VGND sg13g2_decap_8
XFILLER_14_520 VPWR VGND sg13g2_decap_8
XFILLER_42_884 VPWR VGND sg13g2_decap_8
XFILLER_14_597 VPWR VGND sg13g2_decap_8
Xclkbuf_4_5_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_5_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_6_785 VPWR VGND sg13g2_decap_8
X_2450_ _1846_ VPWR _1867_ VGND _1855_ _1866_ sg13g2_o21ai_1
X_2381_ _1654_ VPWR _1798_ VGND _1705_ _1797_ sg13g2_o21ai_1
X_4120_ _1470_ VPWR _1471_ VGND net800 u_ser.shadow_reg\[5\] sg13g2_o21ai_1
X_4051_ _1420_ VPWR _1421_ VGND _1417_ _1419_ sg13g2_o21ai_1
XFILLER_49_461 VPWR VGND sg13g2_decap_8
X_3002_ net708 net782 _0471_ _0501_ VPWR VGND sg13g2_a21o_1
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
XFILLER_25_807 VPWR VGND sg13g2_decap_8
XFILLER_37_656 VPWR VGND sg13g2_decap_8
X_3904_ VGND VPWR net643 _0931_ _1293_ net587 sg13g2_a21oi_1
XFILLER_33_862 VPWR VGND sg13g2_decap_8
X_3835_ net634 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[7\] _1242_
+ _0129_ VPWR VGND sg13g2_a21o_1
XFILLER_20_567 VPWR VGND sg13g2_decap_8
X_3766_ net592 VPWR _1199_ VGND net676 _1028_ sg13g2_o21ai_1
X_2717_ net697 net627 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[0\]
+ _0247_ VPWR VGND sg13g2_nand3_1
X_3697_ _1145_ net608 _1045_ VPWR VGND sg13g2_nand2_1
XFILLER_10_48 VPWR VGND sg13g2_fill_2
X_2648_ _2055_ _2012_ _2054_ VPWR VGND sg13g2_nand2_2
X_2579_ net576 VPWR _1990_ VGND _1984_ _1989_ sg13g2_o21ai_1
XFILLER_0_917 VPWR VGND sg13g2_decap_8
X_4318_ net812 VGND VPWR _0175_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[6\]
+ clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4249_ net827 VGND VPWR _0106_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[0\]
+ clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_16_807 VPWR VGND sg13g2_decap_8
XFILLER_28_645 VPWR VGND sg13g2_decap_8
XFILLER_43_626 VPWR VGND sg13g2_decap_8
XFILLER_11_523 VPWR VGND sg13g2_decap_8
Xclkbuf_5_8__f_sap_3_inst.alu_inst.clk_regs clknet_4_4_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_7_527 VPWR VGND sg13g2_decap_8
XFILLER_13_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_700 VPWR VGND sg13g2_decap_8
XFILLER_3_777 VPWR VGND sg13g2_decap_8
XFILLER_47_921 VPWR VGND sg13g2_decap_8
Xfanout580 net581 net580 VPWR VGND sg13g2_buf_8
XFILLER_19_623 VPWR VGND sg13g2_decap_8
Xfanout591 _0825_ net591 VPWR VGND sg13g2_buf_8
XFILLER_47_998 VPWR VGND sg13g2_decap_8
XFILLER_46_475 VPWR VGND sg13g2_decap_8
XFILLER_34_626 VPWR VGND sg13g2_decap_8
XFILLER_15_840 VPWR VGND sg13g2_decap_8
XFILLER_42_681 VPWR VGND sg13g2_decap_8
XFILLER_30_854 VPWR VGND sg13g2_decap_8
X_3620_ net569 _1077_ _1078_ VPWR VGND sg13g2_and2_1
X_3551_ _1014_ _1015_ _1013_ _1016_ VPWR VGND sg13g2_nand3_1
X_2502_ VGND VPWR _1914_ _1915_ _0032_ _1917_ sg13g2_a21oi_1
XFILLER_6_582 VPWR VGND sg13g2_decap_8
X_3482_ _0780_ _0852_ _0892_ _0950_ VGND VPWR _0949_ sg13g2_nor4_2
X_2433_ net696 _1849_ _1850_ VPWR VGND sg13g2_and2_1
X_2364_ net733 _1780_ _1781_ VPWR VGND sg13g2_nor2_1
X_4103_ _1457_ VPWR _1458_ VGND net779 net699 sg13g2_o21ai_1
X_2295_ _1712_ _1693_ _1631_ _1646_ _1640_ VPWR VGND sg13g2_a22oi_1
XFILLER_38_965 VPWR VGND sg13g2_decap_8
X_4034_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[5\] _1348_
+ _1405_ net795 sg13g2_a21oi_1
XFILLER_25_604 VPWR VGND sg13g2_decap_8
X_4146__4 VPWR net38 clknet_leaf_1_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
XFILLER_40_618 VPWR VGND sg13g2_decap_8
XFILLER_21_832 VPWR VGND sg13g2_decap_8
XFILLER_36_1023 VPWR VGND sg13g2_decap_4
X_3818_ VGND VPWR net688 _1233_ _1705_ _1659_ sg13g2_a21oi_2
XFILLER_4_508 VPWR VGND sg13g2_decap_8
X_3749_ _1184_ VPWR _1185_ VGND net20 net603 sg13g2_o21ai_1
XFILLER_0_714 VPWR VGND sg13g2_decap_8
XFILLER_29_943 VPWR VGND sg13g2_decap_8
XFILLER_16_604 VPWR VGND sg13g2_decap_8
XFILLER_44_946 VPWR VGND sg13g2_decap_8
XFILLER_31_607 VPWR VGND sg13g2_decap_8
XFILLER_12_821 VPWR VGND sg13g2_decap_8
XFILLER_30_139 VPWR VGND sg13g2_fill_1
XFILLER_8_836 VPWR VGND sg13g2_decap_8
XFILLER_12_898 VPWR VGND sg13g2_decap_8
XFILLER_7_335 VPWR VGND sg13g2_fill_2
XFILLER_3_574 VPWR VGND sg13g2_decap_8
XFILLER_39_718 VPWR VGND sg13g2_decap_8
X_2080_ VPWR _1498_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[3\]
+ VGND sg13g2_inv_1
XFILLER_47_795 VPWR VGND sg13g2_decap_8
XFILLER_46_283 VPWR VGND sg13g2_decap_8
XFILLER_19_497 VPWR VGND sg13g2_decap_8
XFILLER_35_946 VPWR VGND sg13g2_decap_8
XFILLER_43_990 VPWR VGND sg13g2_decap_8
X_2982_ _0481_ _0479_ _0482_ VPWR VGND sg13g2_xor2_1
XFILLER_30_651 VPWR VGND sg13g2_decap_8
X_3603_ net613 _0919_ _1064_ VPWR VGND sg13g2_nor2_2
XFILLER_7_891 VPWR VGND sg13g2_decap_8
X_3534_ VGND VPWR _0793_ _0862_ _1000_ net585 sg13g2_a21oi_1
X_3465_ _0933_ net685 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[3\]
+ net687 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2416_ net752 _1635_ net715 _1692_ _1833_ VPWR VGND sg13g2_and4_1
X_3396_ net589 _0863_ _0867_ VPWR VGND sg13g2_nor2_1
X_2347_ VPWR VGND _1597_ net719 _1763_ _1743_ _1764_ _1757_ sg13g2_a221oi_1
X_2278_ _1694_ _1670_ _1691_ _1695_ VPWR VGND sg13g2_a21o_1
X_4017_ _1387_ _1388_ _1383_ _1390_ VPWR VGND _1389_ sg13g2_nand4_1
XFILLER_38_762 VPWR VGND sg13g2_decap_8
XFILLER_26_957 VPWR VGND sg13g2_decap_8
XFILLER_25_478 VPWR VGND sg13g2_decap_8
XFILLER_34_990 VPWR VGND sg13g2_decap_8
XFILLER_5_828 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_29_740 VPWR VGND sg13g2_decap_8
XFILLER_44_743 VPWR VGND sg13g2_decap_8
XFILLER_17_968 VPWR VGND sg13g2_decap_8
XFILLER_16_478 VPWR VGND sg13g2_decap_8
XFILLER_32_938 VPWR VGND sg13g2_decap_8
XFILLER_40_982 VPWR VGND sg13g2_decap_8
XFILLER_8_633 VPWR VGND sg13g2_decap_8
XFILLER_12_695 VPWR VGND sg13g2_decap_8
XFILLER_4_872 VPWR VGND sg13g2_decap_8
X_3250_ VGND VPWR net726 net720 _0721_ _0670_ sg13g2_a21oi_1
Xclkbuf_4_13_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs
+ clknet_4_13_0_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
X_2201_ _1571_ _1617_ _1618_ VPWR VGND sg13g2_nor2_1
X_3181_ VGND VPWR _0650_ _0652_ _0647_ net740 sg13g2_a21oi_2
XFILLER_39_515 VPWR VGND sg13g2_decap_8
X_2132_ VPWR _1550_ net52 VGND sg13g2_inv_1
XFILLER_47_592 VPWR VGND sg13g2_decap_8
XFILLER_35_743 VPWR VGND sg13g2_decap_8
XFILLER_23_949 VPWR VGND sg13g2_decap_8
XFILLER_22_459 VPWR VGND sg13g2_decap_8
X_2965_ VPWR VGND _0465_ net693 _0464_ sap_3_inst.alu_inst.act\[3\] _0466_ _0320_
+ sg13g2_a221oi_1
XFILLER_31_971 VPWR VGND sg13g2_decap_8
X_2896_ _0377_ _0396_ _0397_ _0398_ _0399_ VPWR VGND sg13g2_nor4_1
X_3517_ _0983_ net681 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[5\]
+ net684 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[5\] VPWR VGND sg13g2_a22oi_1
X_3448_ _0917_ _0893_ _0915_ VPWR VGND sg13g2_xnor2_1
X_3379_ _0813_ net591 _0836_ _0847_ _0850_ VPWR VGND sg13g2_and4_1
XFILLER_27_68 VPWR VGND sg13g2_fill_1
XFILLER_14_905 VPWR VGND sg13g2_decap_8
XFILLER_26_754 VPWR VGND sg13g2_decap_8
XFILLER_40_201 VPWR VGND sg13g2_fill_1
XFILLER_41_768 VPWR VGND sg13g2_decap_8
XFILLER_49_1000 VPWR VGND sg13g2_decap_8
XFILLER_5_625 VPWR VGND sg13g2_decap_8
XFILLER_1_842 VPWR VGND sg13g2_decap_8
XFILLER_49_846 VPWR VGND sg13g2_decap_8
XFILLER_48_367 VPWR VGND sg13g2_decap_8
XFILLER_1_1024 VPWR VGND sg13g2_decap_4
XFILLER_44_540 VPWR VGND sg13g2_decap_8
XFILLER_17_765 VPWR VGND sg13g2_decap_8
XFILLER_31_212 VPWR VGND sg13g2_fill_2
XFILLER_32_735 VPWR VGND sg13g2_decap_8
X_2750_ _0276_ VPWR _0277_ VGND _1666_ _1676_ sg13g2_o21ai_1
XFILLER_9_942 VPWR VGND sg13g2_decap_8
XFILLER_31_278 VPWR VGND sg13g2_fill_1
XFILLER_12_492 VPWR VGND sg13g2_decap_8
X_2681_ _0213_ net600 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[2\]
+ net619 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[2\] VPWR VGND
+ sg13g2_a22oi_1
X_4282_ net806 VGND VPWR _0139_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[1\]
+ clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3302_ _0773_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[7\] net641
+ VPWR VGND sg13g2_nand2_1
X_3233_ _0704_ net730 net719 VPWR VGND sg13g2_nand2_1
X_3164_ _0635_ _1762_ _1875_ VPWR VGND sg13g2_nand2_1
XFILLER_27_518 VPWR VGND sg13g2_decap_8
X_2115_ VPWR _1533_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[4\]
+ VGND sg13g2_inv_1
X_3095_ net703 _0591_ _0592_ VPWR VGND sg13g2_nor2_1
XFILLER_35_540 VPWR VGND sg13g2_decap_8
XFILLER_23_746 VPWR VGND sg13g2_decap_8
XFILLER_11_908 VPWR VGND sg13g2_decap_8
X_3997_ VPWR VGND _1371_ net798 _1370_ _1510_ _1372_ net794 sg13g2_a221oi_1
X_2948_ _0449_ net691 net781 net692 net786 VPWR VGND sg13g2_a22oi_1
XFILLER_13_48 VPWR VGND sg13g2_fill_1
X_2879_ _0348_ VPWR _0382_ VGND _0380_ _0381_ sg13g2_o21ai_1
XFILLER_2_617 VPWR VGND sg13g2_decap_8
XFILLER_18_529 VPWR VGND sg13g2_decap_8
XFILLER_14_702 VPWR VGND sg13g2_decap_8
XFILLER_26_551 VPWR VGND sg13g2_decap_8
XFILLER_41_565 VPWR VGND sg13g2_decap_8
XFILLER_14_779 VPWR VGND sg13g2_decap_8
XFILLER_16_1010 VPWR VGND sg13g2_decap_8
XFILLER_10_996 VPWR VGND sg13g2_decap_8
Xclkload19 VPWR clkload19/Y clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs VGND sg13g2_inv_1
XFILLER_6_967 VPWR VGND sg13g2_decap_8
XFILLER_5_499 VPWR VGND sg13g2_decap_8
XFILLER_49_643 VPWR VGND sg13g2_decap_8
XFILLER_37_838 VPWR VGND sg13g2_decap_8
X_3920_ VGND VPWR _1536_ net643 _0151_ _1305_ sg13g2_a21oi_1
XFILLER_17_562 VPWR VGND sg13g2_decap_8
XFILLER_32_532 VPWR VGND sg13g2_decap_8
X_3851_ net654 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[2\] _1255_
+ _0132_ VPWR VGND sg13g2_a21o_1
X_2802_ VGND VPWR _1620_ _0315_ _0316_ _1622_ sg13g2_a21oi_1
XFILLER_20_749 VPWR VGND sg13g2_decap_8
X_3782_ net580 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[0\] _1212_
+ _0106_ VPWR VGND sg13g2_a21o_1
X_2733_ _0254_ _0262_ _0250_ net17 VPWR VGND sg13g2_nand3_1
X_2664_ _0198_ net616 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[3\]
+ net625 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2595_ net757 _1996_ _2004_ VPWR VGND sg13g2_and2_1
X_4334_ net830 VGND VPWR _0191_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[2\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_2
X_4265_ net827 VGND VPWR _0122_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[0\]
+ clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3216_ VGND VPWR _0679_ _0686_ _0687_ _0669_ sg13g2_a21oi_1
X_4196_ net823 VGND VPWR _0053_ sap_3_inst.alu_inst.tmp\[3\] clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
X_3147_ _0623_ VPWR _0060_ VGND _1494_ _1585_ sg13g2_o21ai_1
XFILLER_28_827 VPWR VGND sg13g2_decap_8
XFILLER_43_808 VPWR VGND sg13g2_decap_8
X_3078_ _0575_ _0573_ _0574_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_705 VPWR VGND sg13g2_decap_8
XFILLER_23_543 VPWR VGND sg13g2_decap_8
XFILLER_7_709 VPWR VGND sg13g2_decap_8
XFILLER_46_1014 VPWR VGND sg13g2_decap_8
XFILLER_3_959 VPWR VGND sg13g2_decap_8
XFILLER_49_88 VPWR VGND sg13g2_fill_1
Xfanout751 _1563_ net751 VPWR VGND sg13g2_buf_8
Xfanout740 _1567_ net740 VPWR VGND sg13g2_buf_8
Xfanout773 net774 net773 VPWR VGND sg13g2_buf_1
Xfanout762 net763 net762 VPWR VGND sg13g2_buf_8
Xfanout784 net785 net784 VPWR VGND sg13g2_buf_1
XFILLER_19_805 VPWR VGND sg13g2_decap_8
Xfanout795 _1343_ net795 VPWR VGND sg13g2_buf_1
XFILLER_46_657 VPWR VGND sg13g2_decap_8
XFILLER_34_808 VPWR VGND sg13g2_decap_8
XFILLER_27_882 VPWR VGND sg13g2_decap_8
XFILLER_42_863 VPWR VGND sg13g2_decap_8
XFILLER_14_576 VPWR VGND sg13g2_decap_8
XFILLER_6_764 VPWR VGND sg13g2_decap_8
XFILLER_10_793 VPWR VGND sg13g2_decap_8
X_2380_ net737 _1679_ _1797_ VPWR VGND sg13g2_and2_1
XFILLER_2_981 VPWR VGND sg13g2_decap_8
XFILLER_49_440 VPWR VGND sg13g2_decap_8
X_4050_ VGND VPWR _1539_ net794 _1420_ net798 sg13g2_a21oi_1
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
X_3001_ _0340_ net781 _0500_ _0037_ VPWR VGND sg13g2_a21o_1
XFILLER_36_101 VPWR VGND sg13g2_fill_2
XFILLER_37_635 VPWR VGND sg13g2_decap_8
XFILLER_24_318 VPWR VGND sg13g2_fill_2
XFILLER_18_893 VPWR VGND sg13g2_decap_8
XFILLER_33_841 VPWR VGND sg13g2_decap_8
X_3903_ _1292_ net648 net11 VPWR VGND sg13g2_nand2b_1
X_3834_ _1090_ _1092_ net634 _1242_ VPWR VGND sg13g2_nor3_1
XFILLER_20_546 VPWR VGND sg13g2_decap_8
X_3765_ _1198_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[6\] net656
+ VPWR VGND sg13g2_nand2_1
X_2716_ _0246_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[0\] net615
+ VPWR VGND sg13g2_nand2_1
X_3696_ net636 _1142_ _1143_ _1144_ VPWR VGND sg13g2_nor3_1
X_2647_ _2054_ _2017_ _2018_ VPWR VGND sg13g2_nand2_2
X_2578_ _1986_ _1987_ _1985_ _1989_ VPWR VGND _1988_ sg13g2_nand4_1
X_4317_ net830 VGND VPWR _0174_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[5\]
+ clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4248_ net809 VGND VPWR _0105_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[7\]
+ clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_28_624 VPWR VGND sg13g2_decap_8
X_4179_ net823 VGND VPWR _0036_ sap_3_inst.alu_inst.acc\[3\] clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_43_605 VPWR VGND sg13g2_decap_8
XFILLER_35_57 VPWR VGND sg13g2_fill_2
XFILLER_11_502 VPWR VGND sg13g2_decap_8
XFILLER_24_885 VPWR VGND sg13g2_decap_8
XFILLER_7_506 VPWR VGND sg13g2_decap_8
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_11_579 VPWR VGND sg13g2_decap_8
XFILLER_3_756 VPWR VGND sg13g2_decap_8
XFILLER_47_900 VPWR VGND sg13g2_decap_8
Xfanout592 net593 net592 VPWR VGND sg13g2_buf_8
XFILLER_19_602 VPWR VGND sg13g2_decap_8
Xfanout570 _1941_ net570 VPWR VGND sg13g2_buf_8
Xfanout581 _1211_ net581 VPWR VGND sg13g2_buf_8
XFILLER_47_977 VPWR VGND sg13g2_decap_8
XFILLER_46_454 VPWR VGND sg13g2_decap_8
XFILLER_18_145 VPWR VGND sg13g2_fill_1
XFILLER_19_679 VPWR VGND sg13g2_decap_8
XFILLER_34_605 VPWR VGND sg13g2_decap_8
XFILLER_42_660 VPWR VGND sg13g2_decap_8
XFILLER_15_896 VPWR VGND sg13g2_decap_8
XFILLER_30_833 VPWR VGND sg13g2_decap_8
X_3550_ _1015_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[6\] net669
+ VPWR VGND sg13g2_nand2_1
XFILLER_10_590 VPWR VGND sg13g2_decap_8
XFILLER_6_561 VPWR VGND sg13g2_decap_8
X_2501_ sap_3_inst.alu_flags\[7\] _1915_ _1917_ VPWR VGND sg13g2_nor2_1
X_3481_ _0949_ _0914_ _0940_ VPWR VGND sg13g2_nand2_1
X_2432_ VGND VPWR net666 net707 _1849_ _1844_ sg13g2_a21oi_1
XFILLER_29_1020 VPWR VGND sg13g2_decap_8
X_2363_ _1705_ _1731_ _1779_ _1780_ VPWR VGND sg13g2_nor3_1
X_4102_ _1457_ net699 _0515_ VPWR VGND sg13g2_nand2b_1
X_2294_ VGND VPWR net724 _1709_ _1711_ _1660_ sg13g2_a21oi_1
X_4033_ _1404_ _1340_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[5\]
+ net796 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_2_94 VPWR VGND sg13g2_decap_8
XFILLER_38_944 VPWR VGND sg13g2_decap_8
XFILLER_18_690 VPWR VGND sg13g2_decap_8
XFILLER_36_1002 VPWR VGND sg13g2_decap_8
XFILLER_21_811 VPWR VGND sg13g2_decap_8
XFILLER_21_888 VPWR VGND sg13g2_decap_8
X_3817_ _1231_ VPWR _0121_ VGND _1090_ _1232_ sg13g2_o21ai_1
X_3748_ _1184_ _0303_ net603 VPWR VGND sg13g2_nand2_1
X_3679_ net612 _0993_ _1126_ _1129_ VPWR VGND sg13g2_nor3_1
XFILLER_29_922 VPWR VGND sg13g2_decap_8
XFILLER_44_925 VPWR VGND sg13g2_decap_8
XFILLER_29_999 VPWR VGND sg13g2_decap_8
XFILLER_28_498 VPWR VGND sg13g2_decap_8
XFILLER_43_479 VPWR VGND sg13g2_decap_8
XFILLER_12_800 VPWR VGND sg13g2_decap_8
XFILLER_24_682 VPWR VGND sg13g2_decap_8
XFILLER_8_815 VPWR VGND sg13g2_decap_8
XFILLER_12_877 VPWR VGND sg13g2_decap_8
XFILLER_7_39 VPWR VGND sg13g2_fill_1
XFILLER_3_553 VPWR VGND sg13g2_decap_8
XFILLER_47_774 VPWR VGND sg13g2_decap_8
XFILLER_19_476 VPWR VGND sg13g2_decap_8
XFILLER_35_925 VPWR VGND sg13g2_decap_8
X_2981_ _0481_ _0413_ _0439_ VPWR VGND sg13g2_nand2_2
XFILLER_15_693 VPWR VGND sg13g2_decap_8
XFILLER_30_630 VPWR VGND sg13g2_decap_8
X_3602_ _0075_ _1061_ _1063_ net583 _1519_ VPWR VGND sg13g2_a22oi_1
XFILLER_7_870 VPWR VGND sg13g2_decap_8
X_3533_ VGND VPWR net569 net606 _0999_ _0998_ sg13g2_a21oi_1
X_3464_ _0906_ VPWR _0068_ VGND _0926_ _0932_ sg13g2_o21ai_1
X_2415_ _1832_ net739 _1831_ VPWR VGND sg13g2_nand2_2
X_3395_ VGND VPWR _0866_ _0862_ net591 sg13g2_or2_1
X_2346_ VGND VPWR net731 _1762_ _1763_ net716 sg13g2_a21oi_1
X_2277_ _1629_ _1692_ _1694_ VPWR VGND sg13g2_nor2_1
XFILLER_38_741 VPWR VGND sg13g2_decap_8
X_4016_ _1389_ _1348_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[3\]
+ _1346_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_26_936 VPWR VGND sg13g2_decap_8
XFILLER_25_457 VPWR VGND sg13g2_decap_8
XFILLER_20_162 VPWR VGND sg13g2_fill_2
XFILLER_21_685 VPWR VGND sg13g2_decap_8
XFILLER_5_807 VPWR VGND sg13g2_decap_8
XFILLER_4_306 VPWR VGND sg13g2_fill_1
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_48_549 VPWR VGND sg13g2_decap_8
XFILLER_44_722 VPWR VGND sg13g2_decap_8
XFILLER_17_947 VPWR VGND sg13g2_decap_8
XFILLER_28_284 VPWR VGND sg13g2_decap_4
XFILLER_29_796 VPWR VGND sg13g2_decap_8
XFILLER_44_799 VPWR VGND sg13g2_decap_8
XFILLER_32_917 VPWR VGND sg13g2_decap_8
XFILLER_40_961 VPWR VGND sg13g2_decap_8
XFILLER_8_612 VPWR VGND sg13g2_decap_8
XFILLER_12_674 VPWR VGND sg13g2_decap_8
XFILLER_8_689 VPWR VGND sg13g2_decap_8
XFILLER_4_851 VPWR VGND sg13g2_decap_8
X_4154__12 VPWR net46 clknet_leaf_0_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
X_2200_ net771 net765 net767 _1617_ VPWR VGND sg13g2_nand3_1
X_3180_ VPWR _0651_ _0650_ VGND sg13g2_inv_1
X_2131_ VPWR _1549_ net50 VGND sg13g2_inv_1
XFILLER_47_571 VPWR VGND sg13g2_decap_8
XFILLER_35_722 VPWR VGND sg13g2_decap_8
XFILLER_23_928 VPWR VGND sg13g2_decap_8
XFILLER_34_254 VPWR VGND sg13g2_fill_1
XFILLER_35_799 VPWR VGND sg13g2_decap_8
X_2964_ VGND VPWR _0353_ _0458_ _0465_ net702 sg13g2_a21oi_1
XFILLER_15_490 VPWR VGND sg13g2_decap_8
XFILLER_22_427 VPWR VGND sg13g2_fill_1
XFILLER_22_438 VPWR VGND sg13g2_decap_8
XFILLER_31_950 VPWR VGND sg13g2_decap_8
XFILLER_33_1016 VPWR VGND sg13g2_decap_8
X_2895_ _0382_ VPWR _0398_ VGND net789 _0335_ sg13g2_o21ai_1
XFILLER_33_1027 VPWR VGND sg13g2_fill_2
X_3516_ _0982_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[5\] net596
+ VPWR VGND sg13g2_nand2_1
X_3447_ _0916_ _0914_ _0893_ VPWR VGND sg13g2_nand2b_1
X_3378_ _0836_ _0847_ net591 _0849_ VPWR VGND sg13g2_nand3_1
X_2329_ VGND VPWR net726 _1736_ _1746_ _1745_ sg13g2_a21oi_1
XFILLER_45_519 VPWR VGND sg13g2_decap_8
XFILLER_27_36 VPWR VGND sg13g2_fill_2
XFILLER_26_733 VPWR VGND sg13g2_decap_8
XFILLER_25_254 VPWR VGND sg13g2_decap_4
XFILLER_41_747 VPWR VGND sg13g2_decap_8
XFILLER_9_409 VPWR VGND sg13g2_fill_2
XFILLER_21_482 VPWR VGND sg13g2_decap_8
XFILLER_5_604 VPWR VGND sg13g2_decap_8
XFILLER_1_821 VPWR VGND sg13g2_decap_8
XFILLER_49_825 VPWR VGND sg13g2_decap_8
XFILLER_1_898 VPWR VGND sg13g2_decap_8
XFILLER_48_346 VPWR VGND sg13g2_decap_8
XFILLER_1_1003 VPWR VGND sg13g2_decap_8
XFILLER_36_519 VPWR VGND sg13g2_decap_8
XFILLER_17_744 VPWR VGND sg13g2_decap_8
XFILLER_29_593 VPWR VGND sg13g2_decap_8
XFILLER_32_714 VPWR VGND sg13g2_decap_8
XFILLER_44_596 VPWR VGND sg13g2_decap_8
XFILLER_9_921 VPWR VGND sg13g2_decap_8
X_2680_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[2\] net630
+ net629 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[2\] _0212_ net711
+ sg13g2_a221oi_1
XFILLER_8_486 VPWR VGND sg13g2_decap_8
XFILLER_9_998 VPWR VGND sg13g2_decap_8
X_3301_ _0772_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[7\] net648
+ VPWR VGND sg13g2_nand2_1
X_4281_ net829 VGND VPWR _0138_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[0\]
+ clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3232_ VGND VPWR _0703_ _0702_ _0700_ sg13g2_or2_1
X_3163_ _0634_ net720 _1634_ _1666_ _1644_ VPWR VGND sg13g2_a22oi_1
X_2114_ VPWR _1532_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[4\]
+ VGND sg13g2_inv_1
X_3094_ VGND VPWR _2000_ _0569_ _0591_ _0590_ sg13g2_a21oi_1
XFILLER_23_725 VPWR VGND sg13g2_decap_8
XFILLER_35_596 VPWR VGND sg13g2_decap_8
Xclkbuf_4_6_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_6_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
X_3996_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[1\] _1369_
+ _1350_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[1\] _1371_ _1348_
+ sg13g2_a221oi_1
X_2947_ _0448_ _0361_ _0437_ VPWR VGND sg13g2_nand2b_1
X_2878_ VGND VPWR net748 _0343_ _0381_ _0379_ sg13g2_a21oi_1
XFILLER_18_508 VPWR VGND sg13g2_decap_8
XFILLER_46_839 VPWR VGND sg13g2_decap_8
XFILLER_26_530 VPWR VGND sg13g2_decap_8
XFILLER_41_544 VPWR VGND sg13g2_decap_8
XFILLER_14_758 VPWR VGND sg13g2_decap_8
XFILLER_6_946 VPWR VGND sg13g2_decap_8
XFILLER_10_975 VPWR VGND sg13g2_decap_8
XFILLER_5_478 VPWR VGND sg13g2_decap_8
XFILLER_49_622 VPWR VGND sg13g2_decap_8
XFILLER_1_695 VPWR VGND sg13g2_decap_8
XFILLER_23_1026 VPWR VGND sg13g2_fill_2
XFILLER_37_817 VPWR VGND sg13g2_decap_8
XFILLER_49_699 VPWR VGND sg13g2_decap_8
XFILLER_45_883 VPWR VGND sg13g2_decap_8
XFILLER_17_541 VPWR VGND sg13g2_decap_8
XFILLER_44_393 VPWR VGND sg13g2_decap_4
XFILLER_44_382 VPWR VGND sg13g2_fill_1
XFILLER_44_371 VPWR VGND sg13g2_fill_2
XFILLER_32_511 VPWR VGND sg13g2_decap_8
X_3850_ _0758_ _0929_ _1254_ _1255_ VPWR VGND sg13g2_nor3_1
X_2801_ _1665_ VPWR _0315_ VGND _0309_ _0314_ sg13g2_o21ai_1
XFILLER_20_728 VPWR VGND sg13g2_decap_8
X_3781_ _1057_ _1058_ net580 _1212_ VPWR VGND sg13g2_nor3_1
XFILLER_32_588 VPWR VGND sg13g2_decap_8
X_2732_ net577 VPWR _0262_ VGND _0257_ _0261_ sg13g2_o21ai_1
XFILLER_30_1008 VPWR VGND sg13g2_decap_8
XFILLER_9_795 VPWR VGND sg13g2_decap_8
X_2663_ _0197_ net614 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[3\]
+ net622 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[3\] VPWR VGND sg13g2_a22oi_1
X_2594_ _2003_ _1916_ _2002_ VPWR VGND sg13g2_nand2_1
X_4333_ net835 VGND VPWR _0190_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[1\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_2
XFILLER_5_61 VPWR VGND sg13g2_fill_2
X_4264_ net813 VGND VPWR _0121_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[7\]
+ clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3215_ net714 _0681_ _0683_ _0685_ _0686_ VPWR VGND sg13g2_nor4_1
X_4195_ net824 VGND VPWR _0052_ sap_3_inst.alu_inst.tmp\[2\] clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
XFILLER_28_806 VPWR VGND sg13g2_decap_8
X_3146_ _0623_ net718 net19 VPWR VGND sg13g2_nand2_1
X_3077_ VGND VPWR _0542_ _0554_ _0574_ _0540_ sg13g2_a21oi_1
XFILLER_23_522 VPWR VGND sg13g2_decap_8
XFILLER_36_883 VPWR VGND sg13g2_decap_8
XFILLER_23_599 VPWR VGND sg13g2_decap_8
X_3979_ _1355_ _1349_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[0\]
+ _1347_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_3_938 VPWR VGND sg13g2_decap_8
Xfanout730 _1582_ net730 VPWR VGND sg13g2_buf_8
Xfanout741 _1566_ net741 VPWR VGND sg13g2_buf_8
Xfanout752 _1558_ net752 VPWR VGND sg13g2_buf_8
Xfanout763 sap_3_inst.controller_inst.opcode\[3\] net763 VPWR VGND sg13g2_buf_8
Xfanout774 sap_3_inst.alu_inst.acc\[7\] net774 VPWR VGND sg13g2_buf_8
Xfanout785 sap_3_inst.alu_inst.acc\[3\] net785 VPWR VGND sg13g2_buf_8
XFILLER_18_305 VPWR VGND sg13g2_fill_2
Xfanout796 _1338_ net796 VPWR VGND sg13g2_buf_8
XFILLER_46_636 VPWR VGND sg13g2_decap_8
XFILLER_27_861 VPWR VGND sg13g2_decap_8
XFILLER_42_842 VPWR VGND sg13g2_decap_8
XFILLER_14_555 VPWR VGND sg13g2_decap_8
XFILLER_10_772 VPWR VGND sg13g2_decap_8
XFILLER_6_743 VPWR VGND sg13g2_decap_8
XFILLER_2_960 VPWR VGND sg13g2_decap_8
XFILLER_1_492 VPWR VGND sg13g2_decap_8
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
X_3000_ VPWR VGND _0499_ net599 _0498_ _1991_ _0500_ _0330_ sg13g2_a221oi_1
XFILLER_37_614 VPWR VGND sg13g2_decap_8
XFILLER_49_496 VPWR VGND sg13g2_decap_8
XFILLER_18_872 VPWR VGND sg13g2_decap_8
XFILLER_45_680 VPWR VGND sg13g2_decap_8
XFILLER_33_820 VPWR VGND sg13g2_decap_8
X_3902_ VGND VPWR _1512_ net643 _0147_ _1291_ sg13g2_a21oi_1
X_3833_ _0128_ _1238_ _1241_ VPWR VGND sg13g2_nand2_1
XFILLER_33_897 VPWR VGND sg13g2_decap_8
XFILLER_20_525 VPWR VGND sg13g2_decap_8
X_3764_ _1192_ VPWR _0103_ VGND _1007_ _1197_ sg13g2_o21ai_1
XFILLER_9_592 VPWR VGND sg13g2_decap_8
X_3695_ VPWR VGND _0306_ _0732_ net604 _1914_ _1143_ net668 sg13g2_a221oi_1
X_2715_ _0245_ net619 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[0\]
+ net620 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[0\] VPWR VGND
+ sg13g2_a22oi_1
X_2646_ _2053_ VPWR _0028_ VGND _1487_ _2024_ sg13g2_o21ai_1
X_2577_ _1988_ net601 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[4\]
+ net711 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[4\] VPWR VGND
+ sg13g2_a22oi_1
X_4316_ net815 VGND VPWR _0173_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[4\]
+ clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4247_ net812 VGND VPWR _0104_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[6\]
+ clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4178_ net824 VGND VPWR _0035_ sap_3_inst.alu_inst.acc\[2\] clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_28_603 VPWR VGND sg13g2_decap_8
X_3129_ net17 sap_3_inst.alu_inst.tmp\[0\] net701 _0050_ VPWR VGND sg13g2_mux2_1
XFILLER_36_680 VPWR VGND sg13g2_decap_8
XFILLER_24_864 VPWR VGND sg13g2_decap_8
XFILLER_11_558 VPWR VGND sg13g2_decap_8
XFILLER_3_735 VPWR VGND sg13g2_decap_8
Xfanout582 _1146_ net582 VPWR VGND sg13g2_buf_8
Xfanout593 net594 net593 VPWR VGND sg13g2_buf_2
Xfanout571 net572 net571 VPWR VGND sg13g2_buf_8
XFILLER_47_956 VPWR VGND sg13g2_decap_8
XFILLER_46_433 VPWR VGND sg13g2_decap_8
XFILLER_19_658 VPWR VGND sg13g2_decap_8
XFILLER_18_135 VPWR VGND sg13g2_fill_2
XFILLER_33_127 VPWR VGND sg13g2_fill_1
XFILLER_15_875 VPWR VGND sg13g2_decap_8
XFILLER_30_812 VPWR VGND sg13g2_decap_8
XFILLER_30_889 VPWR VGND sg13g2_decap_8
XFILLER_6_540 VPWR VGND sg13g2_decap_8
X_2500_ _1627_ net722 _1557_ _1916_ VPWR VGND sg13g2_nand3_1
X_3480_ VGND VPWR net665 _0945_ _0948_ _0947_ sg13g2_a21oi_1
X_2431_ _1848_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[7\] net628
+ VPWR VGND sg13g2_nand2_1
X_2362_ VGND VPWR _1693_ net721 _1779_ _1656_ sg13g2_a21oi_1
X_2293_ _1660_ _1709_ _1710_ VPWR VGND sg13g2_nor2_1
X_4101_ _1456_ VPWR _0181_ VGND net578 _1455_ sg13g2_o21ai_1
X_4032_ _1403_ _1351_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[5\]
+ _1350_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_38_923 VPWR VGND sg13g2_decap_8
XFILLER_49_293 VPWR VGND sg13g2_decap_8
XFILLER_49_271 VPWR VGND sg13g2_fill_2
XFILLER_25_639 VPWR VGND sg13g2_decap_8
XFILLER_37_488 VPWR VGND sg13g2_decap_8
XFILLER_24_127 VPWR VGND sg13g2_fill_2
XFILLER_33_694 VPWR VGND sg13g2_decap_8
XFILLER_21_867 VPWR VGND sg13g2_decap_8
X_3816_ net680 VPWR _1232_ VGND net586 _1045_ sg13g2_o21ai_1
X_3747_ VGND VPWR _1183_ _0945_ net588 sg13g2_or2_1
X_3678_ _1127_ VPWR _1128_ VGND net569 net604 sg13g2_o21ai_1
X_2629_ _2038_ net748 _1902_ VPWR VGND sg13g2_nand2_1
Xclkbuf_4_14_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs
+ clknet_4_14_0_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_43_1018 VPWR VGND sg13g2_decap_8
XFILLER_0_749 VPWR VGND sg13g2_decap_8
XFILLER_29_901 VPWR VGND sg13g2_decap_8
XFILLER_44_904 VPWR VGND sg13g2_decap_8
XFILLER_29_978 VPWR VGND sg13g2_decap_8
XFILLER_16_639 VPWR VGND sg13g2_decap_8
XFILLER_28_477 VPWR VGND sg13g2_decap_8
XFILLER_43_458 VPWR VGND sg13g2_decap_8
XFILLER_24_661 VPWR VGND sg13g2_decap_8
XFILLER_12_856 VPWR VGND sg13g2_decap_8
XFILLER_23_160 VPWR VGND sg13g2_fill_1
XFILLER_7_337 VPWR VGND sg13g2_fill_1
XFILLER_3_532 VPWR VGND sg13g2_decap_8
XFILLER_11_93 VPWR VGND sg13g2_fill_2
XFILLER_4_1012 VPWR VGND sg13g2_decap_8
XFILLER_47_753 VPWR VGND sg13g2_decap_8
XFILLER_35_904 VPWR VGND sg13g2_decap_8
XFILLER_36_90 VPWR VGND sg13g2_fill_2
X_2980_ VPWR _0480_ _0479_ VGND sg13g2_inv_1
XFILLER_15_672 VPWR VGND sg13g2_decap_8
XFILLER_21_119 VPWR VGND sg13g2_fill_2
X_3601_ _1062_ _2051_ _1063_ VPWR VGND sg13g2_nor2b_2
XFILLER_30_686 VPWR VGND sg13g2_decap_8
X_3532_ net14 net605 _0998_ VPWR VGND sg13g2_nor2_1
X_3463_ _0742_ VPWR _0932_ VGND net587 _0928_ sg13g2_o21ai_1
X_2414_ _1553_ _1610_ sap_3_inst.controller_inst.opcode\[0\] _1831_ VPWR VGND _1617_
+ sg13g2_nand4_1
X_3394_ _0771_ _0779_ _0786_ _0865_ VGND VPWR _0863_ sg13g2_nor4_2
X_2345_ net760 net757 net763 _1762_ VPWR VGND sg13g2_nand3_1
X_2276_ _1693_ _1553_ _1671_ VPWR VGND sg13g2_nand2_2
XFILLER_38_720 VPWR VGND sg13g2_decap_8
Xclkbuf_1_0__f_sap_3_inst.alu_inst.clk clknet_0_sap_3_inst.alu_inst.clk clknet_1_0__leaf_sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_8
XFILLER_26_915 VPWR VGND sg13g2_decap_8
X_4015_ _1388_ _1350_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[3\]
+ _1349_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_38_797 VPWR VGND sg13g2_decap_8
XFILLER_25_436 VPWR VGND sg13g2_decap_8
XFILLER_41_929 VPWR VGND sg13g2_decap_8
XFILLER_33_480 VPWR VGND sg13g2_fill_2
XFILLER_33_491 VPWR VGND sg13g2_decap_8
XFILLER_21_664 VPWR VGND sg13g2_decap_8
XFILLER_10_1017 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_528 VPWR VGND sg13g2_decap_8
XFILLER_44_701 VPWR VGND sg13g2_decap_8
XFILLER_17_926 VPWR VGND sg13g2_decap_8
XFILLER_29_775 VPWR VGND sg13g2_decap_8
XFILLER_44_778 VPWR VGND sg13g2_decap_8
XFILLER_31_417 VPWR VGND sg13g2_fill_1
XFILLER_40_940 VPWR VGND sg13g2_decap_8
XFILLER_12_653 VPWR VGND sg13g2_decap_8
XFILLER_7_123 VPWR VGND sg13g2_fill_2
XFILLER_8_668 VPWR VGND sg13g2_decap_8
XFILLER_4_830 VPWR VGND sg13g2_decap_8
XFILLER_26_1013 VPWR VGND sg13g2_decap_8
X_2130_ VPWR _1548_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[7\]
+ VGND sg13g2_inv_1
XFILLER_47_550 VPWR VGND sg13g2_decap_8
XFILLER_35_701 VPWR VGND sg13g2_decap_8
XFILLER_23_907 VPWR VGND sg13g2_decap_8
XFILLER_34_222 VPWR VGND sg13g2_fill_1
XFILLER_35_778 VPWR VGND sg13g2_decap_8
X_2963_ _0451_ _0463_ net575 _0464_ VPWR VGND sg13g2_nand3_1
X_2894_ _0390_ _0395_ _0384_ _0397_ VPWR VGND sg13g2_nand3_1
X_3515_ _0959_ VPWR _0070_ VGND _0976_ _0980_ sg13g2_o21ai_1
X_3446_ VPWR _0915_ _0914_ VGND sg13g2_inv_1
X_3377_ _0848_ net589 _0847_ VPWR VGND sg13g2_nand2_2
X_2328_ _1745_ _1649_ _1744_ VPWR VGND sg13g2_nand2_1
X_2259_ net731 _1672_ _1676_ VPWR VGND sg13g2_nor2_1
XFILLER_26_712 VPWR VGND sg13g2_decap_8
XFILLER_38_594 VPWR VGND sg13g2_decap_8
XFILLER_26_789 VPWR VGND sg13g2_decap_8
XFILLER_41_726 VPWR VGND sg13g2_decap_8
XFILLER_22_984 VPWR VGND sg13g2_decap_8
XFILLER_1_800 VPWR VGND sg13g2_decap_8
XFILLER_49_804 VPWR VGND sg13g2_decap_8
XFILLER_1_877 VPWR VGND sg13g2_decap_8
XFILLER_48_325 VPWR VGND sg13g2_decap_8
XFILLER_17_723 VPWR VGND sg13g2_decap_8
XFILLER_29_572 VPWR VGND sg13g2_decap_8
XFILLER_44_575 VPWR VGND sg13g2_decap_8
XFILLER_31_214 VPWR VGND sg13g2_fill_1
XFILLER_9_900 VPWR VGND sg13g2_decap_8
XFILLER_12_450 VPWR VGND sg13g2_fill_2
XFILLER_13_984 VPWR VGND sg13g2_decap_8
XFILLER_9_977 VPWR VGND sg13g2_decap_8
X_3300_ _0771_ _0768_ _0769_ VPWR VGND sg13g2_nand2_1
X_4280_ net809 VGND VPWR _0137_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[7\]
+ clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3231_ _1633_ _0659_ _0701_ _0702_ VPWR VGND sg13g2_nor3_1
X_3162_ VGND VPWR _1634_ _1709_ _0633_ _1653_ sg13g2_a21oi_1
X_2113_ VPWR _1531_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[4\]
+ VGND sg13g2_inv_1
X_3093_ _0585_ _0587_ net575 _0590_ VPWR VGND _0589_ sg13g2_nand4_1
XFILLER_48_892 VPWR VGND sg13g2_decap_8
XFILLER_23_704 VPWR VGND sg13g2_decap_8
XFILLER_35_575 VPWR VGND sg13g2_decap_8
X_3995_ _1370_ _1353_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[1\]
+ _1347_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2946_ _0446_ VPWR _0447_ VGND _0355_ _0439_ sg13g2_o21ai_1
X_2877_ _0380_ net748 _0343_ _0379_ VPWR VGND sg13g2_and3_2
X_3429_ VGND VPWR _0770_ _0868_ _0899_ _0891_ sg13g2_a21oi_1
XFILLER_46_818 VPWR VGND sg13g2_decap_8
XFILLER_41_523 VPWR VGND sg13g2_decap_8
XFILLER_14_737 VPWR VGND sg13g2_decap_8
XFILLER_26_586 VPWR VGND sg13g2_decap_8
XFILLER_22_781 VPWR VGND sg13g2_decap_8
XFILLER_10_954 VPWR VGND sg13g2_decap_8
XFILLER_6_925 VPWR VGND sg13g2_decap_8
XFILLER_5_402 VPWR VGND sg13g2_fill_2
XFILLER_5_457 VPWR VGND sg13g2_decap_8
XFILLER_49_601 VPWR VGND sg13g2_decap_8
XFILLER_1_674 VPWR VGND sg13g2_decap_8
XFILLER_23_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_678 VPWR VGND sg13g2_decap_8
XFILLER_17_520 VPWR VGND sg13g2_decap_8
XFILLER_45_862 VPWR VGND sg13g2_decap_8
XFILLER_17_597 VPWR VGND sg13g2_decap_8
XFILLER_20_707 VPWR VGND sg13g2_decap_8
XFILLER_32_567 VPWR VGND sg13g2_decap_8
X_2800_ _0314_ _0312_ _0313_ VPWR VGND sg13g2_nand2_1
X_3780_ net683 net602 _1211_ VPWR VGND sg13g2_nor2_1
XFILLER_13_781 VPWR VGND sg13g2_decap_8
X_2731_ _0259_ _0260_ _0258_ _0261_ VPWR VGND sg13g2_nand3_1
XFILLER_9_774 VPWR VGND sg13g2_decap_8
X_2662_ VGND VPWR _0196_ _2068_ _1768_ sg13g2_or2_1
X_2593_ _1996_ net704 _2001_ _2002_ VPWR VGND sg13g2_nor3_2
X_4332_ net835 VGND VPWR _0189_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[0\]
+ clknet_3_6__leaf_clk sg13g2_dfrbpq_2
X_4263_ net811 VGND VPWR _0120_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[6\]
+ clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3214_ _0684_ VPWR _0685_ VGND _1660_ _1752_ sg13g2_o21ai_1
X_4194_ net820 VGND VPWR _0051_ sap_3_inst.alu_inst.tmp\[1\] clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
X_3145_ VGND VPWR net717 _2051_ _0059_ _0622_ sg13g2_a21oi_1
X_3076_ VPWR _0573_ _0572_ VGND sg13g2_inv_1
XFILLER_39_199 VPWR VGND sg13g2_fill_2
XFILLER_39_1012 VPWR VGND sg13g2_decap_8
XFILLER_36_862 VPWR VGND sg13g2_decap_8
XFILLER_23_501 VPWR VGND sg13g2_decap_8
XFILLER_23_578 VPWR VGND sg13g2_decap_8
X_3978_ _1354_ _1352_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[0\]
+ net797 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2929_ net575 _0417_ _0431_ VPWR VGND sg13g2_nor2_1
XFILLER_3_917 VPWR VGND sg13g2_decap_8
XFILLER_49_57 VPWR VGND sg13g2_fill_2
Xfanout720 _1752_ net720 VPWR VGND sg13g2_buf_8
Xfanout742 _1566_ net742 VPWR VGND sg13g2_buf_1
Xfanout731 _1582_ net731 VPWR VGND sg13g2_buf_8
Xfanout775 net776 net775 VPWR VGND sg13g2_buf_8
Xfanout753 net754 net753 VPWR VGND sg13g2_buf_8
Xfanout764 sap_3_inst.controller_inst.opcode\[3\] net764 VPWR VGND sg13g2_buf_8
XFILLER_46_615 VPWR VGND sg13g2_decap_8
Xfanout786 net788 net786 VPWR VGND sg13g2_buf_8
Xfanout797 _1337_ net797 VPWR VGND sg13g2_buf_8
XFILLER_27_840 VPWR VGND sg13g2_decap_8
XFILLER_42_821 VPWR VGND sg13g2_decap_8
XFILLER_14_534 VPWR VGND sg13g2_decap_8
XFILLER_42_898 VPWR VGND sg13g2_decap_8
XFILLER_10_751 VPWR VGND sg13g2_decap_8
XFILLER_6_722 VPWR VGND sg13g2_decap_8
XFILLER_5_254 VPWR VGND sg13g2_fill_1
XFILLER_6_799 VPWR VGND sg13g2_decap_8
XFILLER_7_1010 VPWR VGND sg13g2_decap_8
XFILLER_1_471 VPWR VGND sg13g2_decap_8
XFILLER_49_475 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
XFILLER_18_851 VPWR VGND sg13g2_decap_8
XFILLER_24_309 VPWR VGND sg13g2_fill_1
X_3901_ VPWR VGND _1290_ net643 _1103_ net607 _1291_ _0901_ sg13g2_a221oi_1
XFILLER_32_320 VPWR VGND sg13g2_fill_2
X_3832_ _1240_ VPWR _1241_ VGND _1084_ _1140_ sg13g2_o21ai_1
XFILLER_20_504 VPWR VGND sg13g2_decap_8
XFILLER_33_876 VPWR VGND sg13g2_decap_8
XFILLER_9_571 VPWR VGND sg13g2_decap_8
X_3763_ net675 VPWR _1197_ VGND _1194_ _1196_ sg13g2_o21ai_1
X_2714_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[0\] net630
+ net629 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[0\] _0244_ net712
+ sg13g2_a221oi_1
X_3694_ net612 _1041_ _1142_ VPWR VGND sg13g2_nor2_1
X_2645_ _2051_ net710 _2052_ _2053_ VPWR VGND sg13g2_a21o_1
X_2576_ _1987_ net618 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[4\]
+ net631 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4315_ net831 VGND VPWR _0172_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[3\]
+ clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4246_ net814 VGND VPWR _0103_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[5\]
+ clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4177_ net820 VGND VPWR _0034_ sap_3_inst.alu_inst.acc\[1\] clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3128_ _1880_ VPWR _0615_ VGND _1800_ _0614_ sg13g2_o21ai_1
XFILLER_28_659 VPWR VGND sg13g2_decap_8
X_3059_ _0557_ _0520_ _0555_ VPWR VGND sg13g2_nand2_1
XFILLER_42_128 VPWR VGND sg13g2_fill_2
XFILLER_24_843 VPWR VGND sg13g2_decap_8
XFILLER_11_537 VPWR VGND sg13g2_decap_8
XFILLER_13_1026 VPWR VGND sg13g2_fill_2
XFILLER_3_714 VPWR VGND sg13g2_decap_8
Xclkbuf_5_23__f_sap_3_inst.alu_inst.clk_regs clknet_4_11_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
Xfanout583 _1053_ net583 VPWR VGND sg13g2_buf_8
Xfanout572 _0943_ net572 VPWR VGND sg13g2_buf_1
XFILLER_47_935 VPWR VGND sg13g2_decap_8
XFILLER_46_412 VPWR VGND sg13g2_decap_8
XFILLER_19_637 VPWR VGND sg13g2_decap_8
XFILLER_20_1008 VPWR VGND sg13g2_decap_8
Xfanout594 net595 net594 VPWR VGND sg13g2_buf_8
XFILLER_46_489 VPWR VGND sg13g2_decap_8
XFILLER_15_854 VPWR VGND sg13g2_decap_8
XFILLER_42_695 VPWR VGND sg13g2_decap_8
XFILLER_30_868 VPWR VGND sg13g2_decap_8
Xclkbuf_5_12__f_sap_3_inst.alu_inst.clk_regs clknet_4_6_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_6_596 VPWR VGND sg13g2_decap_8
X_2430_ net667 net666 net707 _1843_ _1847_ VPWR VGND sg13g2_and4_1
X_2361_ _1653_ _1682_ _1778_ VPWR VGND sg13g2_nor2_1
XFILLER_37_4 VPWR VGND sg13g2_fill_1
X_2292_ _1709_ _1679_ _1553_ net732 net738 VPWR VGND sg13g2_a22oi_1
X_4100_ _1456_ sap_3_inst.alu_inst.act\[4\] net578 VPWR VGND sg13g2_nand2_1
XFILLER_49_250 VPWR VGND sg13g2_decap_8
XFILLER_38_902 VPWR VGND sg13g2_decap_8
X_4031_ net798 net63 _1402_ _0165_ VPWR VGND sg13g2_a21o_1
XFILLER_2_63 VPWR VGND sg13g2_fill_1
XFILLER_38_979 VPWR VGND sg13g2_decap_8
XFILLER_25_618 VPWR VGND sg13g2_decap_8
XFILLER_33_673 VPWR VGND sg13g2_decap_8
XFILLER_21_846 VPWR VGND sg13g2_decap_8
X_3815_ _1231_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[7\] net657
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_367 VPWR VGND sg13g2_fill_1
X_3746_ _1182_ net595 _0951_ VPWR VGND sg13g2_nand2b_1
X_3677_ _1127_ net14 net604 VPWR VGND sg13g2_nand2_1
X_2628_ net791 net695 _2037_ VPWR VGND sg13g2_nor2_1
X_2559_ _1970_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[4\] net622
+ VPWR VGND sg13g2_nand2_1
XFILLER_0_728 VPWR VGND sg13g2_decap_8
X_4229_ net810 VGND VPWR _0086_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[4\]
+ clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_46_25 VPWR VGND sg13g2_fill_1
XFILLER_29_957 VPWR VGND sg13g2_decap_8
XFILLER_28_456 VPWR VGND sg13g2_decap_8
XFILLER_15_117 VPWR VGND sg13g2_fill_1
XFILLER_16_618 VPWR VGND sg13g2_decap_8
XFILLER_24_640 VPWR VGND sg13g2_decap_8
XFILLER_30_109 VPWR VGND sg13g2_fill_2
XFILLER_12_835 VPWR VGND sg13g2_decap_8
XFILLER_11_345 VPWR VGND sg13g2_fill_2
XFILLER_11_356 VPWR VGND sg13g2_fill_1
XFILLER_3_511 VPWR VGND sg13g2_decap_8
XFILLER_3_588 VPWR VGND sg13g2_decap_8
XFILLER_47_732 VPWR VGND sg13g2_decap_8
XFILLER_15_651 VPWR VGND sg13g2_decap_8
XFILLER_42_492 VPWR VGND sg13g2_decap_8
XFILLER_30_665 VPWR VGND sg13g2_decap_8
X_3600_ VGND VPWR _0848_ _0882_ _1062_ net612 sg13g2_a21oi_1
X_3531_ VGND VPWR net663 _0993_ _0997_ _0996_ sg13g2_a21oi_1
X_3462_ _0931_ _0836_ _0882_ VPWR VGND sg13g2_xnor2_1
X_2413_ VPWR VGND net739 net741 _1829_ net743 _1830_ _1581_ sg13g2_a221oi_1
X_3393_ VGND VPWR _0864_ _0863_ _0786_ sg13g2_or2_1
X_2344_ _1493_ net752 _1761_ VPWR VGND sg13g2_nor2_1
XFILLER_28_0 VPWR VGND sg13g2_fill_1
X_2275_ _1553_ net732 _1692_ VPWR VGND sg13g2_and2_1
X_4014_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[3\] _1351_
+ _1387_ net795 sg13g2_a21oi_1
XFILLER_37_242 VPWR VGND sg13g2_fill_2
XFILLER_25_415 VPWR VGND sg13g2_decap_8
XFILLER_38_776 VPWR VGND sg13g2_decap_8
XFILLER_41_908 VPWR VGND sg13g2_decap_8
XFILLER_20_120 VPWR VGND sg13g2_fill_1
XFILLER_21_643 VPWR VGND sg13g2_decap_8
XFILLER_20_164 VPWR VGND sg13g2_fill_1
X_3729_ _1166_ _1167_ _1094_ _1168_ VPWR VGND sg13g2_nand3_1
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_48_507 VPWR VGND sg13g2_decap_8
XFILLER_17_905 VPWR VGND sg13g2_decap_8
XFILLER_29_754 VPWR VGND sg13g2_decap_8
XFILLER_28_253 VPWR VGND sg13g2_fill_1
XFILLER_44_757 VPWR VGND sg13g2_decap_8
XFILLER_43_212 VPWR VGND sg13g2_fill_2
Xclkbuf_4_7_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_7_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_25_982 VPWR VGND sg13g2_decap_8
XFILLER_12_632 VPWR VGND sg13g2_decap_8
XFILLER_40_996 VPWR VGND sg13g2_decap_8
XFILLER_8_647 VPWR VGND sg13g2_decap_8
XFILLER_4_886 VPWR VGND sg13g2_decap_8
XFILLER_39_529 VPWR VGND sg13g2_decap_8
XFILLER_35_757 VPWR VGND sg13g2_decap_8
X_2962_ VGND VPWR _0444_ _0452_ _0463_ _0462_ sg13g2_a21oi_1
XFILLER_16_982 VPWR VGND sg13g2_decap_8
XFILLER_8_40 VPWR VGND sg13g2_fill_1
X_2893_ _0355_ _0374_ _0396_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_985 VPWR VGND sg13g2_decap_8
XFILLER_8_73 VPWR VGND sg13g2_fill_1
X_3514_ _0802_ VPWR _0981_ VGND net591 _0861_ sg13g2_o21ai_1
X_3445_ _0913_ VPWR _0914_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[2\]
+ net662 sg13g2_o21ai_1
X_3376_ _0841_ _0846_ _0847_ VPWR VGND sg13g2_and2_1
X_2327_ _1744_ net730 VPWR VGND _1669_ sg13g2_nand2b_2
X_2258_ VGND VPWR _1670_ _1674_ _1675_ _1666_ sg13g2_a21oi_1
XFILLER_38_573 VPWR VGND sg13g2_decap_8
X_2189_ net728 _1605_ _1606_ VPWR VGND sg13g2_nor2_1
XFILLER_41_705 VPWR VGND sg13g2_decap_8
XFILLER_14_919 VPWR VGND sg13g2_decap_8
XFILLER_26_768 VPWR VGND sg13g2_decap_8
XFILLER_22_963 VPWR VGND sg13g2_decap_8
XFILLER_5_639 VPWR VGND sg13g2_decap_8
XFILLER_49_1014 VPWR VGND sg13g2_decap_8
XFILLER_1_856 VPWR VGND sg13g2_decap_8
XFILLER_48_304 VPWR VGND sg13g2_decap_8
XFILLER_17_702 VPWR VGND sg13g2_decap_8
XFILLER_29_551 VPWR VGND sg13g2_decap_8
XFILLER_44_554 VPWR VGND sg13g2_decap_8
XFILLER_17_779 VPWR VGND sg13g2_decap_8
XFILLER_32_749 VPWR VGND sg13g2_decap_8
XFILLER_13_963 VPWR VGND sg13g2_decap_8
XFILLER_40_793 VPWR VGND sg13g2_decap_8
XFILLER_9_956 VPWR VGND sg13g2_decap_8
XFILLER_4_683 VPWR VGND sg13g2_decap_8
X_3230_ VGND VPWR _1491_ _1493_ _0701_ _1683_ sg13g2_a21oi_1
X_3161_ _0630_ _0631_ _0629_ _0632_ VPWR VGND sg13g2_nand3_1
X_2112_ VPWR _1530_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[4\]
+ VGND sg13g2_inv_1
XFILLER_48_871 VPWR VGND sg13g2_decap_8
X_3092_ _0589_ _0578_ _0588_ _0576_ _0344_ VPWR VGND sg13g2_a22oi_1
XFILLER_35_554 VPWR VGND sg13g2_decap_8
X_3994_ _1366_ _1367_ _1365_ _1369_ VPWR VGND _1368_ sg13g2_nand4_1
X_2945_ sap_3_inst.alu_inst.tmp\[3\] _0363_ net784 _0446_ VPWR VGND sg13g2_nand3_1
X_2876_ _0379_ _0374_ _0378_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_782 VPWR VGND sg13g2_decap_8
X_3428_ net589 _0897_ _0898_ VPWR VGND sg13g2_nor2_1
X_3359_ _0826_ _0827_ _0828_ _0829_ _0830_ VPWR VGND sg13g2_and4_1
XFILLER_45_307 VPWR VGND sg13g2_fill_2
XFILLER_39_893 VPWR VGND sg13g2_decap_8
XFILLER_26_565 VPWR VGND sg13g2_decap_8
XFILLER_41_502 VPWR VGND sg13g2_decap_8
XFILLER_14_716 VPWR VGND sg13g2_decap_8
XFILLER_41_579 VPWR VGND sg13g2_decap_8
XFILLER_16_1024 VPWR VGND sg13g2_decap_4
XFILLER_22_760 VPWR VGND sg13g2_decap_8
XFILLER_10_933 VPWR VGND sg13g2_decap_8
XFILLER_6_904 VPWR VGND sg13g2_decap_8
XFILLER_1_653 VPWR VGND sg13g2_decap_8
XFILLER_48_101 VPWR VGND sg13g2_fill_1
XFILLER_0_163 VPWR VGND sg13g2_fill_1
XFILLER_49_657 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_45_841 VPWR VGND sg13g2_decap_8
XFILLER_17_576 VPWR VGND sg13g2_decap_8
XFILLER_32_546 VPWR VGND sg13g2_decap_8
XFILLER_13_760 VPWR VGND sg13g2_decap_8
XFILLER_40_590 VPWR VGND sg13g2_decap_8
XFILLER_9_753 VPWR VGND sg13g2_decap_8
X_2730_ _0260_ net615 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[0\]
+ net617 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2661_ _2059_ VPWR _2068_ VGND _2063_ _2067_ sg13g2_o21ai_1
X_2592_ VGND VPWR net725 _1673_ _2001_ net733 sg13g2_a21oi_1
XFILLER_5_41 VPWR VGND sg13g2_fill_1
X_4331_ net817 VGND VPWR net65 sap_3_outputReg_start_sync clknet_3_0__leaf_clk sg13g2_dfrbpq_1
X_4262_ net815 VGND VPWR _0119_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[5\]
+ clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_5_96 VPWR VGND sg13g2_fill_2
XFILLER_5_74 VPWR VGND sg13g2_fill_1
XFILLER_4_480 VPWR VGND sg13g2_decap_8
X_3213_ _1645_ VPWR _0684_ VGND _1612_ _1672_ sg13g2_o21ai_1
XFILLER_39_101 VPWR VGND sg13g2_fill_2
X_4149__7 VPWR net41 clknet_leaf_2_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
X_4193_ net820 VGND VPWR _0050_ sap_3_inst.alu_inst.tmp\[0\] clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
X_3144_ net769 net718 _0622_ VPWR VGND sg13g2_nor2_1
XFILLER_39_145 VPWR VGND sg13g2_fill_2
X_3075_ _0572_ _0571_ VPWR VGND _0570_ sg13g2_nand2b_2
XFILLER_36_841 VPWR VGND sg13g2_decap_8
XFILLER_23_557 VPWR VGND sg13g2_decap_8
X_3977_ _1336_ _1341_ _1353_ VPWR VGND sg13g2_nor2_2
XFILLER_11_719 VPWR VGND sg13g2_decap_8
X_2928_ VGND VPWR _0412_ _0428_ _0430_ _0429_ sg13g2_a21oi_1
X_2859_ net761 _2013_ _2017_ _0363_ VPWR VGND sg13g2_nor3_2
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_8 VPWR VGND sg13g2_fill_2
Xfanout732 _1671_ net732 VPWR VGND sg13g2_buf_8
Xfanout721 _1723_ net721 VPWR VGND sg13g2_buf_8
Xfanout710 _1915_ net710 VPWR VGND sg13g2_buf_8
Xfanout765 sap_3_inst.controller_inst.opcode\[2\] net765 VPWR VGND sg13g2_buf_8
Xfanout776 net777 net776 VPWR VGND sg13g2_buf_8
Xfanout743 _1551_ net743 VPWR VGND sg13g2_buf_8
Xfanout754 sap_3_inst.controller_inst.opcode\[7\] net754 VPWR VGND sg13g2_buf_8
Xfanout787 net788 net787 VPWR VGND sg13g2_buf_1
XFILLER_19_819 VPWR VGND sg13g2_decap_8
Xfanout798 _1313_ net798 VPWR VGND sg13g2_buf_8
XFILLER_39_690 VPWR VGND sg13g2_decap_8
XFILLER_45_148 VPWR VGND sg13g2_fill_1
XFILLER_42_800 VPWR VGND sg13g2_decap_8
XFILLER_14_513 VPWR VGND sg13g2_decap_8
XFILLER_27_896 VPWR VGND sg13g2_decap_8
XFILLER_42_877 VPWR VGND sg13g2_decap_8
XFILLER_10_730 VPWR VGND sg13g2_decap_8
XFILLER_6_701 VPWR VGND sg13g2_decap_8
XFILLER_14_94 VPWR VGND sg13g2_fill_1
XFILLER_6_778 VPWR VGND sg13g2_decap_8
Xclkbuf_4_15_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs
+ clknet_4_15_0_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_2_995 VPWR VGND sg13g2_decap_8
XFILLER_1_450 VPWR VGND sg13g2_decap_8
XFILLER_49_454 VPWR VGND sg13g2_decap_8
XFILLER_18_830 VPWR VGND sg13g2_decap_8
XFILLER_37_649 VPWR VGND sg13g2_decap_8
XFILLER_17_373 VPWR VGND sg13g2_fill_2
X_3900_ net612 VPWR _1290_ VGND _0302_ _1289_ sg13g2_o21ai_1
XFILLER_33_855 VPWR VGND sg13g2_decap_8
X_3831_ VGND VPWR net610 _1239_ _1240_ net634 sg13g2_a21oi_1
X_3762_ _1196_ _1195_ _1002_ VPWR VGND sg13g2_nand2b_1
XFILLER_9_550 VPWR VGND sg13g2_decap_8
X_3693_ _1131_ VPWR _0088_ VGND _1133_ _1141_ sg13g2_o21ai_1
X_2713_ _0241_ _0242_ _0240_ _0243_ VPWR VGND sg13g2_nand3_1
X_2644_ _2024_ VPWR _2052_ VGND sap_3_inst.alu_inst.carry net710 sg13g2_o21ai_1
X_2575_ _1986_ net600 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[4\]
+ net622 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4314_ net819 VGND VPWR _0171_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[2\]
+ clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4245_ net810 VGND VPWR _0102_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[4\]
+ clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4176_ net818 VGND VPWR _0033_ sap_3_inst.alu_inst.acc\[0\] clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3127_ _0614_ net716 _0613_ VPWR VGND sg13g2_nand2_1
XFILLER_28_638 VPWR VGND sg13g2_decap_8
XFILLER_43_619 VPWR VGND sg13g2_decap_8
X_3058_ _0556_ _0542_ _0554_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_822 VPWR VGND sg13g2_decap_8
XFILLER_11_516 VPWR VGND sg13g2_decap_8
XFILLER_24_899 VPWR VGND sg13g2_decap_8
XFILLER_13_1005 VPWR VGND sg13g2_decap_8
Xfanout584 _1053_ net584 VPWR VGND sg13g2_buf_1
XFILLER_47_914 VPWR VGND sg13g2_decap_8
Xfanout573 _0967_ net573 VPWR VGND sg13g2_buf_8
XFILLER_19_616 VPWR VGND sg13g2_decap_8
Xfanout595 _0744_ net595 VPWR VGND sg13g2_buf_8
XFILLER_46_468 VPWR VGND sg13g2_decap_8
XFILLER_34_619 VPWR VGND sg13g2_decap_8
XFILLER_15_833 VPWR VGND sg13g2_decap_8
XFILLER_27_693 VPWR VGND sg13g2_decap_8
XFILLER_42_674 VPWR VGND sg13g2_decap_8
XFILLER_30_847 VPWR VGND sg13g2_decap_8
XFILLER_6_575 VPWR VGND sg13g2_decap_8
X_2360_ _1646_ _1691_ _1640_ _1777_ VPWR VGND sg13g2_nand3_1
X_2291_ _1704_ _1707_ _1708_ VPWR VGND sg13g2_nor2_1
XFILLER_2_792 VPWR VGND sg13g2_decap_8
X_4030_ VGND VPWR _1396_ _1400_ _1402_ _1401_ sg13g2_a21oi_1
XFILLER_38_958 VPWR VGND sg13g2_decap_8
XFILLER_24_129 VPWR VGND sg13g2_fill_1
XFILLER_33_652 VPWR VGND sg13g2_decap_8
XFILLER_36_1016 VPWR VGND sg13g2_decap_8
XFILLER_36_1027 VPWR VGND sg13g2_fill_2
XFILLER_21_825 VPWR VGND sg13g2_decap_8
X_3814_ _0120_ _1204_ _1230_ net657 _1543_ VPWR VGND sg13g2_a22oi_1
X_3745_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[3\] net678 _1181_
+ VPWR VGND sg13g2_nor2_1
X_3676_ net638 _0995_ _1126_ VPWR VGND sg13g2_nor2_1
X_2627_ VPWR VGND _2034_ _1768_ _2031_ _1510_ _2036_ net630 sg13g2_a221oi_1
X_2558_ _1969_ net632 sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[4\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_0_707 VPWR VGND sg13g2_decap_8
X_2489_ _1906_ net614 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[7\]
+ net618 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[7\] VPWR VGND
+ sg13g2_a22oi_1
X_4228_ net828 VGND VPWR _0085_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[3\]
+ clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_29_936 VPWR VGND sg13g2_decap_8
X_4159_ net822 VGND VPWR _0020_ u_ser.shadow_reg\[3\] clknet_3_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_939 VPWR VGND sg13g2_decap_8
XFILLER_12_814 VPWR VGND sg13g2_decap_8
XFILLER_24_696 VPWR VGND sg13g2_decap_8
XFILLER_8_829 VPWR VGND sg13g2_decap_8
XFILLER_3_567 VPWR VGND sg13g2_decap_8
XFILLER_11_95 VPWR VGND sg13g2_fill_1
XFILLER_47_711 VPWR VGND sg13g2_decap_8
XFILLER_46_232 VPWR VGND sg13g2_fill_2
XFILLER_47_788 VPWR VGND sg13g2_decap_8
XFILLER_46_276 VPWR VGND sg13g2_decap_8
XFILLER_35_939 VPWR VGND sg13g2_decap_8
XFILLER_15_630 VPWR VGND sg13g2_decap_8
XFILLER_27_490 VPWR VGND sg13g2_decap_8
XFILLER_36_92 VPWR VGND sg13g2_fill_1
XFILLER_43_983 VPWR VGND sg13g2_decap_8
XFILLER_42_471 VPWR VGND sg13g2_decap_8
XFILLER_30_644 VPWR VGND sg13g2_decap_8
X_3530_ net593 VPWR _0996_ VGND net663 _0995_ sg13g2_o21ai_1
XFILLER_11_880 VPWR VGND sg13g2_decap_8
XFILLER_7_884 VPWR VGND sg13g2_decap_8
X_3461_ net591 _0860_ _0930_ VPWR VGND sg13g2_nor2_1
X_2412_ _1617_ net722 net769 _1829_ VPWR VGND sg13g2_nand3_1
X_3392_ _0803_ _0814_ _0794_ _0863_ VPWR VGND _0859_ sg13g2_nand4_1
X_2343_ VGND VPWR _1760_ _1758_ _1592_ sg13g2_or2_1
X_2274_ VGND VPWR _1691_ net749 _1562_ sg13g2_or2_1
X_4013_ _1386_ _1384_ _1385_ VPWR VGND sg13g2_nand2_1
XFILLER_38_755 VPWR VGND sg13g2_decap_8
XFILLER_19_980 VPWR VGND sg13g2_decap_8
XFILLER_21_622 VPWR VGND sg13g2_decap_8
XFILLER_34_983 VPWR VGND sg13g2_decap_8
XFILLER_21_699 VPWR VGND sg13g2_decap_8
X_3728_ VGND VPWR net655 _1055_ _1167_ _1056_ sg13g2_a21oi_1
X_3659_ net637 _0929_ _1109_ _1111_ _1112_ VPWR VGND sg13g2_or4_1
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_29_733 VPWR VGND sg13g2_decap_8
XFILLER_44_736 VPWR VGND sg13g2_decap_8
XFILLER_25_961 VPWR VGND sg13g2_decap_8
XFILLER_12_611 VPWR VGND sg13g2_decap_8
XFILLER_19_1022 VPWR VGND sg13g2_decap_8
XFILLER_24_493 VPWR VGND sg13g2_decap_8
XFILLER_40_975 VPWR VGND sg13g2_decap_8
XFILLER_8_626 VPWR VGND sg13g2_decap_8
XFILLER_12_688 VPWR VGND sg13g2_decap_8
XFILLER_7_125 VPWR VGND sg13g2_fill_1
XFILLER_4_865 VPWR VGND sg13g2_decap_8
XFILLER_3_353 VPWR VGND sg13g2_fill_2
XFILLER_39_508 VPWR VGND sg13g2_decap_8
XFILLER_21_8 VPWR VGND sg13g2_fill_2
XFILLER_19_232 VPWR VGND sg13g2_fill_1
XFILLER_47_585 VPWR VGND sg13g2_decap_8
XFILLER_35_736 VPWR VGND sg13g2_decap_8
XFILLER_16_961 VPWR VGND sg13g2_decap_8
XFILLER_34_246 VPWR VGND sg13g2_fill_2
XFILLER_43_780 VPWR VGND sg13g2_decap_8
X_2961_ _0461_ VPWR _0462_ VGND net783 _0334_ sg13g2_o21ai_1
XFILLER_31_964 VPWR VGND sg13g2_decap_8
X_2892_ _0393_ _0394_ _0344_ _0395_ VPWR VGND sg13g2_nand3_1
XFILLER_30_452 VPWR VGND sg13g2_fill_2
X_3513_ _0742_ VPWR _0980_ VGND net586 _0979_ sg13g2_o21ai_1
XFILLER_7_681 VPWR VGND sg13g2_decap_8
X_3444_ _0910_ _0911_ _0909_ _0913_ VPWR VGND _0912_ sg13g2_nand4_1
X_3375_ _0842_ _0843_ _0844_ _0845_ _0846_ VPWR VGND sg13g2_nor4_1
X_2326_ _1741_ VPWR _1743_ VGND _1696_ _1742_ sg13g2_o21ai_1
X_2257_ _1629_ _1672_ _1674_ VPWR VGND sg13g2_nor2_1
XFILLER_38_552 VPWR VGND sg13g2_decap_8
X_2188_ _1605_ _1561_ _1603_ VPWR VGND sg13g2_nand2_2
XFILLER_26_747 VPWR VGND sg13g2_decap_8
XFILLER_34_780 VPWR VGND sg13g2_decap_8
XFILLER_22_942 VPWR VGND sg13g2_decap_8
XFILLER_21_496 VPWR VGND sg13g2_decap_8
XFILLER_5_618 VPWR VGND sg13g2_decap_8
XFILLER_1_835 VPWR VGND sg13g2_decap_8
XFILLER_49_839 VPWR VGND sg13g2_decap_8
XFILLER_29_530 VPWR VGND sg13g2_decap_8
XFILLER_44_533 VPWR VGND sg13g2_decap_8
XFILLER_1_1017 VPWR VGND sg13g2_decap_8
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_17_758 VPWR VGND sg13g2_decap_8
XFILLER_32_728 VPWR VGND sg13g2_decap_8
XFILLER_13_942 VPWR VGND sg13g2_decap_8
XFILLER_40_772 VPWR VGND sg13g2_decap_8
XFILLER_9_935 VPWR VGND sg13g2_decap_8
XFILLER_12_485 VPWR VGND sg13g2_decap_8
XFILLER_4_662 VPWR VGND sg13g2_decap_8
X_3160_ _0631_ _1635_ net724 VPWR VGND sg13g2_nand2b_1
X_2111_ _1529_ sap_3_inst.alu_inst.tmp\[7\] VPWR VGND sg13g2_inv_2
X_3091_ _0346_ VPWR _0588_ VGND _0349_ _0552_ sg13g2_o21ai_1
Xhold1 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[0\] VPWR VGND net48
+ sg13g2_dlygate4sd3_1
XFILLER_39_349 VPWR VGND sg13g2_fill_1
XFILLER_48_850 VPWR VGND sg13g2_decap_8
XFILLER_47_382 VPWR VGND sg13g2_decap_8
XFILLER_35_533 VPWR VGND sg13g2_decap_8
XFILLER_23_739 VPWR VGND sg13g2_decap_8
X_3993_ _1368_ _1349_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[1\]
+ net797 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2944_ _0414_ _0444_ _0445_ VPWR VGND sg13g2_nor2_1
XFILLER_31_761 VPWR VGND sg13g2_decap_8
X_2875_ net793 sap_3_inst.alu_inst.tmp\[0\] _0378_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_990 VPWR VGND sg13g2_decap_8
X_3427_ _0897_ _0865_ _0891_ VPWR VGND sg13g2_nand2_1
X_3358_ _0829_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[2\] net673
+ VPWR VGND sg13g2_nand2_1
X_2309_ _1643_ _1651_ _1657_ _1661_ _1726_ VPWR VGND sg13g2_nor4_1
X_3289_ _0760_ _0690_ _0748_ VPWR VGND sg13g2_nand2_1
XFILLER_39_872 VPWR VGND sg13g2_decap_8
XFILLER_26_544 VPWR VGND sg13g2_decap_8
XFILLER_41_558 VPWR VGND sg13g2_decap_8
XFILLER_10_912 VPWR VGND sg13g2_decap_8
XFILLER_16_1003 VPWR VGND sg13g2_decap_8
XFILLER_10_989 VPWR VGND sg13g2_decap_8
XFILLER_1_632 VPWR VGND sg13g2_decap_8
XFILLER_49_636 VPWR VGND sg13g2_decap_8
XFILLER_45_820 VPWR VGND sg13g2_decap_8
XFILLER_17_555 VPWR VGND sg13g2_decap_8
XFILLER_45_897 VPWR VGND sg13g2_decap_8
XFILLER_32_525 VPWR VGND sg13g2_decap_8
XFILLER_9_732 VPWR VGND sg13g2_decap_8
X_2660_ _2065_ _2066_ _2064_ _2067_ VPWR VGND sg13g2_nand3_1
XFILLER_5_20 VPWR VGND sg13g2_fill_2
X_2591_ _1997_ VPWR _2000_ VGND _1760_ _1999_ sg13g2_o21ai_1
XFILLER_5_982 VPWR VGND sg13g2_decap_8
X_4330_ net817 VGND VPWR _0187_ sap_3_outputReg_serial clknet_3_0__leaf_clk sg13g2_dfrbpq_1
X_4261_ net810 VGND VPWR _0118_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[4\]
+ clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3212_ _1495_ _0636_ _0683_ VPWR VGND sg13g2_nor2_1
X_4192_ net818 VGND VPWR _0049_ sap_3_inst.alu_inst.carry clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3143_ sap_3_inst.controller_inst.opcode\[0\] net31 net717 _0058_ VPWR VGND sg13g2_mux2_1
X_3074_ _0571_ net772 sap_3_inst.alu_inst.tmp\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_36_820 VPWR VGND sg13g2_decap_8
XFILLER_35_363 VPWR VGND sg13g2_fill_2
XFILLER_36_897 VPWR VGND sg13g2_decap_8
XFILLER_23_536 VPWR VGND sg13g2_decap_8
X_3976_ _1335_ _1345_ _1352_ VPWR VGND sg13g2_nor2_2
X_2927_ _0409_ _0421_ net575 _0429_ VPWR VGND _0427_ sg13g2_nand4_1
X_2858_ _0361_ VPWR _0362_ VGND net793 sap_3_inst.alu_inst.tmp\[0\] sg13g2_o21ai_1
X_2789_ _0305_ net15 VPWR VGND sg13g2_inv_4
XFILLER_46_1007 VPWR VGND sg13g2_decap_8
Xfanout700 net701 net700 VPWR VGND sg13g2_buf_8
Xfanout733 _1662_ net733 VPWR VGND sg13g2_buf_8
Xfanout722 _1722_ net722 VPWR VGND sg13g2_buf_8
Xfanout711 net713 net711 VPWR VGND sg13g2_buf_8
Xfanout755 net756 net755 VPWR VGND sg13g2_buf_8
Xfanout766 sap_3_inst.controller_inst.opcode\[2\] net766 VPWR VGND sg13g2_buf_1
Xfanout744 sap_3_inst.controller_inst.stage\[3\] net744 VPWR VGND sg13g2_buf_8
Xfanout799 _0185_ net799 VPWR VGND sg13g2_buf_8
Xfanout788 sap_3_inst.alu_inst.acc\[2\] net788 VPWR VGND sg13g2_buf_8
Xfanout777 sap_3_inst.alu_inst.acc\[6\] net777 VPWR VGND sg13g2_buf_8
XFILLER_27_875 VPWR VGND sg13g2_decap_8
XFILLER_42_856 VPWR VGND sg13g2_decap_8
XFILLER_14_569 VPWR VGND sg13g2_decap_8
XFILLER_14_62 VPWR VGND sg13g2_fill_1
XFILLER_10_786 VPWR VGND sg13g2_decap_8
XFILLER_6_757 VPWR VGND sg13g2_decap_8
XFILLER_2_974 VPWR VGND sg13g2_decap_8
XFILLER_49_433 VPWR VGND sg13g2_decap_8
XFILLER_37_628 VPWR VGND sg13g2_decap_8
XFILLER_18_886 VPWR VGND sg13g2_decap_8
XFILLER_45_694 VPWR VGND sg13g2_decap_8
XFILLER_33_834 VPWR VGND sg13g2_decap_8
X_3830_ _1239_ _1022_ net686 VPWR VGND sg13g2_nand2b_1
XFILLER_20_539 VPWR VGND sg13g2_decap_8
X_3761_ net569 _0304_ net603 _1195_ VPWR VGND sg13g2_mux2_1
X_2712_ _0242_ net617 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[0\]
+ net625 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[0\] VPWR VGND sg13g2_a22oi_1
X_3692_ _1135_ _1137_ _1140_ _1141_ VPWR VGND sg13g2_nor3_1
X_4151__9 VPWR net43 clknet_leaf_2_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
X_2643_ net18 _2051_ VPWR VGND sg13g2_inv_2
X_2574_ _1985_ net614 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[4\]
+ net624 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4313_ net824 VGND VPWR _0170_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[1\]
+ clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4244_ net829 VGND VPWR _0101_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[3\]
+ clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4175_ net819 VGND VPWR _0032_ sap_3_inst.alu_flags\[7\] net47 sg13g2_dfrbpq_1
X_3126_ VGND VPWR net730 _1595_ _0613_ _1874_ sg13g2_a21oi_1
XFILLER_28_617 VPWR VGND sg13g2_decap_8
X_3057_ _0554_ _0542_ _0555_ VPWR VGND sg13g2_xor2_1
XFILLER_24_801 VPWR VGND sg13g2_decap_8
XFILLER_36_694 VPWR VGND sg13g2_decap_8
XFILLER_24_878 VPWR VGND sg13g2_decap_8
X_3959_ _1335_ net802 VPWR VGND net801 sg13g2_nand2b_2
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_749 VPWR VGND sg13g2_decap_8
Xfanout574 _0967_ net574 VPWR VGND sg13g2_buf_1
Xfanout596 net597 net596 VPWR VGND sg13g2_buf_8
Xfanout585 _0881_ net585 VPWR VGND sg13g2_buf_8
XFILLER_46_447 VPWR VGND sg13g2_decap_8
XFILLER_15_812 VPWR VGND sg13g2_decap_8
XFILLER_27_672 VPWR VGND sg13g2_decap_8
XFILLER_42_653 VPWR VGND sg13g2_decap_8
XFILLER_15_889 VPWR VGND sg13g2_decap_8
XFILLER_30_826 VPWR VGND sg13g2_decap_8
XFILLER_41_71 VPWR VGND sg13g2_fill_1
XFILLER_6_554 VPWR VGND sg13g2_decap_8
XFILLER_10_583 VPWR VGND sg13g2_decap_8
XFILLER_29_1013 VPWR VGND sg13g2_decap_8
Xclkbuf_5_3__f_sap_3_inst.alu_inst.clk_regs clknet_4_1_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
X_2290_ net733 _1706_ _1707_ VPWR VGND sg13g2_nor2_2
XFILLER_2_771 VPWR VGND sg13g2_decap_8
XFILLER_38_937 VPWR VGND sg13g2_decap_8
XFILLER_37_436 VPWR VGND sg13g2_fill_2
Xclkbuf_4_8_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_8_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_45_491 VPWR VGND sg13g2_decap_8
XFILLER_18_683 VPWR VGND sg13g2_decap_8
XFILLER_33_631 VPWR VGND sg13g2_decap_8
XFILLER_21_804 VPWR VGND sg13g2_decap_8
X_3813_ net657 _1084_ _1230_ VPWR VGND sg13g2_nor2_1
XFILLER_32_196 VPWR VGND sg13g2_fill_2
X_3744_ _0100_ _1177_ _1180_ net655 _1504_ VPWR VGND sg13g2_a22oi_1
X_3675_ _1125_ net609 _1006_ VPWR VGND sg13g2_nand2_1
X_2626_ _2035_ _2031_ _2034_ net630 _1510_ VPWR VGND sg13g2_a22oi_1
X_2557_ VGND VPWR net710 net569 _0030_ _1968_ sg13g2_a21oi_1
X_2488_ VGND VPWR net8 _1884_ _1905_ _1904_ sg13g2_a21oi_1
X_4227_ net828 VGND VPWR _0084_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[2\]
+ clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_28_403 VPWR VGND sg13g2_fill_2
XFILLER_29_915 VPWR VGND sg13g2_decap_8
X_4158_ net821 VGND VPWR _0019_ u_ser.shadow_reg\[2\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_918 VPWR VGND sg13g2_decap_8
X_3109_ net774 sap_3_inst.out\[7\] net706 _0048_ VPWR VGND sg13g2_mux2_1
X_4089_ _1448_ sap_3_inst.alu_inst.act\[1\] net579 VPWR VGND sg13g2_nand2_1
XFILLER_36_480 VPWR VGND sg13g2_fill_2
XFILLER_37_992 VPWR VGND sg13g2_decap_8
XFILLER_36_491 VPWR VGND sg13g2_decap_8
XFILLER_24_675 VPWR VGND sg13g2_decap_8
XFILLER_8_808 VPWR VGND sg13g2_decap_8
XFILLER_3_546 VPWR VGND sg13g2_decap_8
XFILLER_11_52 VPWR VGND sg13g2_fill_2
XFILLER_4_1026 VPWR VGND sg13g2_fill_2
XFILLER_47_767 VPWR VGND sg13g2_decap_8
XFILLER_19_469 VPWR VGND sg13g2_decap_8
XFILLER_35_918 VPWR VGND sg13g2_decap_8
XFILLER_28_981 VPWR VGND sg13g2_decap_8
XFILLER_43_962 VPWR VGND sg13g2_decap_8
XFILLER_42_450 VPWR VGND sg13g2_decap_8
XFILLER_15_686 VPWR VGND sg13g2_decap_8
XFILLER_30_623 VPWR VGND sg13g2_decap_8
XFILLER_7_863 VPWR VGND sg13g2_decap_8
X_3460_ net587 _0928_ _0929_ VPWR VGND sg13g2_nor2_2
XFILLER_42_4 VPWR VGND sg13g2_fill_1
X_2411_ _1569_ VPWR _1828_ VGND _1811_ _1827_ sg13g2_o21ai_1
X_3391_ _0814_ _0859_ _0803_ _0862_ VPWR VGND sg13g2_nand3_1
X_2342_ _1592_ _1758_ _1759_ VPWR VGND sg13g2_nor2_2
XFILLER_42_1010 VPWR VGND sg13g2_decap_8
X_2273_ _1562_ net749 _1690_ VPWR VGND sg13g2_nor2_1
X_4012_ _1385_ _1352_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[3\]
+ _1340_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_38_734 VPWR VGND sg13g2_decap_8
XFILLER_26_929 VPWR VGND sg13g2_decap_8
XFILLER_18_480 VPWR VGND sg13g2_decap_8
XFILLER_34_962 VPWR VGND sg13g2_decap_8
XFILLER_21_601 VPWR VGND sg13g2_decap_8
XFILLER_21_678 VPWR VGND sg13g2_decap_8
X_3727_ _1165_ VPWR _1166_ VGND net31 net603 sg13g2_o21ai_1
X_3658_ VPWR VGND net11 _0732_ net604 net19 _1111_ _0874_ sg13g2_a221oi_1
X_2609_ net760 _1996_ _2018_ VPWR VGND sg13g2_and2_1
X_3589_ VGND VPWR _1545_ net597 _0073_ _1052_ sg13g2_a21oi_1
XFILLER_29_712 VPWR VGND sg13g2_decap_8
XFILLER_28_222 VPWR VGND sg13g2_fill_2
XFILLER_44_715 VPWR VGND sg13g2_decap_8
XFILLER_29_789 VPWR VGND sg13g2_decap_8
XFILLER_16_439 VPWR VGND sg13g2_fill_2
XFILLER_28_288 VPWR VGND sg13g2_fill_1
XFILLER_19_1001 VPWR VGND sg13g2_decap_8
XFILLER_25_940 VPWR VGND sg13g2_decap_8
XFILLER_24_472 VPWR VGND sg13g2_decap_8
XFILLER_40_954 VPWR VGND sg13g2_decap_8
XFILLER_8_605 VPWR VGND sg13g2_decap_8
XFILLER_12_667 VPWR VGND sg13g2_decap_8
XFILLER_4_844 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_26_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_564 VPWR VGND sg13g2_decap_8
XFILLER_35_715 VPWR VGND sg13g2_decap_8
XFILLER_16_940 VPWR VGND sg13g2_decap_8
X_2960_ _0461_ _0460_ _0344_ _0456_ net704 VPWR VGND sg13g2_a22oi_1
X_2891_ _0376_ VPWR _0394_ VGND _1487_ _0343_ sg13g2_o21ai_1
XFILLER_15_483 VPWR VGND sg13g2_decap_8
XFILLER_31_943 VPWR VGND sg13g2_decap_8
XFILLER_33_1009 VPWR VGND sg13g2_decap_8
XFILLER_30_497 VPWR VGND sg13g2_decap_8
XFILLER_8_97 VPWR VGND sg13g2_decap_4
XFILLER_7_660 VPWR VGND sg13g2_decap_8
X_3512_ _0979_ _0944_ net573 VPWR VGND sg13g2_xnor2_1
X_3443_ _0912_ net639 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[2\]
+ net642 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[2\] VPWR VGND sg13g2_a22oi_1
X_3374_ _1518_ net689 _0746_ _0845_ VPWR VGND sg13g2_nor3_1
X_2325_ _1742_ _1640_ _1726_ VPWR VGND sg13g2_nand2_1
X_2256_ _1673_ _1584_ net732 VPWR VGND sg13g2_nand2_2
XFILLER_38_531 VPWR VGND sg13g2_decap_8
X_2187_ net753 net755 net766 _1604_ VPWR VGND sg13g2_nand3_1
XFILLER_26_726 VPWR VGND sg13g2_decap_8
XFILLER_25_258 VPWR VGND sg13g2_fill_1
XFILLER_22_921 VPWR VGND sg13g2_decap_8
XFILLER_21_475 VPWR VGND sg13g2_decap_8
XFILLER_22_998 VPWR VGND sg13g2_decap_8
XFILLER_1_814 VPWR VGND sg13g2_decap_8
XFILLER_49_818 VPWR VGND sg13g2_decap_8
XFILLER_48_339 VPWR VGND sg13g2_decap_8
XFILLER_44_512 VPWR VGND sg13g2_decap_8
XFILLER_17_737 VPWR VGND sg13g2_decap_8
XFILLER_29_586 VPWR VGND sg13g2_decap_8
XFILLER_32_707 VPWR VGND sg13g2_decap_8
XFILLER_44_589 VPWR VGND sg13g2_decap_8
XFILLER_13_921 VPWR VGND sg13g2_decap_8
XFILLER_24_280 VPWR VGND sg13g2_decap_4
XFILLER_40_751 VPWR VGND sg13g2_decap_8
XFILLER_9_914 VPWR VGND sg13g2_decap_8
XFILLER_13_998 VPWR VGND sg13g2_decap_8
XFILLER_8_479 VPWR VGND sg13g2_decap_8
XFILLER_4_641 VPWR VGND sg13g2_decap_8
X_3090_ _0522_ _0586_ _0348_ _0587_ VPWR VGND sg13g2_nand3_1
X_2110_ VPWR _1528_ sap_3_inst.alu_inst.tmp\[6\] VGND sg13g2_inv_1
Xhold2 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[3\] VPWR VGND net49
+ sg13g2_dlygate4sd3_1
XFILLER_47_361 VPWR VGND sg13g2_decap_8
XFILLER_35_512 VPWR VGND sg13g2_decap_8
XFILLER_23_718 VPWR VGND sg13g2_decap_8
X_3992_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[1\] _1352_
+ _1367_ net794 sg13g2_a21oi_1
XFILLER_35_589 VPWR VGND sg13g2_decap_8
X_2943_ _0444_ _0439_ _0442_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_740 VPWR VGND sg13g2_decap_8
X_2874_ net575 _0376_ _0377_ VPWR VGND sg13g2_nor2_1
XFILLER_30_294 VPWR VGND sg13g2_fill_1
X_3426_ _0896_ net594 _0895_ VPWR VGND sg13g2_nand2_1
X_3357_ _0828_ net677 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[2\]
+ net684 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2308_ VGND VPWR net758 _1657_ _1725_ _1651_ sg13g2_a21oi_1
XFILLER_45_309 VPWR VGND sg13g2_fill_1
X_3288_ _0690_ _0748_ _0759_ VPWR VGND sg13g2_and2_1
XFILLER_39_851 VPWR VGND sg13g2_decap_8
X_2239_ _1656_ net758 VPWR VGND net759 sg13g2_nand2b_2
XFILLER_26_523 VPWR VGND sg13g2_decap_8
XFILLER_41_537 VPWR VGND sg13g2_decap_8
XFILLER_22_795 VPWR VGND sg13g2_decap_8
XFILLER_10_968 VPWR VGND sg13g2_decap_8
XFILLER_6_939 VPWR VGND sg13g2_decap_8
XFILLER_1_611 VPWR VGND sg13g2_decap_8
XFILLER_49_615 VPWR VGND sg13g2_decap_8
XFILLER_1_688 VPWR VGND sg13g2_decap_8
XFILLER_23_1019 VPWR VGND sg13g2_decap_8
XFILLER_17_534 VPWR VGND sg13g2_decap_8
XFILLER_45_876 VPWR VGND sg13g2_decap_8
XFILLER_32_504 VPWR VGND sg13g2_decap_8
XFILLER_44_397 VPWR VGND sg13g2_fill_2
XFILLER_44_386 VPWR VGND sg13g2_decap_8
XFILLER_9_711 VPWR VGND sg13g2_decap_8
XFILLER_8_210 VPWR VGND sg13g2_fill_1
XFILLER_13_795 VPWR VGND sg13g2_decap_8
XFILLER_9_788 VPWR VGND sg13g2_decap_8
X_2590_ _1999_ _1998_ _1600_ VPWR VGND sg13g2_nand2b_1
XFILLER_5_961 VPWR VGND sg13g2_decap_8
XFILLER_5_54 VPWR VGND sg13g2_fill_1
XFILLER_5_98 VPWR VGND sg13g2_fill_1
X_4260_ net831 VGND VPWR _0117_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[3\]
+ clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3211_ net715 _0681_ _0682_ VPWR VGND sg13g2_nor2_1
X_4191_ net818 VGND VPWR _0048_ sap_3_inst.out\[7\] clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3142_ VGND VPWR _1529_ net701 _0057_ _0621_ sg13g2_a21oi_1
XFILLER_39_136 VPWR VGND sg13g2_fill_1
X_3073_ net772 sap_3_inst.alu_inst.tmp\[7\] _0570_ VPWR VGND sg13g2_nor2_1
XFILLER_39_1026 VPWR VGND sg13g2_fill_2
XFILLER_23_515 VPWR VGND sg13g2_decap_8
XFILLER_36_876 VPWR VGND sg13g2_decap_8
X_3975_ _1339_ _1341_ _1351_ VPWR VGND sg13g2_nor2_2
X_2926_ _0346_ VPWR _0428_ VGND _0349_ _0380_ sg13g2_o21ai_1
X_2857_ _2013_ _2019_ _0361_ VPWR VGND sg13g2_nor2_2
X_2788_ _0305_ net576 VPWR VGND _1928_ sg13g2_nand2b_2
Xfanout701 _0615_ net701 VPWR VGND sg13g2_buf_8
Xfanout723 _1722_ net723 VPWR VGND sg13g2_buf_1
Xfanout712 net713 net712 VPWR VGND sg13g2_buf_2
X_3409_ _0880_ _0870_ _0879_ VPWR VGND sg13g2_nand2_1
Xfanout734 _1661_ net734 VPWR VGND sg13g2_buf_8
Xfanout767 net768 net767 VPWR VGND sg13g2_buf_8
Xfanout745 sap_3_inst.controller_inst.stage\[2\] net745 VPWR VGND sg13g2_buf_8
Xfanout756 sap_3_inst.controller_inst.opcode\[6\] net756 VPWR VGND sg13g2_buf_8
Xfanout778 net779 net778 VPWR VGND sg13g2_buf_8
Xfanout789 net791 net789 VPWR VGND sg13g2_buf_8
XFILLER_46_629 VPWR VGND sg13g2_decap_8
XFILLER_26_331 VPWR VGND sg13g2_decap_4
XFILLER_27_854 VPWR VGND sg13g2_decap_8
XFILLER_42_835 VPWR VGND sg13g2_decap_8
XFILLER_14_548 VPWR VGND sg13g2_decap_8
XFILLER_22_592 VPWR VGND sg13g2_decap_8
XFILLER_6_736 VPWR VGND sg13g2_decap_8
XFILLER_10_765 VPWR VGND sg13g2_decap_8
XFILLER_5_235 VPWR VGND sg13g2_fill_1
XFILLER_2_953 VPWR VGND sg13g2_decap_8
XFILLER_49_412 VPWR VGND sg13g2_decap_8
XFILLER_7_1024 VPWR VGND sg13g2_decap_4
XFILLER_1_485 VPWR VGND sg13g2_decap_8
XFILLER_37_607 VPWR VGND sg13g2_decap_8
XFILLER_49_489 VPWR VGND sg13g2_decap_8
XFILLER_45_673 VPWR VGND sg13g2_decap_8
XFILLER_18_865 VPWR VGND sg13g2_decap_8
XFILLER_33_813 VPWR VGND sg13g2_decap_8
X_3760_ _0993_ _1193_ _1194_ VPWR VGND sg13g2_nor2_1
XFILLER_20_518 VPWR VGND sg13g2_decap_8
XFILLER_32_378 VPWR VGND sg13g2_fill_1
XFILLER_13_592 VPWR VGND sg13g2_decap_8
X_2711_ _1809_ net627 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[0\]
+ _0241_ VPWR VGND sg13g2_nand3_1
X_3691_ VGND VPWR _1140_ _1139_ net609 sg13g2_or2_1
XFILLER_9_585 VPWR VGND sg13g2_decap_8
X_2642_ _2036_ _2039_ _2040_ _2051_ VGND VPWR _2050_ sg13g2_nor4_2
X_2573_ _1984_ _1857_ _1983_ VPWR VGND sg13g2_nand2_1
X_4312_ net829 VGND VPWR _0169_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[0\]
+ clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4243_ net806 VGND VPWR _0100_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[2\]
+ clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4174_ net805 VGND VPWR _0031_ sap_3_inst.alu_flags\[6\] net46 sg13g2_dfrbpq_1
X_3125_ VGND VPWR _0607_ _0611_ _0049_ _0612_ sg13g2_a21oi_1
X_3056_ _0507_ VPWR _0554_ VGND _0506_ _0518_ sg13g2_o21ai_1
XFILLER_42_109 VPWR VGND sg13g2_fill_1
XFILLER_36_673 VPWR VGND sg13g2_decap_8
XFILLER_23_312 VPWR VGND sg13g2_fill_2
XFILLER_24_857 VPWR VGND sg13g2_decap_8
X_3958_ VGND VPWR _0155_ _1334_ _0160_ _1324_ sg13g2_a21oi_1
X_3889_ VGND VPWR net672 _1081_ _0143_ _1282_ sg13g2_a21oi_1
X_2909_ _0410_ VPWR _0411_ VGND _0374_ _0378_ sg13g2_o21ai_1
XFILLER_3_728 VPWR VGND sg13g2_decap_8
Xfanout575 _0354_ net575 VPWR VGND sg13g2_buf_8
XFILLER_47_949 VPWR VGND sg13g2_decap_8
Xfanout597 _0741_ net597 VPWR VGND sg13g2_buf_8
Xfanout586 net587 net586 VPWR VGND sg13g2_buf_8
XFILLER_46_426 VPWR VGND sg13g2_decap_8
XFILLER_27_651 VPWR VGND sg13g2_decap_8
XFILLER_42_632 VPWR VGND sg13g2_decap_8
XFILLER_15_868 VPWR VGND sg13g2_decap_8
XFILLER_30_805 VPWR VGND sg13g2_decap_8
XFILLER_25_73 VPWR VGND sg13g2_fill_1
XFILLER_10_562 VPWR VGND sg13g2_decap_8
XFILLER_6_533 VPWR VGND sg13g2_decap_8
XFILLER_2_750 VPWR VGND sg13g2_decap_8
XFILLER_2_22 VPWR VGND sg13g2_fill_1
XFILLER_49_264 VPWR VGND sg13g2_decap_8
XFILLER_38_916 VPWR VGND sg13g2_decap_8
XFILLER_49_286 VPWR VGND sg13g2_decap_8
XFILLER_18_662 VPWR VGND sg13g2_decap_8
XFILLER_46_993 VPWR VGND sg13g2_decap_8
XFILLER_45_470 VPWR VGND sg13g2_decap_8
XFILLER_33_610 VPWR VGND sg13g2_decap_8
XFILLER_32_131 VPWR VGND sg13g2_fill_2
X_3812_ _1228_ VPWR _0119_ VGND _1007_ _1229_ sg13g2_o21ai_1
XFILLER_33_687 VPWR VGND sg13g2_decap_8
X_3743_ VPWR VGND _1179_ net655 _1110_ net608 _1180_ _0928_ sg13g2_a221oi_1
X_3674_ net610 _1006_ _1124_ VPWR VGND sg13g2_and2_1
X_2625_ _2025_ _2027_ _2032_ _2033_ _2034_ VPWR VGND sg13g2_and4_1
X_2556_ sap_3_inst.alu_flags\[5\] net710 _1968_ VPWR VGND sg13g2_nor2_1
X_2487_ VGND VPWR net695 _1903_ _1904_ _1901_ sg13g2_a21oi_1
X_4226_ net805 VGND VPWR _0083_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4157_ net821 VGND VPWR _0018_ u_ser.shadow_reg\[1\] clknet_3_2__leaf_clk sg13g2_dfrbpq_1
X_3108_ net775 sap_3_inst.out\[6\] net706 _0047_ VPWR VGND sg13g2_mux2_1
Xclkbuf_5_27__f_sap_3_inst.alu_inst.clk_regs clknet_4_13_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
X_4088_ _1446_ VPWR _1447_ VGND net790 net698 sg13g2_o21ai_1
XFILLER_37_971 VPWR VGND sg13g2_decap_8
XFILLER_43_429 VPWR VGND sg13g2_decap_4
X_3039_ _0536_ _0502_ _0535_ _0537_ VPWR VGND sg13g2_a21o_1
XFILLER_24_654 VPWR VGND sg13g2_decap_8
XFILLER_12_849 VPWR VGND sg13g2_decap_8
XFILLER_23_186 VPWR VGND sg13g2_fill_2
XFILLER_20_882 VPWR VGND sg13g2_decap_8
XFILLER_3_525 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_fill_2
XFILLER_4_1005 VPWR VGND sg13g2_decap_8
XFILLER_47_746 VPWR VGND sg13g2_decap_8
Xclkbuf_5_16__f_sap_3_inst.alu_inst.clk_regs clknet_4_8_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_28_960 VPWR VGND sg13g2_decap_8
XFILLER_43_941 VPWR VGND sg13g2_decap_8
XFILLER_15_665 VPWR VGND sg13g2_decap_8
XFILLER_30_602 VPWR VGND sg13g2_decap_8
XFILLER_30_679 VPWR VGND sg13g2_decap_8
XFILLER_7_842 VPWR VGND sg13g2_decap_8
X_2410_ net719 _1825_ _1826_ _1827_ VPWR VGND sg13g2_nor3_1
X_3390_ _0861_ _0814_ _0859_ VPWR VGND sg13g2_nand2_2
X_2341_ net750 VPWR _1758_ VGND _1573_ _1616_ sg13g2_o21ai_1
X_2272_ _1649_ VPWR _1689_ VGND _1687_ _1688_ sg13g2_o21ai_1
X_4011_ _1384_ _1353_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[3\]
+ _1347_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_38_713 VPWR VGND sg13g2_decap_8
XFILLER_26_908 VPWR VGND sg13g2_decap_8
XFILLER_25_429 VPWR VGND sg13g2_decap_8
XFILLER_46_790 VPWR VGND sg13g2_decap_8
XFILLER_34_941 VPWR VGND sg13g2_decap_8
XFILLER_20_134 VPWR VGND sg13g2_fill_1
XFILLER_21_657 VPWR VGND sg13g2_decap_8
X_3726_ _1165_ _0301_ net603 VPWR VGND sg13g2_nand2_1
X_3657_ _1110_ _0227_ net668 VPWR VGND sg13g2_nand2_1
X_2608_ _2015_ VPWR _2017_ VGND net733 _1673_ sg13g2_o21ai_1
X_3588_ VPWR VGND net607 _1051_ _1048_ _1042_ _1052_ _1044_ sg13g2_a221oi_1
X_2539_ _1946_ _1950_ _1944_ _1952_ VPWR VGND _1951_ sg13g2_nand4_1
XFILLER_0_539 VPWR VGND sg13g2_decap_8
X_4209_ net813 VGND VPWR _0066_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[0\]
+ clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_17_919 VPWR VGND sg13g2_decap_8
XFILLER_29_768 VPWR VGND sg13g2_decap_8
XFILLER_24_451 VPWR VGND sg13g2_decap_8
XFILLER_25_996 VPWR VGND sg13g2_decap_8
XFILLER_40_933 VPWR VGND sg13g2_decap_8
XFILLER_12_646 VPWR VGND sg13g2_decap_8
XFILLER_4_823 VPWR VGND sg13g2_decap_8
XFILLER_26_1006 VPWR VGND sg13g2_decap_8
XFILLER_47_543 VPWR VGND sg13g2_decap_8
XFILLER_34_204 VPWR VGND sg13g2_fill_1
XFILLER_34_248 VPWR VGND sg13g2_fill_1
XFILLER_15_462 VPWR VGND sg13g2_decap_8
XFILLER_16_996 VPWR VGND sg13g2_decap_8
X_2890_ _0342_ _0374_ net748 _0393_ VPWR VGND sg13g2_nand3_1
XFILLER_31_922 VPWR VGND sg13g2_decap_8
XFILLER_31_999 VPWR VGND sg13g2_decap_8
X_3511_ net590 net571 net573 _0978_ VPWR VGND sg13g2_nor3_1
X_3442_ _0911_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[2\] net670
+ VPWR VGND sg13g2_nand2_1
X_3373_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[1\] net670 _0844_
+ VPWR VGND sg13g2_and2_1
X_2324_ _1738_ _1739_ _1729_ _1741_ VPWR VGND _1740_ sg13g2_nand4_1
X_2255_ net738 net732 _1672_ VPWR VGND sg13g2_and2_1
XFILLER_38_510 VPWR VGND sg13g2_decap_8
X_2186_ _1603_ net765 net753 net755 VPWR VGND sg13g2_and3_2
XFILLER_26_705 VPWR VGND sg13g2_decap_8
XFILLER_38_587 VPWR VGND sg13g2_decap_8
XFILLER_25_226 VPWR VGND sg13g2_fill_2
XFILLER_41_719 VPWR VGND sg13g2_decap_8
XFILLER_22_900 VPWR VGND sg13g2_decap_8
XFILLER_22_977 VPWR VGND sg13g2_decap_8
X_3709_ _1154_ _1065_ VPWR VGND _0925_ sg13g2_nand2b_2
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_48_318 VPWR VGND sg13g2_decap_8
XFILLER_17_716 VPWR VGND sg13g2_decap_8
XFILLER_29_565 VPWR VGND sg13g2_decap_8
XFILLER_44_568 VPWR VGND sg13g2_decap_8
XFILLER_13_900 VPWR VGND sg13g2_decap_8
XFILLER_40_730 VPWR VGND sg13g2_decap_8
XFILLER_25_793 VPWR VGND sg13g2_decap_8
XFILLER_13_977 VPWR VGND sg13g2_decap_8
XFILLER_8_436 VPWR VGND sg13g2_fill_1
XFILLER_8_447 VPWR VGND sg13g2_fill_1
XFILLER_4_620 VPWR VGND sg13g2_decap_8
XFILLER_3_141 VPWR VGND sg13g2_fill_1
XFILLER_4_697 VPWR VGND sg13g2_decap_8
Xhold3 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[2\] VPWR VGND net50
+ sg13g2_dlygate4sd3_1
XFILLER_47_340 VPWR VGND sg13g2_decap_8
XFILLER_48_885 VPWR VGND sg13g2_decap_8
X_3991_ _1366_ _1351_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[1\]
+ net796 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[1\] VPWR VGND sg13g2_a22oi_1
XFILLER_35_568 VPWR VGND sg13g2_decap_8
X_2942_ _0440_ _0442_ _0443_ VPWR VGND sg13g2_nor2_1
XFILLER_16_793 VPWR VGND sg13g2_decap_8
X_2873_ _0374_ _0341_ _0376_ VPWR VGND sg13g2_xor2_1
XFILLER_31_796 VPWR VGND sg13g2_decap_8
X_3425_ _0884_ VPWR _0895_ VGND net660 _0894_ sg13g2_o21ai_1
X_3356_ _0827_ net681 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[2\]
+ net688 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[2\] VPWR VGND sg13g2_a22oi_1
X_2307_ VGND VPWR _1617_ net722 _1724_ _1590_ sg13g2_a21oi_1
X_3287_ _0758_ _0666_ _0690_ VPWR VGND sg13g2_nand2_2
XFILLER_39_830 VPWR VGND sg13g2_decap_8
X_2238_ net761 net757 _1655_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_502 VPWR VGND sg13g2_decap_8
X_2169_ net747 net746 _1586_ VPWR VGND sg13g2_nor2b_2
XFILLER_41_516 VPWR VGND sg13g2_decap_8
XFILLER_26_579 VPWR VGND sg13g2_decap_8
XFILLER_22_774 VPWR VGND sg13g2_decap_8
XFILLER_6_918 VPWR VGND sg13g2_decap_8
XFILLER_10_947 VPWR VGND sg13g2_decap_8
XFILLER_1_667 VPWR VGND sg13g2_decap_8
XFILLER_48_115 VPWR VGND sg13g2_fill_1
XFILLER_17_513 VPWR VGND sg13g2_decap_8
XFILLER_45_855 VPWR VGND sg13g2_decap_8
XFILLER_25_590 VPWR VGND sg13g2_decap_8
XFILLER_13_774 VPWR VGND sg13g2_decap_8
XFILLER_9_767 VPWR VGND sg13g2_decap_8
XFILLER_5_940 VPWR VGND sg13g2_decap_8
XFILLER_4_494 VPWR VGND sg13g2_decap_8
X_3210_ VGND VPWR _0279_ _0680_ _0681_ _1752_ sg13g2_a21oi_1
X_4190_ net821 VGND VPWR _0047_ sap_3_inst.out\[6\] clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3141_ net24 net701 _0621_ VPWR VGND sg13g2_nor2_1
X_3072_ _0569_ _0567_ _0568_ VPWR VGND sg13g2_xnor2_1
XFILLER_48_682 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk_div_out clk_div_out clknet_0_clk_div_out VPWR VGND sg13g2_buf_8
XFILLER_36_855 VPWR VGND sg13g2_decap_8
XFILLER_47_192 VPWR VGND sg13g2_fill_1
XFILLER_39_1005 VPWR VGND sg13g2_decap_8
X_3974_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[0\] sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[1\]
+ _1341_ _1350_ VPWR VGND sg13g2_nor3_2
XFILLER_16_590 VPWR VGND sg13g2_decap_8
X_2925_ VPWR VGND net783 _0426_ net691 net789 _0427_ net692 sg13g2_a221oi_1
X_2856_ VPWR VGND net789 net703 net691 net692 _0360_ _0358_ sg13g2_a221oi_1
XFILLER_31_593 VPWR VGND sg13g2_decap_8
X_2787_ net14 _0304_ VPWR VGND sg13g2_inv_2
Xfanout713 _1796_ net713 VPWR VGND sg13g2_buf_8
Xfanout724 _1631_ net724 VPWR VGND sg13g2_buf_8
Xfanout702 net703 net702 VPWR VGND sg13g2_buf_8
X_3408_ VGND VPWR _0877_ _0878_ _0879_ net596 sg13g2_a21oi_1
Xfanout735 _1652_ net735 VPWR VGND sg13g2_buf_8
Xfanout757 net758 net757 VPWR VGND sg13g2_buf_8
Xfanout746 sap_3_inst.controller_inst.stage\[1\] net746 VPWR VGND sg13g2_buf_8
XFILLER_46_608 VPWR VGND sg13g2_decap_8
Xfanout779 net780 net779 VPWR VGND sg13g2_buf_2
Xfanout768 net769 net768 VPWR VGND sg13g2_buf_8
X_3339_ _1499_ net662 _0810_ VPWR VGND sg13g2_nor2_1
Xclkbuf_4_9_0_sap_3_inst.alu_inst.clk_regs clknet_0_sap_3_inst.alu_inst.clk_regs clknet_4_9_0_sap_3_inst.alu_inst.clk_regs
+ VPWR VGND sg13g2_buf_8
XFILLER_27_833 VPWR VGND sg13g2_decap_8
XFILLER_42_814 VPWR VGND sg13g2_decap_8
XFILLER_14_527 VPWR VGND sg13g2_decap_8
XFILLER_41_346 VPWR VGND sg13g2_fill_2
XFILLER_22_571 VPWR VGND sg13g2_decap_8
XFILLER_10_744 VPWR VGND sg13g2_decap_8
XFILLER_6_715 VPWR VGND sg13g2_decap_8
XFILLER_30_63 VPWR VGND sg13g2_fill_2
XFILLER_2_932 VPWR VGND sg13g2_decap_8
XFILLER_7_1003 VPWR VGND sg13g2_decap_8
XFILLER_1_464 VPWR VGND sg13g2_decap_8
XFILLER_49_468 VPWR VGND sg13g2_decap_8
XFILLER_18_844 VPWR VGND sg13g2_decap_8
XFILLER_45_652 VPWR VGND sg13g2_decap_8
XFILLER_33_869 VPWR VGND sg13g2_decap_8
XFILLER_41_880 VPWR VGND sg13g2_decap_8
XFILLER_13_571 VPWR VGND sg13g2_decap_8
X_2710_ _0240_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[0\] net623
+ VPWR VGND sg13g2_nand2_1
XFILLER_9_564 VPWR VGND sg13g2_decap_8
X_3690_ _0720_ _0731_ _0864_ _1138_ _1139_ VPWR VGND sg13g2_and4_1
X_2641_ VGND VPWR _2044_ _2049_ _2050_ _1720_ sg13g2_a21oi_1
X_2572_ _1983_ net616 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[4\]
+ net628 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[4\] VPWR VGND sg13g2_a22oi_1
X_4311_ net833 VGND VPWR _0168_ sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[7\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
X_4242_ net805 VGND VPWR _0099_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4173_ net804 VGND VPWR _0030_ sap_3_inst.alu_flags\[5\] net45 sg13g2_dfrbpq_1
X_3124_ sap_3_inst.alu_inst.carry _0608_ _0612_ VPWR VGND sg13g2_nor2_1
X_3055_ _0553_ _0522_ _0547_ VPWR VGND sg13g2_xnor2_1
XFILLER_36_652 VPWR VGND sg13g2_decap_8
XFILLER_24_836 VPWR VGND sg13g2_decap_8
XFILLER_35_184 VPWR VGND sg13g2_fill_2
X_3957_ _1334_ _1333_ _1315_ _1318_ net48 VPWR VGND sg13g2_a22oi_1
X_2908_ _0410_ net790 sap_3_inst.alu_inst.tmp\[1\] VPWR VGND sg13g2_nand2b_1
X_3888_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[5\] net672 _1282_
+ VPWR VGND sg13g2_nor2_1
XFILLER_13_1019 VPWR VGND sg13g2_decap_8
X_2839_ _0343_ net792 sap_3_inst.alu_inst.tmp\[0\] VPWR VGND sg13g2_xnor2_1
XFILLER_3_707 VPWR VGND sg13g2_decap_8
XFILLER_4_8 VPWR VGND sg13g2_fill_1
XFILLER_47_928 VPWR VGND sg13g2_decap_8
XFILLER_46_405 VPWR VGND sg13g2_decap_8
Xfanout598 net599 net598 VPWR VGND sg13g2_buf_2
Xfanout587 net588 net587 VPWR VGND sg13g2_buf_8
Xfanout576 _1721_ net576 VPWR VGND sg13g2_buf_8
XFILLER_27_630 VPWR VGND sg13g2_decap_8
XFILLER_42_611 VPWR VGND sg13g2_decap_8
XFILLER_15_847 VPWR VGND sg13g2_decap_8
XFILLER_26_184 VPWR VGND sg13g2_fill_2
XFILLER_42_688 VPWR VGND sg13g2_decap_8
XFILLER_10_541 VPWR VGND sg13g2_decap_8
XFILLER_6_512 VPWR VGND sg13g2_decap_8
XFILLER_6_589 VPWR VGND sg13g2_decap_8
XFILLER_2_34 VPWR VGND sg13g2_fill_2
XFILLER_46_972 VPWR VGND sg13g2_decap_8
XFILLER_18_641 VPWR VGND sg13g2_decap_8
XFILLER_33_666 VPWR VGND sg13g2_decap_8
X_3811_ _1229_ net681 _1079_ VPWR VGND sg13g2_nand2_1
XFILLER_14_891 VPWR VGND sg13g2_decap_8
XFILLER_21_839 VPWR VGND sg13g2_decap_8
X_3742_ VGND VPWR _1179_ _1178_ net11 sg13g2_or2_1
X_3673_ _0086_ _1120_ _1123_ net636 _1534_ VPWR VGND sg13g2_a22oi_1
X_2624_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[1\] net630
+ net624 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[1\] _2033_ net713
+ sg13g2_a221oi_1
X_2555_ net22 net569 VPWR VGND sg13g2_inv_2
X_2486_ _1903_ sap_3_inst.alu_flags\[7\] _1902_ VPWR VGND sg13g2_nand2_1
X_4225_ net816 VGND VPWR _0082_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[0\]
+ clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4156_ net817 VGND VPWR _0017_ u_ser.shadow_reg\[0\] clknet_3_1__leaf_clk sg13g2_dfrbpq_1
X_3107_ net779 sap_3_inst.out\[5\] net706 _0046_ VPWR VGND sg13g2_mux2_1
XFILLER_28_449 VPWR VGND sg13g2_decap_8
X_4087_ _1446_ _0379_ net698 VPWR VGND sg13g2_nand2_1
XFILLER_37_950 VPWR VGND sg13g2_decap_8
X_3038_ _0501_ VPWR _0536_ VGND net778 net709 sg13g2_o21ai_1
XFILLER_24_633 VPWR VGND sg13g2_decap_8
XFILLER_12_828 VPWR VGND sg13g2_decap_8
XFILLER_20_861 VPWR VGND sg13g2_decap_8
XFILLER_3_504 VPWR VGND sg13g2_decap_8
XFILLER_11_65 VPWR VGND sg13g2_fill_2
XFILLER_47_725 VPWR VGND sg13g2_decap_8
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
XFILLER_43_920 VPWR VGND sg13g2_decap_8
XFILLER_34_408 VPWR VGND sg13g2_fill_2
XFILLER_15_644 VPWR VGND sg13g2_decap_8
XFILLER_43_997 VPWR VGND sg13g2_decap_8
XFILLER_42_485 VPWR VGND sg13g2_decap_8
XFILLER_30_658 VPWR VGND sg13g2_decap_8
XFILLER_7_821 VPWR VGND sg13g2_decap_8
XFILLER_11_894 VPWR VGND sg13g2_decap_8
XFILLER_7_898 VPWR VGND sg13g2_decap_8
X_2340_ _1675_ _1746_ _1756_ _1757_ VPWR VGND sg13g2_nor3_1
X_2271_ _1688_ _1682_ _1685_ VPWR VGND sg13g2_nand2_1
X_4010_ _1383_ _1338_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[3\]
+ _1337_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_37_257 VPWR VGND sg13g2_fill_1
XFILLER_38_769 VPWR VGND sg13g2_decap_8
XFILLER_19_994 VPWR VGND sg13g2_decap_8
XFILLER_34_920 VPWR VGND sg13g2_decap_8
XFILLER_37_279 VPWR VGND sg13g2_fill_1
XFILLER_34_997 VPWR VGND sg13g2_decap_8
XFILLER_21_636 VPWR VGND sg13g2_decap_8
X_3725_ net655 net668 _1164_ VPWR VGND sg13g2_nor2_1
X_3656_ VGND VPWR _0917_ _1108_ _1109_ net613 sg13g2_a21oi_1
X_3587_ _1051_ _0742_ _1050_ VPWR VGND sg13g2_nand2_1
X_2607_ VPWR VGND net762 _2014_ _1996_ net734 _2016_ _1672_ sg13g2_a221oi_1
XFILLER_0_518 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_sap_3_inst.alu_inst.clk clknet_1_0__leaf_sap_3_inst.alu_inst.clk clknet_leaf_0_sap_3_inst.alu_inst.clk
+ VPWR VGND sg13g2_buf_8
X_2538_ _1951_ net615 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[5\]
+ _1853_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[5\] VPWR VGND sg13g2_a22oi_1
X_2469_ _1600_ net725 _1886_ VPWR VGND sg13g2_nor2_2
X_4208_ net808 VGND VPWR _0065_ sap_3_inst.controller_inst.opcode\[7\] clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_29_747 VPWR VGND sg13g2_decap_8
X_4139_ net800 _1465_ _1484_ VPWR VGND sg13g2_nor2_1
XFILLER_28_224 VPWR VGND sg13g2_fill_1
XFILLER_24_430 VPWR VGND sg13g2_decap_8
XFILLER_40_912 VPWR VGND sg13g2_decap_8
XFILLER_25_975 VPWR VGND sg13g2_decap_8
XFILLER_11_113 VPWR VGND sg13g2_fill_1
XFILLER_12_625 VPWR VGND sg13g2_decap_8
XFILLER_40_989 VPWR VGND sg13g2_decap_8
XFILLER_11_157 VPWR VGND sg13g2_fill_1
XFILLER_4_802 VPWR VGND sg13g2_decap_8
XFILLER_4_879 VPWR VGND sg13g2_decap_8
XFILLER_47_522 VPWR VGND sg13g2_decap_8
XFILLER_47_599 VPWR VGND sg13g2_decap_8
XFILLER_16_975 VPWR VGND sg13g2_decap_8
XFILLER_31_901 VPWR VGND sg13g2_decap_8
XFILLER_43_794 VPWR VGND sg13g2_decap_8
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_31_978 VPWR VGND sg13g2_decap_8
X_3510_ net571 net574 _0977_ VPWR VGND sg13g2_nor2_1
XFILLER_11_691 VPWR VGND sg13g2_decap_8
XFILLER_7_695 VPWR VGND sg13g2_decap_8
X_3441_ _0910_ net649 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[2\]
+ net673 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[2\] VPWR VGND sg13g2_a22oi_1
X_3372_ _1517_ net689 _0749_ _0843_ VPWR VGND sg13g2_nor3_1
X_2323_ _1704_ _1710_ _1728_ _1730_ _1740_ VPWR VGND sg13g2_nor4_1
X_2254_ sap_3_inst.controller_inst.stage\[2\] net744 _1671_ VPWR VGND sg13g2_nor2b_2
X_2185_ _1600_ VPWR _1602_ VGND net751 _1596_ sg13g2_o21ai_1
XFILLER_19_0 VPWR VGND sg13g2_fill_1
XFILLER_38_566 VPWR VGND sg13g2_decap_8
XFILLER_19_791 VPWR VGND sg13g2_decap_8
XFILLER_34_794 VPWR VGND sg13g2_decap_8
XFILLER_22_956 VPWR VGND sg13g2_decap_8
XFILLER_33_282 VPWR VGND sg13g2_fill_2
XFILLER_49_1007 VPWR VGND sg13g2_decap_8
X_3708_ VPWR _0091_ _1153_ VGND sg13g2_inv_1
X_3639_ _1094_ net595 _0855_ VPWR VGND sg13g2_nand2_1
XFILLER_1_849 VPWR VGND sg13g2_decap_8
XFILLER_29_544 VPWR VGND sg13g2_decap_8
XFILLER_44_547 VPWR VGND sg13g2_decap_8
XFILLER_25_772 VPWR VGND sg13g2_decap_8
XFILLER_13_956 VPWR VGND sg13g2_decap_8
XFILLER_40_786 VPWR VGND sg13g2_decap_8
XFILLER_9_949 VPWR VGND sg13g2_decap_8
XFILLER_32_1022 VPWR VGND sg13g2_decap_8
XFILLER_12_499 VPWR VGND sg13g2_decap_8
XFILLER_4_676 VPWR VGND sg13g2_decap_8
XFILLER_0_882 VPWR VGND sg13g2_decap_8
Xhold4 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[5\] VPWR VGND net51
+ sg13g2_dlygate4sd3_1
XFILLER_48_864 VPWR VGND sg13g2_decap_8
XFILLER_47_396 VPWR VGND sg13g2_decap_8
XFILLER_35_547 VPWR VGND sg13g2_decap_8
X_3990_ _1365_ _1346_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[1\]
+ _1340_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2941_ VGND VPWR _0405_ _0411_ _0442_ _0441_ sg13g2_a21oi_1
XFILLER_16_772 VPWR VGND sg13g2_decap_8
XFILLER_43_591 VPWR VGND sg13g2_decap_8
XFILLER_15_293 VPWR VGND sg13g2_fill_2
X_2872_ _0375_ _0374_ _0341_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_775 VPWR VGND sg13g2_decap_8
XFILLER_7_492 VPWR VGND sg13g2_decap_8
X_3424_ _0894_ _0853_ _0891_ VPWR VGND sg13g2_xnor2_1
X_3355_ _0690_ _0748_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[2\]
+ _0826_ VPWR VGND sg13g2_nand3_1
X_2306_ _1723_ _1553_ net736 VPWR VGND sg13g2_nand2_2
X_3286_ VPWR VGND _0689_ _0665_ _0688_ _0648_ _0757_ _0651_ sg13g2_a221oi_1
X_2237_ _1654_ _1650_ net735 VPWR VGND sg13g2_nand2_2
XFILLER_39_886 VPWR VGND sg13g2_decap_8
XFILLER_38_352 VPWR VGND sg13g2_fill_2
X_2168_ _1491_ _1555_ _1585_ VPWR VGND sg13g2_nor2_2
XFILLER_14_709 VPWR VGND sg13g2_decap_8
X_2099_ VPWR _1517_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[1\]
+ VGND sg13g2_inv_1
XFILLER_26_558 VPWR VGND sg13g2_decap_8
XFILLER_16_1017 VPWR VGND sg13g2_decap_8
XFILLER_22_753 VPWR VGND sg13g2_decap_8
XFILLER_34_591 VPWR VGND sg13g2_decap_8
XFILLER_10_926 VPWR VGND sg13g2_decap_8
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_134 VPWR VGND sg13g2_decap_4
XFILLER_1_646 VPWR VGND sg13g2_decap_8
XFILLER_45_834 VPWR VGND sg13g2_decap_8
XFILLER_28_96 VPWR VGND sg13g2_fill_2
XFILLER_17_569 VPWR VGND sg13g2_decap_8
XFILLER_32_539 VPWR VGND sg13g2_decap_8
XFILLER_13_753 VPWR VGND sg13g2_decap_8
XFILLER_40_583 VPWR VGND sg13g2_decap_8
XFILLER_9_746 VPWR VGND sg13g2_decap_8
XFILLER_12_274 VPWR VGND sg13g2_fill_1
XFILLER_5_996 VPWR VGND sg13g2_decap_8
XFILLER_4_473 VPWR VGND sg13g2_decap_8
X_3140_ _0620_ VPWR _0056_ VGND net570 net700 sg13g2_o21ai_1
XFILLER_48_661 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_fill_1
X_3071_ _0568_ net772 net709 VPWR VGND sg13g2_xnor2_1
XFILLER_36_834 VPWR VGND sg13g2_decap_8
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
X_3973_ net801 net802 _1339_ _1349_ VPWR VGND sg13g2_nor3_2
X_2924_ _0426_ net704 _0424_ _0425_ VPWR VGND sg13g2_and3_1
XFILLER_31_572 VPWR VGND sg13g2_decap_8
X_2855_ _2016_ _0339_ _0359_ VPWR VGND sg13g2_nor2_2
Xclk_div_param_inst__1__1 VPWR net35 clknet_1_1__leaf_clk_div_out VGND sg13g2_inv_1
X_2786_ _0304_ net576 VPWR VGND _1953_ sg13g2_nand2b_2
Xfanout714 net715 net714 VPWR VGND sg13g2_buf_8
Xfanout703 _0320_ net703 VPWR VGND sg13g2_buf_8
X_3407_ VGND VPWR net9 _0875_ _0878_ _0732_ sg13g2_a21oi_1
Xfanout736 _1610_ net736 VPWR VGND sg13g2_buf_8
Xfanout725 _1613_ net725 VPWR VGND sg13g2_buf_8
Xfanout758 sap_3_inst.controller_inst.opcode\[5\] net758 VPWR VGND sg13g2_buf_8
Xfanout747 sap_3_inst.controller_inst.stage\[0\] net747 VPWR VGND sg13g2_buf_8
X_3338_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[3\] net639 _0809_
+ VPWR VGND sg13g2_and2_1
Xfanout769 sap_3_inst.controller_inst.opcode\[1\] net769 VPWR VGND sg13g2_buf_1
X_3269_ _1556_ _1870_ _0328_ _0739_ _0740_ VPWR VGND sg13g2_nor4_1
XFILLER_27_812 VPWR VGND sg13g2_decap_8
XFILLER_39_683 VPWR VGND sg13g2_decap_8
XFILLER_14_506 VPWR VGND sg13g2_decap_8
XFILLER_27_889 VPWR VGND sg13g2_decap_8
XFILLER_22_550 VPWR VGND sg13g2_decap_8
XFILLER_10_723 VPWR VGND sg13g2_decap_8
XFILLER_2_911 VPWR VGND sg13g2_decap_8
XFILLER_2_988 VPWR VGND sg13g2_decap_8
XFILLER_49_447 VPWR VGND sg13g2_decap_8
XFILLER_36_108 VPWR VGND sg13g2_fill_1
XFILLER_45_631 VPWR VGND sg13g2_decap_8
XFILLER_18_823 VPWR VGND sg13g2_decap_8
XFILLER_17_344 VPWR VGND sg13g2_fill_2
XFILLER_33_848 VPWR VGND sg13g2_decap_8
XFILLER_13_550 VPWR VGND sg13g2_decap_8
XFILLER_9_543 VPWR VGND sg13g2_decap_8
X_2640_ _2045_ _2046_ _2047_ _2048_ _2049_ VPWR VGND sg13g2_and4_1
X_2571_ _1982_ _1980_ _1981_ _1884_ net5 VPWR VGND sg13g2_a22oi_1
XFILLER_5_793 VPWR VGND sg13g2_decap_8
X_4310_ net835 VGND VPWR _0167_ sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[6\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_1
X_4241_ net828 VGND VPWR _0098_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[0\]
+ clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_4172_ net805 VGND VPWR _0029_ sap_3_inst.alu_flags\[4\] net44 sg13g2_dfrbpq_1
X_3123_ _0610_ _0608_ _0611_ VPWR VGND sg13g2_nor2b_1
X_3054_ _0547_ _0522_ _0552_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_119 VPWR VGND sg13g2_decap_4
XFILLER_36_631 VPWR VGND sg13g2_decap_8
XFILLER_24_815 VPWR VGND sg13g2_decap_8
XFILLER_35_163 VPWR VGND sg13g2_fill_1
XFILLER_11_509 VPWR VGND sg13g2_decap_8
X_3956_ VGND VPWR _1326_ _1328_ _1333_ _1332_ sg13g2_a21oi_1
X_2907_ _0406_ _0408_ _0409_ VPWR VGND sg13g2_nor2_1
X_3887_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[4\] _1160_ net672
+ _0142_ VPWR VGND sg13g2_mux2_1
X_2838_ sap_3_inst.alu_inst.tmp\[0\] net792 _0342_ VPWR VGND sg13g2_xor2_1
X_2769_ _0295_ _1578_ _0296_ VPWR VGND _0294_ sg13g2_nand3b_1
XFILLER_47_907 VPWR VGND sg13g2_decap_8
Xfanout599 _0340_ net599 VPWR VGND sg13g2_buf_8
XFILLER_19_609 VPWR VGND sg13g2_decap_8
Xfanout588 _0858_ net588 VPWR VGND sg13g2_buf_8
Xfanout577 _1721_ net577 VPWR VGND sg13g2_buf_1
XFILLER_39_480 VPWR VGND sg13g2_decap_8
XFILLER_15_826 VPWR VGND sg13g2_decap_8
XFILLER_27_686 VPWR VGND sg13g2_decap_8
XFILLER_14_314 VPWR VGND sg13g2_fill_2
XFILLER_14_347 VPWR VGND sg13g2_fill_1
XFILLER_42_667 VPWR VGND sg13g2_decap_8
XFILLER_10_520 VPWR VGND sg13g2_decap_8
XFILLER_22_391 VPWR VGND sg13g2_fill_1
XFILLER_6_568 VPWR VGND sg13g2_decap_8
XFILLER_10_597 VPWR VGND sg13g2_decap_8
XFILLER_29_1027 VPWR VGND sg13g2_fill_2
XFILLER_2_785 VPWR VGND sg13g2_decap_8
XFILLER_18_620 VPWR VGND sg13g2_decap_8
XFILLER_46_951 VPWR VGND sg13g2_decap_8
XFILLER_17_141 VPWR VGND sg13g2_fill_2
XFILLER_18_697 VPWR VGND sg13g2_decap_8
XFILLER_33_645 VPWR VGND sg13g2_decap_8
XFILLER_36_1009 VPWR VGND sg13g2_decap_8
XFILLER_21_818 VPWR VGND sg13g2_decap_8
X_3810_ _1228_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[5\] net658
+ VPWR VGND sg13g2_nand2_1
XFILLER_14_870 VPWR VGND sg13g2_decap_8
X_3741_ _0732_ net603 _1178_ VPWR VGND sg13g2_nor2_1
X_3672_ net636 _1118_ _1122_ _1123_ VPWR VGND sg13g2_nor3_1
X_2623_ _2032_ net615 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[1\]
+ net617 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[1\] VPWR VGND sg13g2_a22oi_1
X_2554_ _1954_ _1957_ _1958_ _1967_ VGND VPWR _1966_ sg13g2_nor4_2
XFILLER_49_0 VPWR VGND sg13g2_decap_4
XFILLER_5_590 VPWR VGND sg13g2_decap_8
X_2485_ net752 _1636_ _1693_ _1902_ VPWR VGND sg13g2_nor3_2
X_4224_ net814 VGND VPWR _0081_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[7\]
+ clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_29_929 VPWR VGND sg13g2_decap_8
X_3106_ _0597_ VPWR _0045_ VGND _1509_ net706 sg13g2_o21ai_1
X_4086_ VGND VPWR _1525_ net579 _0177_ _1445_ sg13g2_a21oi_1
X_3037_ _0535_ net775 net708 VPWR VGND sg13g2_xnor2_1
XFILLER_24_612 VPWR VGND sg13g2_decap_8
XFILLER_36_450 VPWR VGND sg13g2_fill_1
XFILLER_12_807 VPWR VGND sg13g2_decap_8
XFILLER_24_689 VPWR VGND sg13g2_decap_8
XFILLER_20_840 VPWR VGND sg13g2_decap_8
X_3939_ VGND VPWR net803 _0155_ _0156_ _1319_ sg13g2_a21oi_1
XFILLER_47_704 VPWR VGND sg13g2_decap_8
Xclkbuf_5_7__f_sap_3_inst.alu_inst.clk_regs clknet_4_3_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_28_995 VPWR VGND sg13g2_decap_8
XFILLER_15_623 VPWR VGND sg13g2_decap_8
XFILLER_27_483 VPWR VGND sg13g2_decap_8
XFILLER_43_976 VPWR VGND sg13g2_decap_8
XFILLER_42_464 VPWR VGND sg13g2_decap_8
XFILLER_30_637 VPWR VGND sg13g2_decap_8
XFILLER_7_800 VPWR VGND sg13g2_decap_8
XFILLER_11_873 VPWR VGND sg13g2_decap_8
XFILLER_7_877 VPWR VGND sg13g2_decap_8
XFILLER_6_387 VPWR VGND sg13g2_fill_1
X_2270_ _1687_ _1630_ _1670_ VPWR VGND sg13g2_nand2_1
XFILLER_2_582 VPWR VGND sg13g2_decap_8
XFILLER_42_1024 VPWR VGND sg13g2_decap_4
XFILLER_38_748 VPWR VGND sg13g2_decap_8
XFILLER_19_973 VPWR VGND sg13g2_decap_8
XFILLER_18_494 VPWR VGND sg13g2_decap_8
XFILLER_34_976 VPWR VGND sg13g2_decap_8
XFILLER_21_615 VPWR VGND sg13g2_decap_8
X_3724_ _1146_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[7\] _1163_
+ _0097_ VPWR VGND sg13g2_a21o_1
X_3655_ _1108_ net637 _0919_ VPWR VGND sg13g2_nand2_1
X_2606_ VGND VPWR net762 _1996_ _2015_ _2014_ sg13g2_a21oi_1
X_3586_ VGND VPWR net24 net606 _1050_ _1049_ sg13g2_a21oi_1
X_2537_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[5\] net632
+ _1860_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[5\] _1950_ _1859_
+ sg13g2_a221oi_1
X_2468_ _1569_ _1617_ _1723_ _1885_ VPWR VGND sg13g2_nor3_1
X_4207_ net808 VGND VPWR _0064_ sap_3_inst.controller_inst.opcode\[6\] clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_2399_ _1816_ _1703_ _1814_ VPWR VGND sg13g2_nand2b_1
XFILLER_29_726 VPWR VGND sg13g2_decap_8
X_4138_ VPWR _0192_ _1483_ VGND sg13g2_inv_1
XFILLER_44_729 VPWR VGND sg13g2_decap_8
X_4069_ _1433_ VPWR _0172_ VGND net646 _1159_ sg13g2_o21ai_1
XFILLER_12_604 VPWR VGND sg13g2_decap_8
XFILLER_19_1015 VPWR VGND sg13g2_decap_8
XFILLER_25_954 VPWR VGND sg13g2_decap_8
XFILLER_24_486 VPWR VGND sg13g2_decap_8
XFILLER_40_968 VPWR VGND sg13g2_decap_8
XFILLER_8_619 VPWR VGND sg13g2_decap_8
XFILLER_4_858 VPWR VGND sg13g2_decap_8
XFILLER_3_324 VPWR VGND sg13g2_fill_2
XFILLER_47_501 VPWR VGND sg13g2_decap_8
XFILLER_47_578 VPWR VGND sg13g2_decap_8
XFILLER_35_729 VPWR VGND sg13g2_decap_8
XFILLER_27_280 VPWR VGND sg13g2_fill_1
XFILLER_28_792 VPWR VGND sg13g2_decap_8
XFILLER_16_954 VPWR VGND sg13g2_decap_8
XFILLER_43_773 VPWR VGND sg13g2_decap_8
XFILLER_15_497 VPWR VGND sg13g2_decap_8
XFILLER_31_957 VPWR VGND sg13g2_decap_8
XFILLER_11_670 VPWR VGND sg13g2_decap_8
XFILLER_7_674 VPWR VGND sg13g2_decap_8
X_3440_ _0909_ net662 _0907_ _0908_ VPWR VGND sg13g2_and3_1
X_3371_ _1519_ _0667_ net689 _0842_ VPWR VGND sg13g2_nor3_1
X_2322_ _1677_ _1701_ _1734_ _1737_ _1739_ VPWR VGND sg13g2_nor4_1
X_2253_ _1670_ net730 _1669_ VPWR VGND sg13g2_nand2_2
X_2184_ _1598_ _1600_ _1601_ VPWR VGND sg13g2_nor2b_2
XFILLER_38_545 VPWR VGND sg13g2_decap_8
XFILLER_19_770 VPWR VGND sg13g2_decap_8
XFILLER_22_935 VPWR VGND sg13g2_decap_8
XFILLER_34_773 VPWR VGND sg13g2_decap_8
XFILLER_21_489 VPWR VGND sg13g2_decap_8
X_3707_ _1153_ _1151_ _1152_ net582 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[1\]
+ VPWR VGND sg13g2_a22oi_1
X_3638_ net584 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[7\] _1093_
+ _0081_ VPWR VGND sg13g2_a21o_1
X_3569_ VGND VPWR _1539_ net597 _0072_ _1033_ sg13g2_a21oi_1
XFILLER_1_828 VPWR VGND sg13g2_decap_8
XFILLER_0_338 VPWR VGND sg13g2_fill_1
XFILLER_29_523 VPWR VGND sg13g2_decap_8
XFILLER_44_526 VPWR VGND sg13g2_decap_8
XFILLER_25_751 VPWR VGND sg13g2_decap_8
XFILLER_13_935 VPWR VGND sg13g2_decap_8
XFILLER_40_765 VPWR VGND sg13g2_decap_8
XFILLER_9_928 VPWR VGND sg13g2_decap_8
XFILLER_12_478 VPWR VGND sg13g2_decap_8
XFILLER_32_1001 VPWR VGND sg13g2_decap_8
XFILLER_4_655 VPWR VGND sg13g2_decap_8
XFILLER_3_121 VPWR VGND sg13g2_fill_1
XFILLER_0_861 VPWR VGND sg13g2_decap_8
XFILLER_48_843 VPWR VGND sg13g2_decap_8
Xhold5 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[6\] VPWR VGND net52
+ sg13g2_dlygate4sd3_1
XFILLER_47_375 VPWR VGND sg13g2_decap_8
XFILLER_35_526 VPWR VGND sg13g2_decap_8
XFILLER_16_751 VPWR VGND sg13g2_decap_8
XFILLER_43_570 VPWR VGND sg13g2_decap_8
X_2940_ sap_3_inst.alu_inst.tmp\[2\] net787 _0441_ VPWR VGND sg13g2_nor2b_1
X_2871_ sap_3_inst.alu_inst.tmp\[1\] net789 _0374_ VPWR VGND sg13g2_xor2_1
XFILLER_31_754 VPWR VGND sg13g2_decap_8
XFILLER_8_983 VPWR VGND sg13g2_decap_8
X_3423_ _0780_ _0852_ _0892_ _0893_ VPWR VGND sg13g2_or3_1
X_3354_ _0815_ _0816_ _0819_ _0825_ VGND VPWR _0824_ sg13g2_nor4_2
X_2305_ _1554_ _1611_ _1722_ VPWR VGND sg13g2_nor2_1
X_3285_ _0756_ net662 _0752_ _0755_ VPWR VGND sg13g2_and3_1
X_2236_ _1649_ _1651_ _1653_ VPWR VGND sg13g2_nor2_2
XFILLER_39_865 VPWR VGND sg13g2_decap_8
X_2167_ net746 net747 _1584_ VPWR VGND sg13g2_nor2b_2
XFILLER_26_537 VPWR VGND sg13g2_decap_8
X_2098_ VPWR _1516_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[1\]
+ VGND sg13g2_inv_1
XFILLER_34_570 VPWR VGND sg13g2_decap_8
XFILLER_22_732 VPWR VGND sg13g2_decap_8
XFILLER_10_905 VPWR VGND sg13g2_decap_8
Xclkbuf_regs_0_clk_div_two sap_3_inst.alu_inst.clk sap_3_inst.alu_inst.clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_1_625 VPWR VGND sg13g2_decap_8
XFILLER_49_629 VPWR VGND sg13g2_decap_8
XFILLER_45_813 VPWR VGND sg13g2_decap_8
XFILLER_28_42 VPWR VGND sg13g2_fill_1
XFILLER_17_548 VPWR VGND sg13g2_decap_8
XFILLER_44_378 VPWR VGND sg13g2_decap_4
XFILLER_44_367 VPWR VGND sg13g2_decap_4
XFILLER_32_518 VPWR VGND sg13g2_decap_8
XFILLER_13_732 VPWR VGND sg13g2_decap_8
XFILLER_40_562 VPWR VGND sg13g2_decap_8
XFILLER_9_725 VPWR VGND sg13g2_decap_8
XFILLER_5_975 VPWR VGND sg13g2_decap_8
XFILLER_4_452 VPWR VGND sg13g2_decap_8
X_3070_ _0567_ _0534_ _0537_ VPWR VGND sg13g2_nand2_1
XFILLER_48_640 VPWR VGND sg13g2_decap_8
XFILLER_36_813 VPWR VGND sg13g2_decap_8
XFILLER_35_312 VPWR VGND sg13g2_fill_1
XFILLER_23_529 VPWR VGND sg13g2_decap_8
XFILLER_44_890 VPWR VGND sg13g2_decap_8
X_3972_ net801 net802 _1345_ _1348_ VPWR VGND sg13g2_nor3_2
X_2923_ _0387_ _0385_ _0423_ _0425_ VPWR VGND sg13g2_a21o_1
XFILLER_31_551 VPWR VGND sg13g2_decap_8
X_2854_ net748 _2018_ _0358_ VPWR VGND sg13g2_and2_1
X_2785_ net13 net576 _1969_ _1978_ VPWR VGND sg13g2_and3_2
XFILLER_8_780 VPWR VGND sg13g2_decap_8
Xfanout704 _2000_ net704 VPWR VGND sg13g2_buf_8
Xfanout715 _1664_ net715 VPWR VGND sg13g2_buf_1
X_3406_ _0877_ net31 net605 VPWR VGND sg13g2_nand2_1
Xfanout748 sap_3_inst.alu_flags\[1\] net748 VPWR VGND sg13g2_buf_8
Xfanout726 net727 net726 VPWR VGND sg13g2_buf_8
Xfanout737 _1586_ net737 VPWR VGND sg13g2_buf_8
X_3337_ _0805_ _0806_ _0804_ _0808_ VPWR VGND _0807_ sg13g2_nand4_1
Xfanout759 net761 net759 VPWR VGND sg13g2_buf_8
X_3268_ VGND VPWR _1569_ _0738_ _0739_ net741 sg13g2_a21oi_1
XFILLER_39_662 VPWR VGND sg13g2_decap_8
X_2219_ _1636_ _1603_ _1623_ VPWR VGND sg13g2_nand2_2
X_3199_ _0670_ _1649_ _1670_ VPWR VGND sg13g2_nand2_1
XFILLER_27_868 VPWR VGND sg13g2_decap_8
XFILLER_42_849 VPWR VGND sg13g2_decap_8
XFILLER_35_890 VPWR VGND sg13g2_decap_8
XFILLER_10_702 VPWR VGND sg13g2_decap_8
XFILLER_10_779 VPWR VGND sg13g2_decap_8
XFILLER_2_967 VPWR VGND sg13g2_decap_8
XFILLER_49_426 VPWR VGND sg13g2_decap_8
XFILLER_1_499 VPWR VGND sg13g2_decap_8
XFILLER_18_802 VPWR VGND sg13g2_decap_8
XFILLER_45_610 VPWR VGND sg13g2_decap_8
XFILLER_18_879 VPWR VGND sg13g2_decap_8
XFILLER_45_687 VPWR VGND sg13g2_decap_8
XFILLER_33_827 VPWR VGND sg13g2_decap_8
XFILLER_9_522 VPWR VGND sg13g2_decap_8
XFILLER_9_599 VPWR VGND sg13g2_decap_8
X_2570_ _1902_ sap_3_inst.alu_flags\[4\] _1900_ _1981_ VPWR VGND sg13g2_a21o_1
XFILLER_5_772 VPWR VGND sg13g2_decap_8
X_4240_ net814 VGND VPWR _0097_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[7\]
+ clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_4_271 VPWR VGND sg13g2_fill_1
X_4171_ net807 VGND VPWR _0004_ sap_3_inst.controller_inst.stage\[3\] net43 sg13g2_dfrbpq_1
X_3122_ VPWR VGND _0345_ _0570_ _0609_ _0571_ _0610_ _0574_ sg13g2_a221oi_1
XFILLER_49_993 VPWR VGND sg13g2_decap_8
X_3053_ _0543_ _0544_ _0541_ _0551_ VPWR VGND _0550_ sg13g2_nand4_1
XFILLER_36_610 VPWR VGND sg13g2_decap_8
XFILLER_36_687 VPWR VGND sg13g2_decap_8
XFILLER_35_186 VPWR VGND sg13g2_fill_1
X_3955_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[7\] _1327_
+ _1332_ _1331_ sg13g2_a21oi_1
X_2906_ _0407_ VPWR _0408_ VGND net786 _0334_ sg13g2_o21ai_1
XFILLER_32_882 VPWR VGND sg13g2_decap_8
X_3886_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[3\] _1216_ net672
+ _0141_ VPWR VGND sg13g2_mux2_1
X_2837_ _0341_ net792 sap_3_inst.alu_inst.tmp\[0\] VPWR VGND sg13g2_nand2_1
X_2768_ net723 VPWR _0295_ VGND net742 _1568_ sg13g2_o21ai_1
X_2699_ _0230_ _0228_ _0229_ VPWR VGND sg13g2_xnor2_1
Xfanout578 net579 net578 VPWR VGND sg13g2_buf_8
Xfanout589 net591 net589 VPWR VGND sg13g2_buf_8
XFILLER_15_805 VPWR VGND sg13g2_decap_8
XFILLER_27_665 VPWR VGND sg13g2_decap_8
XFILLER_42_646 VPWR VGND sg13g2_decap_8
XFILLER_25_43 VPWR VGND sg13g2_fill_2
XFILLER_26_186 VPWR VGND sg13g2_fill_1
XFILLER_30_819 VPWR VGND sg13g2_decap_8
XFILLER_23_893 VPWR VGND sg13g2_decap_8
XFILLER_10_576 VPWR VGND sg13g2_decap_8
XFILLER_6_547 VPWR VGND sg13g2_decap_8
XFILLER_29_1006 VPWR VGND sg13g2_decap_8
XFILLER_9_0 VPWR VGND sg13g2_fill_2
XFILLER_2_764 VPWR VGND sg13g2_decap_8
XFILLER_1_274 VPWR VGND sg13g2_fill_2
XFILLER_46_930 VPWR VGND sg13g2_decap_8
XFILLER_18_676 VPWR VGND sg13g2_decap_8
XFILLER_45_484 VPWR VGND sg13g2_decap_8
XFILLER_17_175 VPWR VGND sg13g2_fill_2
XFILLER_17_186 VPWR VGND sg13g2_fill_1
XFILLER_33_624 VPWR VGND sg13g2_decap_8
X_3740_ _1177_ net594 _0917_ VPWR VGND sg13g2_nand2_1
X_3671_ VGND VPWR _1991_ _1097_ _1122_ _1121_ sg13g2_a21oi_1
XFILLER_12_1010 VPWR VGND sg13g2_decap_8
X_2622_ _2026_ _2028_ _2029_ _2030_ _2031_ VPWR VGND sg13g2_and4_1
X_2553_ VGND VPWR _1961_ _1965_ _1966_ _1720_ sg13g2_a21oi_1
X_2484_ net774 net695 _1901_ VPWR VGND sg13g2_nor2_1
X_4223_ net811 VGND VPWR _0080_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[6\]
+ clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_29_908 VPWR VGND sg13g2_decap_8
X_3105_ _0597_ sap_3_inst.out\[4\] net706 VPWR VGND sg13g2_nand2_1
X_4085_ net579 _1444_ _1445_ VPWR VGND sg13g2_nor2_1
XFILLER_49_790 VPWR VGND sg13g2_decap_8
X_3036_ _0534_ net775 net708 VPWR VGND sg13g2_nand2_1
XFILLER_37_985 VPWR VGND sg13g2_decap_8
XFILLER_24_668 VPWR VGND sg13g2_decap_8
XFILLER_23_178 VPWR VGND sg13g2_fill_2
X_3938_ net803 _1315_ _1319_ VPWR VGND sg13g2_nor2_1
X_3869_ VGND VPWR net609 _1021_ _1270_ net653 sg13g2_a21oi_1
XFILLER_20_896 VPWR VGND sg13g2_decap_8
XFILLER_3_539 VPWR VGND sg13g2_decap_8
XFILLER_4_1019 VPWR VGND sg13g2_decap_8
XFILLER_15_602 VPWR VGND sg13g2_decap_8
XFILLER_27_462 VPWR VGND sg13g2_decap_8
XFILLER_28_974 VPWR VGND sg13g2_decap_8
XFILLER_36_64 VPWR VGND sg13g2_fill_1
XFILLER_43_955 VPWR VGND sg13g2_decap_8
XFILLER_42_443 VPWR VGND sg13g2_decap_8
XFILLER_15_679 VPWR VGND sg13g2_decap_8
XFILLER_30_616 VPWR VGND sg13g2_decap_8
XFILLER_11_852 VPWR VGND sg13g2_decap_8
XFILLER_23_690 VPWR VGND sg13g2_decap_8
XFILLER_10_351 VPWR VGND sg13g2_fill_2
XFILLER_7_856 VPWR VGND sg13g2_decap_8
XFILLER_2_561 VPWR VGND sg13g2_decap_8
XFILLER_42_1003 VPWR VGND sg13g2_decap_8
XFILLER_38_727 VPWR VGND sg13g2_decap_8
XFILLER_19_952 VPWR VGND sg13g2_decap_8
XFILLER_18_473 VPWR VGND sg13g2_decap_8
XFILLER_34_955 VPWR VGND sg13g2_decap_8
XFILLER_33_498 VPWR VGND sg13g2_decap_8
X_3723_ _1090_ _1092_ net582 _1163_ VPWR VGND sg13g2_nor3_1
X_3654_ VPWR _0083_ _1107_ VGND sg13g2_inv_1
X_2605_ _1600_ _1831_ _2014_ VPWR VGND sg13g2_nor2_2
X_3585_ _0306_ net605 _1049_ VPWR VGND sg13g2_nor2_1
X_2536_ _1947_ _1948_ _1945_ _1949_ VPWR VGND sg13g2_nand3_1
X_2467_ VGND VPWR _1884_ _1883_ net718 sg13g2_or2_1
X_4206_ net804 VGND VPWR _0063_ sap_3_inst.controller_inst.opcode\[5\] clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
X_2398_ _1814_ _1703_ _1815_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_705 VPWR VGND sg13g2_decap_8
X_4137_ _1483_ _1480_ net801 _1479_ net797 VPWR VGND sg13g2_a22oi_1
XFILLER_44_708 VPWR VGND sg13g2_decap_8
X_4068_ _1433_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[3\] net645
+ VPWR VGND sg13g2_nand2_1
X_3019_ VGND VPWR _0475_ _0489_ _0518_ _0473_ sg13g2_a21oi_1
XFILLER_25_933 VPWR VGND sg13g2_decap_8
XFILLER_37_782 VPWR VGND sg13g2_decap_8
XFILLER_24_465 VPWR VGND sg13g2_decap_8
XFILLER_40_947 VPWR VGND sg13g2_decap_8
XFILLER_20_693 VPWR VGND sg13g2_decap_8
XFILLER_4_837 VPWR VGND sg13g2_decap_8
XFILLER_47_557 VPWR VGND sg13g2_decap_8
XFILLER_35_708 VPWR VGND sg13g2_decap_8
XFILLER_16_933 VPWR VGND sg13g2_decap_8
XFILLER_28_771 VPWR VGND sg13g2_decap_8
XFILLER_34_218 VPWR VGND sg13g2_decap_4
XFILLER_43_752 VPWR VGND sg13g2_decap_8
XFILLER_15_476 VPWR VGND sg13g2_decap_8
XFILLER_31_936 VPWR VGND sg13g2_decap_8
XFILLER_10_170 VPWR VGND sg13g2_fill_1
XFILLER_7_653 VPWR VGND sg13g2_decap_8
XFILLER_6_174 VPWR VGND sg13g2_fill_1
X_3370_ _0837_ _0838_ _0839_ _0840_ _0841_ VPWR VGND sg13g2_and4_1
X_2321_ VGND VPWR _1629_ _1659_ _1738_ net730 sg13g2_a21oi_1
X_2252_ _1669_ net762 _1668_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_4 VPWR VGND sg13g2_fill_1
X_2183_ net765 _1570_ _1492_ _1600_ VPWR VGND sg13g2_nand3_1
XFILLER_38_524 VPWR VGND sg13g2_decap_8
XFILLER_26_719 VPWR VGND sg13g2_decap_8
XFILLER_34_752 VPWR VGND sg13g2_decap_8
XFILLER_22_914 VPWR VGND sg13g2_decap_8
XFILLER_21_468 VPWR VGND sg13g2_decap_8
X_3706_ net582 _1150_ _1152_ VPWR VGND sg13g2_nor2_1
XFILLER_30_980 VPWR VGND sg13g2_decap_8
X_3637_ net584 _1090_ _1092_ _1093_ VPWR VGND sg13g2_nor3_1
X_3568_ net597 _1024_ _1030_ _1032_ _1033_ VPWR VGND sg13g2_nor4_1
XFILLER_1_807 VPWR VGND sg13g2_decap_8
X_2519_ _1934_ net624 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[6\]
+ net631 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[6\] VPWR VGND sg13g2_a22oi_1
X_3499_ _0964_ _0965_ _0963_ _0966_ VPWR VGND sg13g2_nand3_1
XFILLER_29_502 VPWR VGND sg13g2_decap_8
XFILLER_44_505 VPWR VGND sg13g2_decap_8
XFILLER_29_579 VPWR VGND sg13g2_decap_8
XFILLER_25_730 VPWR VGND sg13g2_decap_8
XFILLER_13_914 VPWR VGND sg13g2_decap_8
XFILLER_40_744 VPWR VGND sg13g2_decap_8
XFILLER_9_907 VPWR VGND sg13g2_decap_8
XFILLER_33_98 VPWR VGND sg13g2_fill_2
XFILLER_20_490 VPWR VGND sg13g2_decap_8
XFILLER_4_634 VPWR VGND sg13g2_decap_8
XFILLER_3_100 VPWR VGND sg13g2_fill_1
XFILLER_0_840 VPWR VGND sg13g2_decap_8
XFILLER_48_822 VPWR VGND sg13g2_decap_8
Xhold6 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[7\] VPWR VGND net53
+ sg13g2_dlygate4sd3_1
XFILLER_47_354 VPWR VGND sg13g2_decap_8
XFILLER_35_505 VPWR VGND sg13g2_decap_8
XFILLER_48_899 VPWR VGND sg13g2_decap_8
XFILLER_16_730 VPWR VGND sg13g2_decap_8
X_2870_ _0373_ net789 sap_3_inst.alu_inst.tmp\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_15_295 VPWR VGND sg13g2_fill_1
XFILLER_31_733 VPWR VGND sg13g2_decap_8
XFILLER_8_962 VPWR VGND sg13g2_decap_8
XFILLER_7_461 VPWR VGND sg13g2_decap_4
X_3422_ VGND VPWR _0892_ _0891_ _0770_ sg13g2_or2_1
X_3353_ _0820_ _0821_ _0822_ _0823_ _0824_ VPWR VGND sg13g2_or4_1
X_2304_ VPWR _1721_ _1720_ VGND sg13g2_inv_1
X_3284_ _0755_ net677 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[0\]
+ net688 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2235_ _1575_ _1604_ _1641_ _1652_ VPWR VGND sg13g2_or3_1
XFILLER_39_844 VPWR VGND sg13g2_decap_8
X_2166_ _1583_ net743 _1580_ VPWR VGND sg13g2_nand2_2
XFILLER_26_516 VPWR VGND sg13g2_decap_8
XFILLER_0_1022 VPWR VGND sg13g2_decap_8
X_2097_ VPWR _1515_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[1\]
+ VGND sg13g2_inv_1
XFILLER_22_711 VPWR VGND sg13g2_decap_8
X_2999_ VGND VPWR sap_3_inst.alu_inst.act\[4\] net702 _0499_ net693 sg13g2_a21oi_1
XFILLER_22_788 VPWR VGND sg13g2_decap_8
XFILLER_1_604 VPWR VGND sg13g2_decap_8
XFILLER_49_608 VPWR VGND sg13g2_decap_8
XFILLER_29_354 VPWR VGND sg13g2_fill_2
XFILLER_17_527 VPWR VGND sg13g2_decap_8
XFILLER_45_869 VPWR VGND sg13g2_decap_8
XFILLER_13_711 VPWR VGND sg13g2_decap_8
XFILLER_40_541 VPWR VGND sg13g2_decap_8
XFILLER_9_704 VPWR VGND sg13g2_decap_8
XFILLER_13_788 VPWR VGND sg13g2_decap_8
XFILLER_5_954 VPWR VGND sg13g2_decap_8
XFILLER_5_47 VPWR VGND sg13g2_fill_1
XFILLER_48_696 VPWR VGND sg13g2_decap_8
XFILLER_39_1019 VPWR VGND sg13g2_decap_8
XFILLER_36_869 VPWR VGND sg13g2_decap_8
X_3971_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[0\] sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[1\]
+ _1335_ _1347_ VPWR VGND sg13g2_nor3_2
XFILLER_23_508 VPWR VGND sg13g2_decap_8
X_2922_ _0387_ _0423_ _0385_ _0424_ VPWR VGND sg13g2_nand3_1
XFILLER_31_530 VPWR VGND sg13g2_decap_8
X_2853_ _2017_ _0339_ _0357_ VPWR VGND sg13g2_nor2_1
X_2784_ VPWR net12 _0303_ VGND sg13g2_inv_1
Xfanout705 _0274_ net705 VPWR VGND sg13g2_buf_8
X_3405_ _0876_ net664 net668 VPWR VGND sg13g2_nand2b_1
Xfanout727 _1583_ net727 VPWR VGND sg13g2_buf_8
Xfanout749 _1625_ net749 VPWR VGND sg13g2_buf_2
Xfanout716 _1601_ net716 VPWR VGND sg13g2_buf_8
Xfanout738 _1584_ net738 VPWR VGND sg13g2_buf_8
X_3336_ _0807_ net677 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[3\]
+ net682 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[3\] VPWR VGND sg13g2_a22oi_1
X_3267_ VGND VPWR _0738_ _0737_ _0643_ sg13g2_or2_1
XFILLER_22_1012 VPWR VGND sg13g2_decap_8
XFILLER_39_641 VPWR VGND sg13g2_decap_8
X_3198_ net714 net705 _0630_ _0631_ _0669_ VPWR VGND sg13g2_and4_1
X_2218_ _1604_ _1624_ _1635_ VPWR VGND sg13g2_nor2_2
XFILLER_38_140 VPWR VGND sg13g2_fill_1
X_2149_ net751 net750 _1566_ VPWR VGND sg13g2_nor2_1
XFILLER_26_324 VPWR VGND sg13g2_decap_8
XFILLER_27_847 VPWR VGND sg13g2_decap_8
XFILLER_42_828 VPWR VGND sg13g2_decap_8
XFILLER_22_585 VPWR VGND sg13g2_decap_8
XFILLER_10_758 VPWR VGND sg13g2_decap_8
XFILLER_6_729 VPWR VGND sg13g2_decap_8
XFILLER_2_946 VPWR VGND sg13g2_decap_8
XFILLER_49_405 VPWR VGND sg13g2_decap_8
XFILLER_7_1017 VPWR VGND sg13g2_decap_8
XFILLER_39_31 VPWR VGND sg13g2_fill_2
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_478 VPWR VGND sg13g2_decap_8
XFILLER_18_858 VPWR VGND sg13g2_decap_8
XFILLER_45_666 VPWR VGND sg13g2_decap_8
XFILLER_33_806 VPWR VGND sg13g2_decap_8
XFILLER_26_880 VPWR VGND sg13g2_decap_8
XFILLER_9_501 VPWR VGND sg13g2_decap_8
XFILLER_41_894 VPWR VGND sg13g2_decap_8
XFILLER_13_585 VPWR VGND sg13g2_decap_8
XFILLER_9_578 VPWR VGND sg13g2_decap_8
XFILLER_5_751 VPWR VGND sg13g2_decap_8
XFILLER_4_261 VPWR VGND sg13g2_fill_1
XFILLER_45_1023 VPWR VGND sg13g2_decap_4
X_4170_ net807 VGND VPWR _0003_ sap_3_inst.controller_inst.stage\[2\] net42 sg13g2_dfrbpq_2
X_3121_ _0609_ _2022_ _0351_ VPWR VGND sg13g2_nand2_1
XFILLER_49_972 VPWR VGND sg13g2_decap_8
X_3052_ VGND VPWR _0347_ _0547_ _0550_ _0549_ sg13g2_a21oi_1
XFILLER_48_493 VPWR VGND sg13g2_decap_8
XFILLER_36_666 VPWR VGND sg13g2_decap_8
XFILLER_17_891 VPWR VGND sg13g2_decap_8
XFILLER_32_861 VPWR VGND sg13g2_decap_8
X_3954_ sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[2\] VPWR _1331_ VGND
+ sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[1\] _1330_ sg13g2_o21ai_1
X_2905_ _0361_ VPWR _0407_ VGND net787 sap_3_inst.alu_inst.tmp\[2\] sg13g2_o21ai_1
X_3885_ VPWR _0140_ _1281_ VGND sg13g2_inv_1
X_2836_ _0340_ _0332_ _0338_ VPWR VGND sg13g2_nand2_2
X_2767_ net742 net739 _0292_ _0293_ _0294_ VPWR VGND sg13g2_nor4_1
X_2698_ net782 net780 _0229_ VPWR VGND sg13g2_xor2_1
Xfanout579 _1442_ net579 VPWR VGND sg13g2_buf_8
X_3319_ _0790_ net669 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[5\]
+ net672 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4299_ net834 VGND VPWR _0156_ sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[0\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_46_419 VPWR VGND sg13g2_decap_8
XFILLER_27_644 VPWR VGND sg13g2_decap_8
XFILLER_26_154 VPWR VGND sg13g2_fill_2
XFILLER_42_625 VPWR VGND sg13g2_decap_8
XFILLER_23_872 VPWR VGND sg13g2_decap_8
XFILLER_41_54 VPWR VGND sg13g2_fill_1
XFILLER_6_526 VPWR VGND sg13g2_decap_8
XFILLER_10_555 VPWR VGND sg13g2_decap_8
XFILLER_2_743 VPWR VGND sg13g2_decap_8
XFILLER_49_257 VPWR VGND sg13g2_decap_8
XFILLER_38_909 VPWR VGND sg13g2_decap_8
XFILLER_46_986 VPWR VGND sg13g2_decap_8
XFILLER_45_463 VPWR VGND sg13g2_decap_8
XFILLER_18_655 VPWR VGND sg13g2_decap_8
XFILLER_33_603 VPWR VGND sg13g2_decap_8
XFILLER_41_691 VPWR VGND sg13g2_decap_8
X_3670_ net13 _1097_ _1121_ VPWR VGND sg13g2_nor2_1
X_2621_ _2030_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[1\] net619
+ VPWR VGND sg13g2_nand2_1
X_2552_ _1857_ _1960_ _1963_ _1964_ _1965_ VPWR VGND sg13g2_and4_1
X_4222_ net830 VGND VPWR _0079_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[5\]
+ clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_2483_ _1900_ net695 VPWR VGND sg13g2_inv_2
X_3104_ net783 sap_3_inst.out\[3\] net705 _0044_ VPWR VGND sg13g2_mux2_1
X_4084_ VGND VPWR _0343_ net698 _1444_ _1443_ sg13g2_a21oi_1
X_3035_ net598 net779 _0533_ _0038_ VPWR VGND sg13g2_a21o_1
XFILLER_48_290 VPWR VGND sg13g2_decap_8
XFILLER_37_964 VPWR VGND sg13g2_decap_8
XFILLER_24_647 VPWR VGND sg13g2_decap_8
X_3937_ _0155_ _1314_ _1318_ VPWR VGND sg13g2_nand2_2
X_3868_ net586 _1083_ _0305_ _1269_ VPWR VGND sg13g2_nand3_1
XFILLER_20_875 VPWR VGND sg13g2_decap_8
X_2819_ _1662_ VPWR _0323_ VGND _1558_ _1628_ sg13g2_o21ai_1
X_3799_ VPWR _0114_ _1221_ VGND sg13g2_inv_1
XFILLER_3_518 VPWR VGND sg13g2_decap_8
XFILLER_47_739 VPWR VGND sg13g2_decap_8
XFILLER_28_953 VPWR VGND sg13g2_decap_8
XFILLER_27_441 VPWR VGND sg13g2_decap_8
XFILLER_43_934 VPWR VGND sg13g2_decap_8
XFILLER_42_433 VPWR VGND sg13g2_fill_1
XFILLER_14_146 VPWR VGND sg13g2_fill_1
XFILLER_15_658 VPWR VGND sg13g2_decap_8
XFILLER_42_499 VPWR VGND sg13g2_decap_8
XFILLER_11_831 VPWR VGND sg13g2_decap_8
XFILLER_7_835 VPWR VGND sg13g2_decap_8
XFILLER_2_540 VPWR VGND sg13g2_decap_8
XFILLER_38_706 VPWR VGND sg13g2_decap_8
XFILLER_19_931 VPWR VGND sg13g2_decap_8
XFILLER_46_783 VPWR VGND sg13g2_decap_8
XFILLER_34_934 VPWR VGND sg13g2_decap_8
X_3722_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[6\] _1162_ _1147_
+ _0096_ VPWR VGND sg13g2_mux2_1
X_3653_ _1107_ _1103_ _1106_ net636 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[1\]
+ VPWR VGND sg13g2_a22oi_1
X_2604_ _2013_ _2004_ _2007_ VPWR VGND sg13g2_nand2_2
XFILLER_6_890 VPWR VGND sg13g2_decap_8
X_3584_ _1045_ _1047_ net660 _1048_ VPWR VGND sg13g2_mux2_1
X_2535_ _1948_ net625 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[5\]
+ net628 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[5\] VPWR VGND sg13g2_a22oi_1
X_2466_ VGND VPWR _1881_ _1882_ _1883_ _1870_ sg13g2_a21oi_1
X_4205_ net804 VGND VPWR _0062_ sap_3_inst.controller_inst.opcode\[4\] clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4136_ VPWR _0191_ _1482_ VGND sg13g2_inv_1
X_2397_ _1814_ net736 _1553_ _1580_ net743 VPWR VGND sg13g2_a22oi_1
X_4067_ net645 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[2\] _1432_
+ _0171_ VPWR VGND sg13g2_a21o_1
XFILLER_37_761 VPWR VGND sg13g2_decap_8
X_3018_ VGND VPWR _0347_ _0515_ _0517_ _0516_ sg13g2_a21oi_1
XFILLER_25_912 VPWR VGND sg13g2_decap_8
XFILLER_24_444 VPWR VGND sg13g2_decap_8
XFILLER_40_926 VPWR VGND sg13g2_decap_8
XFILLER_25_989 VPWR VGND sg13g2_decap_8
XFILLER_12_639 VPWR VGND sg13g2_decap_8
XFILLER_20_672 VPWR VGND sg13g2_decap_8
XFILLER_4_816 VPWR VGND sg13g2_decap_8
XFILLER_47_536 VPWR VGND sg13g2_decap_8
XFILLER_28_750 VPWR VGND sg13g2_decap_8
XFILLER_16_912 VPWR VGND sg13g2_decap_8
XFILLER_43_731 VPWR VGND sg13g2_decap_8
XFILLER_16_989 VPWR VGND sg13g2_decap_8
XFILLER_31_915 VPWR VGND sg13g2_decap_8
XFILLER_7_632 VPWR VGND sg13g2_decap_8
XFILLER_3_882 VPWR VGND sg13g2_decap_8
X_2320_ net735 _1736_ _1737_ VPWR VGND sg13g2_nor2_1
X_2251_ net757 sap_3_inst.alu_flags\[0\] sap_3_inst.alu_flags\[2\] net748 sap_3_inst.alu_flags\[3\]
+ net760 _1668_ VPWR VGND sg13g2_mux4_1
XFILLER_38_503 VPWR VGND sg13g2_decap_8
X_2182_ _1599_ _1594_ _1597_ VPWR VGND sg13g2_nand2_1
XFILLER_46_580 VPWR VGND sg13g2_decap_8
XFILLER_34_731 VPWR VGND sg13g2_decap_8
XFILLER_33_252 VPWR VGND sg13g2_fill_2
X_3705_ _1151_ net607 _0883_ VPWR VGND sg13g2_nand2_1
X_3636_ _1092_ _1091_ VPWR VGND sg13g2_inv_2
X_3567_ VGND VPWR net570 net605 _1032_ _1031_ sg13g2_a21oi_1
X_2518_ _1933_ net614 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[6\]
+ net600 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[6\] VPWR VGND sg13g2_a22oi_1
X_3498_ _0965_ net669 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[4\]
+ net641 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_25_1010 VPWR VGND sg13g2_decap_8
X_2449_ _1861_ _1863_ _1858_ _1866_ VPWR VGND _1865_ sg13g2_nand4_1
X_4119_ _1470_ net800 u_ser.shadow_reg\[6\] VPWR VGND sg13g2_nand2b_1
XFILLER_17_709 VPWR VGND sg13g2_decap_8
XFILLER_29_558 VPWR VGND sg13g2_decap_8
XFILLER_12_403 VPWR VGND sg13g2_fill_1
XFILLER_25_786 VPWR VGND sg13g2_decap_8
XFILLER_40_723 VPWR VGND sg13g2_decap_8
XFILLER_33_88 VPWR VGND sg13g2_fill_2
XFILLER_4_613 VPWR VGND sg13g2_decap_8
XFILLER_3_178 VPWR VGND sg13g2_fill_1
XFILLER_3_156 VPWR VGND sg13g2_fill_1
XFILLER_48_801 VPWR VGND sg13g2_decap_8
XFILLER_0_896 VPWR VGND sg13g2_decap_8
Xhold7 sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[1\] VPWR VGND net54
+ sg13g2_dlygate4sd3_1
XFILLER_48_878 VPWR VGND sg13g2_decap_8
XFILLER_47_333 VPWR VGND sg13g2_decap_8
XFILLER_16_786 VPWR VGND sg13g2_decap_8
XFILLER_31_712 VPWR VGND sg13g2_decap_8
XFILLER_8_941 VPWR VGND sg13g2_decap_8
XFILLER_31_789 VPWR VGND sg13g2_decap_8
X_3421_ _0891_ _0888_ _0890_ net665 _1510_ VPWR VGND sg13g2_a22oi_1
X_3352_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[0\] net670 _0823_
+ VPWR VGND sg13g2_and2_1
X_2303_ _1556_ _1719_ _1720_ VPWR VGND sg13g2_nor2_2
X_3283_ _0754_ _0666_ _0707_ VPWR VGND sg13g2_nand2_1
X_2234_ _1575_ _1604_ _1641_ _1651_ VPWR VGND sg13g2_nor3_2
XFILLER_39_823 VPWR VGND sg13g2_decap_8
X_2165_ _1552_ _1581_ _1582_ VPWR VGND sg13g2_nor2_2
XFILLER_0_1001 VPWR VGND sg13g2_decap_8
X_2096_ VPWR _1514_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[1\]
+ VGND sg13g2_inv_1
XFILLER_41_509 VPWR VGND sg13g2_decap_8
XFILLER_0_81 VPWR VGND sg13g2_decap_4
XFILLER_21_222 VPWR VGND sg13g2_fill_2
XFILLER_22_767 VPWR VGND sg13g2_decap_8
X_2998_ _0498_ _0497_ net702 VPWR VGND sg13g2_nand2b_1
X_3619_ _1077_ net595 _0995_ VPWR VGND sg13g2_nand2_1
XFILLER_0_115 VPWR VGND sg13g2_fill_2
XFILLER_0_104 VPWR VGND sg13g2_decap_4
XFILLER_17_506 VPWR VGND sg13g2_decap_8
XFILLER_45_848 VPWR VGND sg13g2_decap_8
XFILLER_40_520 VPWR VGND sg13g2_decap_8
XFILLER_25_583 VPWR VGND sg13g2_decap_8
XFILLER_13_767 VPWR VGND sg13g2_decap_8
XFILLER_40_597 VPWR VGND sg13g2_decap_8
XFILLER_8_204 VPWR VGND sg13g2_fill_1
XFILLER_5_933 VPWR VGND sg13g2_decap_8
XFILLER_4_487 VPWR VGND sg13g2_decap_8
XFILLER_0_693 VPWR VGND sg13g2_decap_8
XFILLER_48_675 VPWR VGND sg13g2_decap_8
XFILLER_36_848 VPWR VGND sg13g2_decap_8
X_3970_ _1341_ _1345_ _1346_ VPWR VGND sg13g2_nor2_2
X_2921_ _0423_ net786 net709 VPWR VGND sg13g2_xnor2_1
XFILLER_16_583 VPWR VGND sg13g2_decap_8
X_2852_ net575 _0355_ _0346_ _0356_ VPWR VGND sg13g2_nand3_1
XFILLER_31_586 VPWR VGND sg13g2_decap_8
X_2783_ _0303_ net577 VPWR VGND _2068_ sg13g2_nand2b_2
X_3404_ net660 net668 _0875_ VPWR VGND sg13g2_nor2_2
Xfanout706 _0274_ net706 VPWR VGND sg13g2_buf_8
Xfanout728 net729 net728 VPWR VGND sg13g2_buf_8
Xfanout739 _1568_ net739 VPWR VGND sg13g2_buf_8
Xfanout717 net718 net717 VPWR VGND sg13g2_buf_8
X_3335_ _0806_ net684 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[3\]
+ net687 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[3\] VPWR VGND sg13g2_a22oi_1
X_3266_ _0319_ _0736_ _0737_ VPWR VGND sg13g2_nor2_1
XFILLER_39_620 VPWR VGND sg13g2_decap_8
X_2217_ _1634_ _1587_ net736 VPWR VGND sg13g2_nand2_2
X_3197_ _0668_ net705 _0630_ VPWR VGND sg13g2_nand2_1
XFILLER_27_826 VPWR VGND sg13g2_decap_8
X_2148_ _1565_ net756 net754 VPWR VGND sg13g2_nand2b_1
XFILLER_39_697 VPWR VGND sg13g2_decap_8
XFILLER_42_807 VPWR VGND sg13g2_decap_8
X_2079_ VPWR _1497_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[3\]
+ VGND sg13g2_inv_1
XFILLER_22_564 VPWR VGND sg13g2_decap_8
XFILLER_6_708 VPWR VGND sg13g2_decap_8
XFILLER_10_737 VPWR VGND sg13g2_decap_8
XFILLER_2_925 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_fill_1
XFILLER_1_457 VPWR VGND sg13g2_decap_8
XFILLER_45_645 VPWR VGND sg13g2_decap_8
XFILLER_18_837 VPWR VGND sg13g2_decap_8
XFILLER_41_873 VPWR VGND sg13g2_decap_8
XFILLER_40_372 VPWR VGND sg13g2_fill_1
XFILLER_13_564 VPWR VGND sg13g2_decap_8
XFILLER_9_557 VPWR VGND sg13g2_decap_8
XFILLER_5_730 VPWR VGND sg13g2_decap_8
XFILLER_45_1002 VPWR VGND sg13g2_decap_8
X_3120_ _2002_ _2023_ _0608_ VPWR VGND sg13g2_nor2_1
XFILLER_49_951 VPWR VGND sg13g2_decap_8
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_48_472 VPWR VGND sg13g2_decap_8
X_3051_ _0548_ VPWR _0549_ VGND net775 _0334_ sg13g2_o21ai_1
XFILLER_36_645 VPWR VGND sg13g2_decap_8
XFILLER_24_829 VPWR VGND sg13g2_decap_8
XFILLER_17_870 VPWR VGND sg13g2_decap_8
XFILLER_32_840 VPWR VGND sg13g2_decap_8
X_3953_ _1329_ VPWR _1330_ VGND net803 sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[5\]
+ sg13g2_o21ai_1
X_2904_ _0404_ VPWR _0406_ VGND _0355_ _0405_ sg13g2_o21ai_1
X_3884_ _1281_ _1154_ _1280_ _0758_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[2\]
+ VPWR VGND sg13g2_a22oi_1
X_2835_ _0339_ _2005_ _2006_ VPWR VGND sg13g2_nand2_1
X_2766_ VGND VPWR net731 _1758_ _0293_ _1896_ sg13g2_a21oi_1
X_2697_ _0228_ net774 net777 VPWR VGND sg13g2_xnor2_1
X_3318_ _0789_ net642 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[5\]
+ net665 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[5\] VPWR VGND sg13g2_a22oi_1
Xfanout569 _1967_ net569 VPWR VGND sg13g2_buf_8
X_4298_ net834 VGND VPWR _0155_ sap_3_inst.reg_file_inst.array_serializer_inst.state\[1\]
+ clknet_3_4__leaf_clk sg13g2_dfrbpq_1
X_3249_ _0715_ _0717_ _0714_ _0720_ VPWR VGND _0718_ sg13g2_nand4_1
XFILLER_27_623 VPWR VGND sg13g2_decap_8
XFILLER_39_494 VPWR VGND sg13g2_decap_8
XFILLER_42_604 VPWR VGND sg13g2_decap_8
XFILLER_23_851 VPWR VGND sg13g2_decap_8
XFILLER_10_534 VPWR VGND sg13g2_decap_8
XFILLER_6_505 VPWR VGND sg13g2_decap_8
X_2133__2 VPWR net36 clknet_leaf_1_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
XFILLER_9_2 VPWR VGND sg13g2_fill_1
XFILLER_2_722 VPWR VGND sg13g2_decap_8
XFILLER_2_799 VPWR VGND sg13g2_decap_8
XFILLER_18_634 VPWR VGND sg13g2_decap_8
XFILLER_46_965 VPWR VGND sg13g2_decap_8
XFILLER_45_442 VPWR VGND sg13g2_decap_8
XFILLER_33_659 VPWR VGND sg13g2_decap_8
XFILLER_41_670 VPWR VGND sg13g2_decap_8
XFILLER_14_884 VPWR VGND sg13g2_decap_8
X_2620_ _2029_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[1\] net620
+ VPWR VGND sg13g2_nand2_1
X_2551_ _1964_ net601 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[5\]
+ net628 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[5\] VPWR VGND sg13g2_a22oi_1
X_2482_ VGND VPWR _1885_ _1899_ _1898_ _1569_ sg13g2_a21oi_2
X_4221_ net815 VGND VPWR _0078_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[4\]
+ clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3103_ net786 sap_3_inst.out\[2\] net705 _0043_ VPWR VGND sg13g2_mux2_1
X_4083_ net793 net698 _1443_ VPWR VGND sg13g2_nor2_1
X_3034_ VPWR VGND _0532_ net598 _0531_ net569 _0533_ _0330_ sg13g2_a221oi_1
XFILLER_37_943 VPWR VGND sg13g2_decap_8
XFILLER_24_626 VPWR VGND sg13g2_decap_8
X_3936_ _1318_ _1315_ _1317_ VPWR VGND sg13g2_nand2_1
XFILLER_20_854 VPWR VGND sg13g2_decap_8
X_3867_ net585 _1018_ _1267_ _1268_ VPWR VGND sg13g2_nor3_1
X_2818_ _0322_ net716 _1773_ VPWR VGND sg13g2_nand2b_1
X_3798_ _1221_ _0870_ _1220_ net657 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[0\]
+ VPWR VGND sg13g2_a22oi_1
X_2749_ _1690_ VPWR _0276_ VGND net731 _1692_ sg13g2_o21ai_1
XFILLER_11_36 VPWR VGND sg13g2_fill_1
XFILLER_47_718 VPWR VGND sg13g2_decap_8
XFILLER_28_932 VPWR VGND sg13g2_decap_8
XFILLER_43_913 VPWR VGND sg13g2_decap_8
XFILLER_14_125 VPWR VGND sg13g2_fill_1
XFILLER_15_637 VPWR VGND sg13g2_decap_8
XFILLER_27_497 VPWR VGND sg13g2_decap_8
XFILLER_42_478 VPWR VGND sg13g2_decap_8
Xclkbuf_5_22__f_sap_3_inst.alu_inst.clk_regs clknet_4_11_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_35_1023 VPWR VGND sg13g2_decap_4
XFILLER_11_810 VPWR VGND sg13g2_decap_8
XFILLER_7_814 VPWR VGND sg13g2_decap_8
XFILLER_11_887 VPWR VGND sg13g2_decap_8
XFILLER_2_596 VPWR VGND sg13g2_decap_8
XFILLER_19_910 VPWR VGND sg13g2_decap_8
XFILLER_46_762 VPWR VGND sg13g2_decap_8
XFILLER_45_272 VPWR VGND sg13g2_fill_2
XFILLER_19_987 VPWR VGND sg13g2_decap_8
XFILLER_34_913 VPWR VGND sg13g2_decap_8
Xclkbuf_5_11__f_sap_3_inst.alu_inst.clk_regs clknet_4_5_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_21_629 VPWR VGND sg13g2_decap_8
XFILLER_14_681 VPWR VGND sg13g2_decap_8
X_3721_ _1083_ _1085_ net570 _1162_ VPWR VGND sg13g2_nand3_1
XFILLER_9_140 VPWR VGND sg13g2_fill_1
X_3652_ VPWR VGND _1105_ net636 _1104_ net607 _1106_ _0900_ sg13g2_a221oi_1
X_2603_ _2005_ _2009_ _2012_ VPWR VGND sg13g2_nor2_2
X_3583_ _0868_ _1046_ _1047_ VPWR VGND sg13g2_nor2b_2
X_2534_ net697 net626 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[5\]
+ _1947_ VPWR VGND sg13g2_nand3_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_2465_ VGND VPWR _1592_ net723 _1882_ net741 sg13g2_a21oi_1
X_2396_ net714 _1812_ _1637_ _1813_ VPWR VGND sg13g2_nand3_1
X_4204_ net804 VGND VPWR _0061_ sap_3_inst.controller_inst.opcode\[3\] clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
X_4135_ _1482_ _1480_ net802 _1479_ net796 VPWR VGND sg13g2_a22oi_1
X_4066_ VPWR VGND _0730_ net645 _1065_ net611 _1432_ _0931_ sg13g2_a221oi_1
XFILLER_37_740 VPWR VGND sg13g2_decap_8
X_3017_ net780 _0336_ _0516_ VPWR VGND sg13g2_nor2_1
XFILLER_24_423 VPWR VGND sg13g2_decap_8
XFILLER_25_968 VPWR VGND sg13g2_decap_8
XFILLER_40_905 VPWR VGND sg13g2_decap_8
XFILLER_12_618 VPWR VGND sg13g2_decap_8
XFILLER_20_651 VPWR VGND sg13g2_decap_8
X_3919_ net643 _1124_ _1303_ _1304_ _1305_ VPWR VGND sg13g2_nor4_1
XFILLER_47_515 VPWR VGND sg13g2_decap_8
XFILLER_19_239 VPWR VGND sg13g2_fill_2
XFILLER_43_710 VPWR VGND sg13g2_decap_8
XFILLER_16_968 VPWR VGND sg13g2_decap_8
XFILLER_43_787 VPWR VGND sg13g2_decap_8
XFILLER_24_990 VPWR VGND sg13g2_decap_8
XFILLER_8_59 VPWR VGND sg13g2_fill_1
XFILLER_7_611 VPWR VGND sg13g2_decap_8
XFILLER_11_684 VPWR VGND sg13g2_decap_8
XFILLER_7_688 VPWR VGND sg13g2_decap_8
XFILLER_3_861 VPWR VGND sg13g2_decap_8
X_4153__11 VPWR net45 clknet_leaf_0_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
X_2250_ sap_3_inst.controller_inst.opcode\[5\] net760 _1667_ VPWR VGND sg13g2_nor2b_2
X_2181_ net751 _1596_ _1598_ VPWR VGND sg13g2_nor2_1
XFILLER_38_559 VPWR VGND sg13g2_decap_8
XFILLER_19_784 VPWR VGND sg13g2_decap_8
XFILLER_34_710 VPWR VGND sg13g2_decap_8
XFILLER_34_787 VPWR VGND sg13g2_decap_8
XFILLER_22_949 VPWR VGND sg13g2_decap_8
X_3704_ _1063_ _1149_ _1150_ VPWR VGND sg13g2_and2_1
X_3635_ _1091_ net610 _1047_ VPWR VGND sg13g2_nand2b_1
X_3566_ net15 net605 _1031_ VPWR VGND sg13g2_nor2_1
X_3497_ _0964_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[4\] net638
+ VPWR VGND sg13g2_nand2_1
X_2517_ _1932_ _1930_ _1931_ _1884_ net7 VPWR VGND sg13g2_a22oi_1
X_2448_ _1865_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[7\] net614
+ VPWR VGND sg13g2_nand2_1
X_2379_ _1653_ _1706_ _1796_ VPWR VGND sg13g2_nor2_1
XFILLER_29_537 VPWR VGND sg13g2_decap_8
X_4118_ u_ser.shadow_reg\[7\] u_ser.bit_pos\[1\] _1469_ VPWR VGND net800 sg13g2_nand3b_1
X_4049_ _1414_ _1415_ _1413_ _1419_ VPWR VGND _1418_ sg13g2_nand4_1
XFILLER_24_220 VPWR VGND sg13g2_fill_1
XFILLER_40_702 VPWR VGND sg13g2_decap_8
XFILLER_24_231 VPWR VGND sg13g2_fill_2
XFILLER_25_765 VPWR VGND sg13g2_decap_8
XFILLER_13_949 VPWR VGND sg13g2_decap_8
XFILLER_40_779 VPWR VGND sg13g2_decap_8
XFILLER_24_297 VPWR VGND sg13g2_fill_1
XFILLER_21_993 VPWR VGND sg13g2_decap_8
XFILLER_32_1015 VPWR VGND sg13g2_decap_8
XFILLER_4_669 VPWR VGND sg13g2_decap_8
XFILLER_0_875 VPWR VGND sg13g2_decap_8
XFILLER_47_312 VPWR VGND sg13g2_decap_8
Xhold8 _0157_ VPWR VGND net55 sg13g2_dlygate4sd3_1
XFILLER_48_857 VPWR VGND sg13g2_decap_8
XFILLER_47_389 VPWR VGND sg13g2_decap_8
XFILLER_16_765 VPWR VGND sg13g2_decap_8
XFILLER_43_584 VPWR VGND sg13g2_decap_8
XFILLER_31_768 VPWR VGND sg13g2_decap_8
XFILLER_8_920 VPWR VGND sg13g2_decap_8
XFILLER_12_982 VPWR VGND sg13g2_decap_8
XFILLER_11_481 VPWR VGND sg13g2_decap_8
XFILLER_8_997 VPWR VGND sg13g2_decap_8
XFILLER_7_485 VPWR VGND sg13g2_decap_8
XFILLER_48_1011 VPWR VGND sg13g2_decap_8
X_3420_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[1\] _0889_
+ net670 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[1\] _0890_ net641
+ sg13g2_a221oi_1
X_3351_ _1524_ _0667_ net690 _0822_ VPWR VGND sg13g2_nor3_1
X_2302_ VGND VPWR net740 _1718_ _1719_ _1589_ sg13g2_a21oi_1
X_3282_ _0652_ _0665_ _0708_ _0753_ VPWR VGND sg13g2_nor3_1
XFILLER_39_802 VPWR VGND sg13g2_decap_8
X_2233_ _1650_ _1603_ VPWR VGND _1576_ sg13g2_nand2b_2
XFILLER_39_879 VPWR VGND sg13g2_decap_8
X_2164_ _1581_ net747 sap_3_inst.controller_inst.stage\[1\] VPWR VGND sg13g2_nand2_2
XFILLER_0_60 VPWR VGND sg13g2_decap_8
XFILLER_19_581 VPWR VGND sg13g2_decap_8
X_2095_ VPWR _1513_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[1\]
+ VGND sg13g2_inv_1
XFILLER_34_584 VPWR VGND sg13g2_decap_8
XFILLER_10_919 VPWR VGND sg13g2_decap_8
XFILLER_22_746 VPWR VGND sg13g2_decap_8
X_2997_ _0490_ _0496_ net575 _0497_ VPWR VGND sg13g2_mux2_1
X_3618_ _0078_ _1075_ _1076_ net584 _1535_ VPWR VGND sg13g2_a22oi_1
X_3549_ _1014_ net640 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[6\]
+ net641 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_0_127 VPWR VGND sg13g2_decap_8
XFILLER_1_639 VPWR VGND sg13g2_decap_8
XFILLER_45_827 VPWR VGND sg13g2_decap_8
XFILLER_29_367 VPWR VGND sg13g2_fill_1
XFILLER_12_212 VPWR VGND sg13g2_fill_1
XFILLER_25_562 VPWR VGND sg13g2_decap_8
XFILLER_13_746 VPWR VGND sg13g2_decap_8
XFILLER_40_576 VPWR VGND sg13g2_decap_8
XFILLER_9_739 VPWR VGND sg13g2_decap_8
XFILLER_12_256 VPWR VGND sg13g2_fill_1
XFILLER_8_249 VPWR VGND sg13g2_fill_1
XFILLER_21_790 VPWR VGND sg13g2_decap_8
XFILLER_5_912 VPWR VGND sg13g2_decap_8
XFILLER_5_989 VPWR VGND sg13g2_decap_8
XFILLER_4_466 VPWR VGND sg13g2_decap_8
XFILLER_0_672 VPWR VGND sg13g2_decap_8
XFILLER_48_654 VPWR VGND sg13g2_decap_8
XFILLER_36_827 VPWR VGND sg13g2_decap_8
X_2920_ _0422_ net786 net708 VPWR VGND sg13g2_nand2_1
XFILLER_16_562 VPWR VGND sg13g2_decap_8
X_2851_ _0355_ _2012_ _0333_ VPWR VGND sg13g2_nand2_2
XFILLER_31_565 VPWR VGND sg13g2_decap_8
X_2782_ VPWR VGND _0215_ _1720_ _0211_ _1501_ net11 net633 sg13g2_a221oi_1
XFILLER_7_260 VPWR VGND sg13g2_fill_1
XFILLER_8_794 VPWR VGND sg13g2_decap_8
X_3403_ VPWR VGND _0873_ _0644_ _0288_ _1551_ _0874_ net737 sg13g2_a221oi_1
Xfanout729 _1583_ net729 VPWR VGND sg13g2_buf_8
Xfanout718 _1585_ net718 VPWR VGND sg13g2_buf_8
Xfanout707 _1830_ net707 VPWR VGND sg13g2_buf_2
X_3334_ _0690_ _0748_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[3\]
+ _0805_ VPWR VGND sg13g2_nand3_1
X_3265_ _1873_ _0733_ _0734_ _0735_ _0736_ VPWR VGND sg13g2_nor4_1
X_2216_ _1587_ net736 _1633_ VPWR VGND sg13g2_and2_1
X_3196_ _0667_ _0653_ _0664_ VPWR VGND sg13g2_nand2_2
XFILLER_27_805 VPWR VGND sg13g2_decap_8
XFILLER_39_676 VPWR VGND sg13g2_decap_8
X_2147_ net753 _1496_ _1564_ VPWR VGND sg13g2_nor2_1
X_2078_ VPWR _1496_ net756 VGND sg13g2_inv_1
XFILLER_22_543 VPWR VGND sg13g2_decap_8
XFILLER_10_716 VPWR VGND sg13g2_decap_8
XFILLER_2_904 VPWR VGND sg13g2_decap_8
XFILLER_18_816 VPWR VGND sg13g2_decap_8
XFILLER_45_624 VPWR VGND sg13g2_decap_8
XFILLER_44_112 VPWR VGND sg13g2_fill_2
XFILLER_17_326 VPWR VGND sg13g2_fill_1
XFILLER_32_307 VPWR VGND sg13g2_fill_1
XFILLER_38_1021 VPWR VGND sg13g2_decap_8
XFILLER_41_852 VPWR VGND sg13g2_decap_8
XFILLER_13_543 VPWR VGND sg13g2_decap_8
XFILLER_9_536 VPWR VGND sg13g2_decap_8
XFILLER_5_786 VPWR VGND sg13g2_decap_8
XFILLER_49_930 VPWR VGND sg13g2_decap_8
X_3050_ _0548_ net691 net772 _0357_ net780 VPWR VGND sg13g2_a22oi_1
XFILLER_48_451 VPWR VGND sg13g2_decap_8
XFILLER_36_624 VPWR VGND sg13g2_decap_8
XFILLER_24_808 VPWR VGND sg13g2_decap_8
X_3952_ _1329_ net803 _1550_ VPWR VGND sg13g2_nand2_1
X_2903_ _0405_ net786 sap_3_inst.alu_inst.tmp\[2\] VPWR VGND sg13g2_xnor2_1
X_3883_ net654 _1155_ _1280_ VPWR VGND sg13g2_nor2_1
X_2834_ _2055_ _0337_ _2004_ _0338_ VPWR VGND sg13g2_nand3_1
XFILLER_32_896 VPWR VGND sg13g2_decap_8
XFILLER_8_591 VPWR VGND sg13g2_decap_8
X_2765_ _1760_ _0289_ _0290_ _0291_ _0292_ VPWR VGND sg13g2_nor4_1
X_2696_ net19 _0227_ VPWR VGND sg13g2_inv_4
X_3317_ _0788_ net678 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[5\]
+ net684 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4297_ net833 VGND VPWR _0154_ sap_3_inst.reg_file_inst.array_serializer_inst.state\[0\]
+ clknet_3_5__leaf_clk sg13g2_dfrbpq_2
X_3248_ _0714_ _0715_ _0717_ _0718_ _0719_ VPWR VGND sg13g2_and4_1
XFILLER_27_602 VPWR VGND sg13g2_decap_8
X_3179_ _1869_ _0649_ _1555_ _0650_ VPWR VGND sg13g2_nand3_1
XFILLER_39_473 VPWR VGND sg13g2_decap_8
XFILLER_15_819 VPWR VGND sg13g2_decap_8
XFILLER_27_679 VPWR VGND sg13g2_decap_8
XFILLER_26_156 VPWR VGND sg13g2_fill_1
XFILLER_23_830 VPWR VGND sg13g2_decap_8
XFILLER_10_513 VPWR VGND sg13g2_decap_8
XFILLER_2_701 VPWR VGND sg13g2_decap_8
XFILLER_2_778 VPWR VGND sg13g2_decap_8
XFILLER_46_944 VPWR VGND sg13g2_decap_8
XFILLER_45_421 VPWR VGND sg13g2_decap_8
XFILLER_18_613 VPWR VGND sg13g2_decap_8
XFILLER_45_498 VPWR VGND sg13g2_decap_8
XFILLER_33_638 VPWR VGND sg13g2_decap_8
XFILLER_14_863 VPWR VGND sg13g2_decap_8
XFILLER_12_1024 VPWR VGND sg13g2_decap_4
X_2550_ _1959_ _1962_ _1963_ VPWR VGND sg13g2_and2_1
XFILLER_5_583 VPWR VGND sg13g2_decap_8
X_2481_ VGND VPWR _1759_ _1892_ _1898_ _1897_ sg13g2_a21oi_1
XFILLER_49_4 VPWR VGND sg13g2_fill_2
X_4220_ net830 VGND VPWR _0077_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[3\]
+ clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3102_ net789 sap_3_inst.out\[1\] net705 _0042_ VPWR VGND sg13g2_mux2_1
X_4082_ _1441_ VPWR _1442_ VGND _0331_ _1439_ sg13g2_o21ai_1
X_3033_ VGND VPWR sap_3_inst.alu_inst.act\[5\] _0320_ _0532_ net693 sg13g2_a21oi_1
XFILLER_37_922 VPWR VGND sg13g2_decap_8
XFILLER_24_605 VPWR VGND sg13g2_decap_8
XFILLER_37_999 VPWR VGND sg13g2_decap_8
XFILLER_36_498 VPWR VGND sg13g2_decap_8
X_3935_ _1317_ sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[2\] _1316_
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_833 VPWR VGND sg13g2_decap_8
XFILLER_32_693 VPWR VGND sg13g2_decap_8
X_3866_ _1004_ _1017_ _1267_ VPWR VGND sg13g2_nor2b_1
X_2817_ _1598_ _1760_ _1763_ _0321_ VPWR VGND sg13g2_nor3_1
X_3797_ net658 _1057_ _1220_ VPWR VGND sg13g2_nor2_1
X_2748_ VGND VPWR net726 _1682_ _0275_ _1650_ sg13g2_a21oi_1
XFILLER_11_59 VPWR VGND sg13g2_fill_1
X_2679_ _0209_ _0210_ _0211_ VPWR VGND sg13g2_and2_1
XFILLER_28_911 VPWR VGND sg13g2_decap_8
XFILLER_15_616 VPWR VGND sg13g2_decap_8
XFILLER_27_476 VPWR VGND sg13g2_decap_8
XFILLER_28_988 VPWR VGND sg13g2_decap_8
XFILLER_43_969 VPWR VGND sg13g2_decap_8
XFILLER_42_457 VPWR VGND sg13g2_decap_8
XFILLER_35_1002 VPWR VGND sg13g2_decap_8
XFILLER_10_321 VPWR VGND sg13g2_fill_2
XFILLER_10_343 VPWR VGND sg13g2_fill_2
XFILLER_11_866 VPWR VGND sg13g2_decap_8
XFILLER_2_575 VPWR VGND sg13g2_decap_8
XFILLER_42_1017 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_741 VPWR VGND sg13g2_decap_8
XFILLER_19_966 VPWR VGND sg13g2_decap_8
XFILLER_18_487 VPWR VGND sg13g2_decap_8
XFILLER_34_969 VPWR VGND sg13g2_decap_8
XFILLER_21_608 VPWR VGND sg13g2_decap_8
X_3720_ _1161_ VPWR _0095_ VGND _1081_ net582 sg13g2_o21ai_1
XFILLER_14_660 VPWR VGND sg13g2_decap_8
X_3651_ VGND VPWR net18 _1097_ _1105_ _0732_ sg13g2_a21oi_1
X_2602_ net704 _2010_ _2011_ VPWR VGND sg13g2_nor2_1
X_3582_ _0779_ VPWR _1046_ VGND net589 _0864_ sg13g2_o21ai_1
X_2533_ _1946_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[5\] net712
+ VPWR VGND sg13g2_nand2_1
X_2464_ _1879_ _1880_ _1759_ _1881_ VPWR VGND sg13g2_nand3_1
X_2395_ _1667_ _1753_ _1635_ _1812_ VPWR VGND sg13g2_nand3_1
X_4203_ net808 VGND VPWR _0060_ sap_3_inst.controller_inst.opcode\[2\] clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4134_ _1480_ _1481_ _0190_ VPWR VGND sg13g2_and2_1
XFILLER_29_719 VPWR VGND sg13g2_decap_8
XFILLER_3_1022 VPWR VGND sg13g2_decap_8
X_4065_ _0170_ _1063_ _1431_ net645 _1511_ VPWR VGND sg13g2_a22oi_1
X_3016_ _0513_ _0508_ _0515_ VPWR VGND sg13g2_xor2_1
XFILLER_24_402 VPWR VGND sg13g2_decap_8
XFILLER_19_1008 VPWR VGND sg13g2_decap_8
XFILLER_25_947 VPWR VGND sg13g2_decap_8
XFILLER_36_273 VPWR VGND sg13g2_fill_2
XFILLER_37_796 VPWR VGND sg13g2_decap_8
XFILLER_24_479 VPWR VGND sg13g2_decap_8
XFILLER_20_630 VPWR VGND sg13g2_decap_8
X_3918_ _1001_ VPWR _1304_ VGND _0304_ _1285_ sg13g2_o21ai_1
X_3849_ VGND VPWR _0927_ _1252_ _1254_ _1253_ sg13g2_a21oi_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_28_785 VPWR VGND sg13g2_decap_8
XFILLER_16_947 VPWR VGND sg13g2_decap_8
XFILLER_43_766 VPWR VGND sg13g2_decap_8
XFILLER_42_287 VPWR VGND sg13g2_fill_2
XFILLER_11_663 VPWR VGND sg13g2_decap_8
XFILLER_7_667 VPWR VGND sg13g2_decap_8
XFILLER_3_840 VPWR VGND sg13g2_decap_8
X_2180_ _1561_ net731 net765 _1597_ VPWR VGND _1595_ sg13g2_nand4_1
XFILLER_38_538 VPWR VGND sg13g2_decap_8
XFILLER_19_763 VPWR VGND sg13g2_decap_8
XFILLER_34_766 VPWR VGND sg13g2_decap_8
XFILLER_15_980 VPWR VGND sg13g2_decap_8
XFILLER_21_416 VPWR VGND sg13g2_fill_1
XFILLER_22_928 VPWR VGND sg13g2_decap_8
X_3703_ _0731_ VPWR _1149_ VGND _0719_ _0847_ sg13g2_o21ai_1
XFILLER_30_994 VPWR VGND sg13g2_decap_8
X_3634_ net24 _1087_ _1089_ _1090_ VPWR VGND sg13g2_nor3_2
X_3565_ VGND VPWR net663 _1027_ _1030_ _1029_ sg13g2_a21oi_1
X_3496_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[4\] _0962_
+ net647 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[4\] _0963_ net674
+ sg13g2_a221oi_1
X_2516_ _1902_ sap_3_inst.alu_flags\[6\] _1900_ _1931_ VPWR VGND sg13g2_a21o_1
X_2447_ VPWR VGND _1842_ _1808_ _1832_ net666 _1864_ net707 sg13g2_a221oi_1
X_2378_ VGND VPWR _1630_ _1670_ _1795_ _1794_ sg13g2_a21oi_1
XFILLER_29_516 VPWR VGND sg13g2_decap_8
X_4117_ _1468_ VPWR _0186_ VGND _1488_ u_ser.state\[1\] sg13g2_o21ai_1
XFILLER_44_519 VPWR VGND sg13g2_decap_8
X_4048_ _1418_ _1349_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[6\]
+ net796 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_25_744 VPWR VGND sg13g2_decap_8
XFILLER_37_593 VPWR VGND sg13g2_decap_8
XFILLER_13_928 VPWR VGND sg13g2_decap_8
XFILLER_24_265 VPWR VGND sg13g2_fill_2
XFILLER_40_758 VPWR VGND sg13g2_decap_8
XFILLER_12_438 VPWR VGND sg13g2_fill_2
XFILLER_21_972 VPWR VGND sg13g2_decap_8
XFILLER_4_648 VPWR VGND sg13g2_decap_8
XFILLER_0_854 VPWR VGND sg13g2_decap_8
XFILLER_48_836 VPWR VGND sg13g2_decap_8
Xhold9 u_ser.shadow_reg\[2\] VPWR VGND net56 sg13g2_dlygate4sd3_1
XFILLER_47_368 VPWR VGND sg13g2_decap_8
XFILLER_35_519 VPWR VGND sg13g2_decap_8
XFILLER_28_582 VPWR VGND sg13g2_decap_8
XFILLER_16_744 VPWR VGND sg13g2_decap_8
XFILLER_43_563 VPWR VGND sg13g2_decap_8
XFILLER_31_747 VPWR VGND sg13g2_decap_8
XFILLER_12_961 VPWR VGND sg13g2_decap_8
XFILLER_30_279 VPWR VGND sg13g2_fill_2
XFILLER_23_90 VPWR VGND sg13g2_decap_4
XFILLER_8_976 VPWR VGND sg13g2_decap_8
X_3350_ _1523_ net690 _0746_ _0821_ VPWR VGND sg13g2_nor3_1
X_2301_ _1590_ VPWR _1718_ VGND _1599_ _1717_ sg13g2_o21ai_1
XFILLER_2_180 VPWR VGND sg13g2_fill_2
X_3281_ _0752_ net681 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[0\]
+ net684 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2232_ _1576_ _1604_ _1649_ VPWR VGND sg13g2_nor2_2
X_2163_ net747 net746 _1580_ VPWR VGND sg13g2_and2_1
XFILLER_39_858 VPWR VGND sg13g2_decap_8
XFILLER_19_560 VPWR VGND sg13g2_decap_8
X_2094_ VPWR _1512_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[1\]
+ VGND sg13g2_inv_1
XFILLER_22_725 VPWR VGND sg13g2_decap_8
XFILLER_34_563 VPWR VGND sg13g2_decap_8
XFILLER_21_224 VPWR VGND sg13g2_fill_1
X_2996_ _0495_ VPWR _0496_ VGND _0471_ _0472_ sg13g2_o21ai_1
XFILLER_30_791 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_clk_div_out clknet_0_clk_div_out clknet_1_1__leaf_clk_div_out VPWR
+ VGND sg13g2_buf_8
X_3617_ net583 _1074_ _1076_ VPWR VGND sg13g2_nor2_1
X_3548_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[6\] _1012_
+ net647 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[6\] _1013_ net671
+ sg13g2_a221oi_1
XFILLER_0_117 VPWR VGND sg13g2_fill_1
XFILLER_1_618 VPWR VGND sg13g2_decap_8
X_3479_ net611 VPWR _0947_ VGND net665 _0946_ sg13g2_o21ai_1
XFILLER_45_806 VPWR VGND sg13g2_decap_8
XFILLER_25_541 VPWR VGND sg13g2_decap_8
XFILLER_13_725 VPWR VGND sg13g2_decap_8
XFILLER_9_718 VPWR VGND sg13g2_decap_8
XFILLER_40_555 VPWR VGND sg13g2_decap_8
XFILLER_5_968 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_fill_2
XFILLER_4_445 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_48_633 VPWR VGND sg13g2_decap_8
XFILLER_36_806 VPWR VGND sg13g2_decap_8
XFILLER_29_880 VPWR VGND sg13g2_decap_8
XFILLER_16_541 VPWR VGND sg13g2_decap_8
XFILLER_44_883 VPWR VGND sg13g2_decap_8
X_2850_ _0337_ _0351_ _2055_ _0354_ VPWR VGND _0352_ sg13g2_nand4_1
XFILLER_31_544 VPWR VGND sg13g2_decap_8
XFILLER_15_1022 VPWR VGND sg13g2_decap_8
X_2781_ VPWR net10 _0302_ VGND sg13g2_inv_1
XFILLER_8_773 VPWR VGND sg13g2_decap_8
XFILLER_11_290 VPWR VGND sg13g2_fill_2
X_3402_ _1620_ VPWR _0873_ VGND _0669_ _0872_ sg13g2_o21ai_1
X_3333_ _0804_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[3\] net672
+ VPWR VGND sg13g2_nand2_1
Xfanout708 net709 net708 VPWR VGND sg13g2_buf_8
Xfanout719 _1760_ net719 VPWR VGND sg13g2_buf_8
X_3264_ _0735_ _0635_ _0695_ VPWR VGND sg13g2_nand2_1
X_2215_ _1628_ net724 _1632_ VPWR VGND sg13g2_nor2_1
X_3195_ _0652_ _0665_ _0666_ VPWR VGND sg13g2_nor2_2
XFILLER_22_1026 VPWR VGND sg13g2_fill_2
XFILLER_39_655 VPWR VGND sg13g2_decap_8
X_2146_ net765 net768 _1563_ VPWR VGND net771 sg13g2_nand3b_1
X_2077_ VPWR _1495_ net758 VGND sg13g2_inv_1
XFILLER_35_883 VPWR VGND sg13g2_decap_8
XFILLER_22_522 VPWR VGND sg13g2_decap_8
XFILLER_14_48 VPWR VGND sg13g2_fill_1
X_2979_ _0477_ _0478_ _0479_ VPWR VGND sg13g2_and2_1
XFILLER_22_599 VPWR VGND sg13g2_decap_8
XFILLER_49_419 VPWR VGND sg13g2_decap_8
XFILLER_45_603 VPWR VGND sg13g2_decap_8
XFILLER_38_1000 VPWR VGND sg13g2_decap_8
XFILLER_41_831 VPWR VGND sg13g2_decap_8
XFILLER_13_522 VPWR VGND sg13g2_decap_8
XFILLER_26_894 VPWR VGND sg13g2_decap_8
XFILLER_9_515 VPWR VGND sg13g2_decap_8
XFILLER_13_599 VPWR VGND sg13g2_decap_8
XFILLER_5_765 VPWR VGND sg13g2_decap_8
XFILLER_1_982 VPWR VGND sg13g2_decap_8
XFILLER_49_986 VPWR VGND sg13g2_decap_8
XFILLER_48_430 VPWR VGND sg13g2_decap_8
XFILLER_36_603 VPWR VGND sg13g2_decap_8
X_3951_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[3\] sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[2\]
+ _1327_ sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[4\] _1328_ _1316_
+ sg13g2_a221oi_1
XFILLER_44_680 VPWR VGND sg13g2_decap_8
X_2902_ sap_3_inst.alu_inst.tmp\[2\] _0363_ net786 _0404_ VPWR VGND sg13g2_nand3_1
X_3882_ _1278_ VPWR _0139_ VGND _1150_ _1279_ sg13g2_o21ai_1
XFILLER_32_875 VPWR VGND sg13g2_decap_8
X_2833_ net704 _0336_ _0337_ VPWR VGND sg13g2_nor2b_2
X_2764_ net728 _1600_ _1762_ _0291_ VPWR VGND sg13g2_nor3_1
XFILLER_8_570 VPWR VGND sg13g2_decap_8
X_2695_ _0216_ _0218_ _0219_ _0226_ net19 VPWR VGND sg13g2_or4_1
X_3316_ _0787_ net681 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[5\]
+ net686 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[5\] VPWR VGND sg13g2_a22oi_1
X_4296_ net809 VGND VPWR _0153_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[7\]
+ clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3247_ VGND VPWR _0718_ _1744_ _1650_ sg13g2_or2_1
X_3178_ _0649_ net741 _1823_ VPWR VGND sg13g2_nand2_1
XFILLER_27_658 VPWR VGND sg13g2_decap_8
X_2129_ VPWR _1547_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[7\]
+ VGND sg13g2_inv_1
XFILLER_42_639 VPWR VGND sg13g2_decap_8
XFILLER_35_680 VPWR VGND sg13g2_decap_8
XFILLER_41_149 VPWR VGND sg13g2_fill_2
XFILLER_23_886 VPWR VGND sg13g2_decap_8
XFILLER_10_569 VPWR VGND sg13g2_decap_8
XFILLER_2_757 VPWR VGND sg13g2_decap_8
XFILLER_1_245 VPWR VGND sg13g2_fill_1
XFILLER_46_923 VPWR VGND sg13g2_decap_8
XFILLER_45_400 VPWR VGND sg13g2_decap_8
XFILLER_18_669 VPWR VGND sg13g2_decap_8
XFILLER_45_477 VPWR VGND sg13g2_decap_8
XFILLER_33_617 VPWR VGND sg13g2_decap_8
XFILLER_14_842 VPWR VGND sg13g2_decap_8
XFILLER_26_691 VPWR VGND sg13g2_decap_8
XFILLER_12_1003 VPWR VGND sg13g2_decap_8
XFILLER_5_562 VPWR VGND sg13g2_decap_8
X_2480_ VGND VPWR _1564_ _1894_ _1897_ _1896_ sg13g2_a21oi_1
X_3101_ _0596_ VPWR _0041_ VGND _1508_ net705 sg13g2_o21ai_1
X_4081_ _1440_ net694 _2002_ _1441_ VPWR VGND sg13g2_mux2_1
XFILLER_37_901 VPWR VGND sg13g2_decap_8
XFILLER_49_783 VPWR VGND sg13g2_decap_8
X_3032_ _0530_ VPWR _0531_ VGND _0505_ _0529_ sg13g2_o21ai_1
XFILLER_37_978 VPWR VGND sg13g2_decap_8
X_3934_ sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[1\] sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[0\]
+ _1316_ VPWR VGND sg13g2_and2_1
XFILLER_20_812 VPWR VGND sg13g2_decap_8
XFILLER_32_672 VPWR VGND sg13g2_decap_8
X_3865_ _0135_ _1125_ _1266_ net653 _1537_ VPWR VGND sg13g2_a22oi_1
X_2816_ _1895_ VPWR _0320_ VGND _1890_ _0319_ sg13g2_o21ai_1
XFILLER_20_889 VPWR VGND sg13g2_decap_8
X_3796_ _0113_ _1218_ _1219_ net581 _1547_ VPWR VGND sg13g2_a22oi_1
X_2747_ _1667_ _1893_ _1626_ _0274_ VPWR VGND sg13g2_nand3_1
XFILLER_11_27 VPWR VGND sg13g2_fill_2
X_2678_ _0210_ net620 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[2\]
+ net623 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[2\] VPWR VGND sg13g2_a22oi_1
X_4279_ net811 VGND VPWR _0136_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[6\]
+ clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_28_967 VPWR VGND sg13g2_decap_8
XFILLER_27_455 VPWR VGND sg13g2_decap_8
XFILLER_43_948 VPWR VGND sg13g2_decap_8
XFILLER_30_609 VPWR VGND sg13g2_decap_8
XFILLER_23_683 VPWR VGND sg13g2_decap_8
XFILLER_11_845 VPWR VGND sg13g2_decap_8
XFILLER_7_849 VPWR VGND sg13g2_decap_8
XFILLER_2_554 VPWR VGND sg13g2_decap_8
XFILLER_37_219 VPWR VGND sg13g2_fill_2
XFILLER_46_720 VPWR VGND sg13g2_decap_8
XFILLER_19_945 VPWR VGND sg13g2_decap_8
XFILLER_18_455 VPWR VGND sg13g2_decap_4
XFILLER_46_797 VPWR VGND sg13g2_decap_8
XFILLER_34_948 VPWR VGND sg13g2_decap_8
Xclkbuf_5_2__f_sap_3_inst.alu_inst.clk_regs clknet_4_1_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_9_175 VPWR VGND sg13g2_fill_2
X_3650_ VGND VPWR _1104_ net668 _0302_ sg13g2_or2_1
X_2601_ _2010_ _2005_ _2007_ VPWR VGND sg13g2_nand2_2
X_3581_ _1040_ _1020_ _1045_ VPWR VGND sg13g2_xor2_1
X_2532_ _1945_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[5\] net621
+ VPWR VGND sg13g2_nand2_1
X_2463_ _1880_ _1602_ _1829_ VPWR VGND sg13g2_nand2_1
X_4202_ net804 VGND VPWR _0059_ sap_3_inst.controller_inst.opcode\[1\] clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_2394_ VGND VPWR net768 _1765_ _1811_ _1759_ sg13g2_a21oi_1
X_4133_ _1479_ sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[0\] sap_3_inst.reg_file_inst.array_serializer_inst.word_index\[1\]
+ _1481_ VPWR VGND sg13g2_a21o_1
XFILLER_3_50 VPWR VGND sg13g2_fill_1
XFILLER_3_1001 VPWR VGND sg13g2_decap_8
X_4064_ net645 _1060_ _1431_ VPWR VGND sg13g2_nor2_1
XFILLER_49_580 VPWR VGND sg13g2_decap_8
X_3015_ _0508_ _0513_ _0514_ VPWR VGND sg13g2_nor2_1
X_4147__5 VPWR net39 clknet_leaf_2_sap_3_inst.alu_inst.clk VGND sg13g2_inv_1
XFILLER_25_926 VPWR VGND sg13g2_decap_8
XFILLER_37_775 VPWR VGND sg13g2_decap_8
XFILLER_24_458 VPWR VGND sg13g2_decap_8
XFILLER_11_119 VPWR VGND sg13g2_fill_1
XFILLER_33_981 VPWR VGND sg13g2_decap_8
X_3917_ _0993_ _1302_ _1303_ VPWR VGND sg13g2_nor2_1
X_3848_ net11 _0857_ _1064_ _1253_ VPWR VGND sg13g2_or3_1
XFILLER_20_686 VPWR VGND sg13g2_decap_8
X_3779_ _1205_ _1210_ _0105_ VPWR VGND sg13g2_nor2b_1
XFILLER_16_926 VPWR VGND sg13g2_decap_8
XFILLER_28_764 VPWR VGND sg13g2_decap_8
XFILLER_43_745 VPWR VGND sg13g2_decap_8
XFILLER_15_469 VPWR VGND sg13g2_decap_8
XFILLER_31_929 VPWR VGND sg13g2_decap_8
XFILLER_11_642 VPWR VGND sg13g2_decap_8
XFILLER_23_480 VPWR VGND sg13g2_decap_8
XFILLER_7_646 VPWR VGND sg13g2_decap_8
XFILLER_6_167 VPWR VGND sg13g2_fill_2
XFILLER_3_896 VPWR VGND sg13g2_decap_8
XFILLER_2_384 VPWR VGND sg13g2_fill_2
XFILLER_38_517 VPWR VGND sg13g2_decap_8
XFILLER_19_742 VPWR VGND sg13g2_decap_8
XFILLER_46_594 VPWR VGND sg13g2_decap_8
XFILLER_22_907 VPWR VGND sg13g2_decap_8
XFILLER_34_745 VPWR VGND sg13g2_decap_8
XFILLER_21_439 VPWR VGND sg13g2_fill_1
XFILLER_30_973 VPWR VGND sg13g2_decap_8
X_3702_ _1148_ VPWR _0090_ VGND _1522_ _1147_ sg13g2_o21ai_1
X_3633_ net587 VPWR _1089_ VGND net585 _1088_ sg13g2_o21ai_1
X_3564_ net592 VPWR _1029_ VGND net663 _1028_ sg13g2_o21ai_1
X_3495_ _0960_ _0961_ net661 _0962_ VPWR VGND sg13g2_nand3_1
X_2515_ VGND VPWR _1930_ _1899_ net777 sg13g2_or2_1
X_2446_ net667 net626 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[7\]
+ _1863_ VPWR VGND sg13g2_nand3_1
XFILLER_25_1024 VPWR VGND sg13g2_decap_4
X_4116_ _1465_ VPWR _1468_ VGND _1490_ _1466_ sg13g2_o21ai_1
X_2377_ _1638_ _1649_ _1794_ VPWR VGND sg13g2_nor2_1
X_4047_ _1417_ _1412_ _1416_ VPWR VGND sg13g2_nand2_1
XFILLER_25_723 VPWR VGND sg13g2_decap_8
XFILLER_37_572 VPWR VGND sg13g2_decap_8
XFILLER_13_907 VPWR VGND sg13g2_decap_8
XFILLER_24_244 VPWR VGND sg13g2_fill_2
XFILLER_40_737 VPWR VGND sg13g2_decap_8
XFILLER_21_951 VPWR VGND sg13g2_decap_8
XFILLER_20_483 VPWR VGND sg13g2_decap_8
XFILLER_4_627 VPWR VGND sg13g2_decap_8
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_48_815 VPWR VGND sg13g2_decap_8
XFILLER_47_347 VPWR VGND sg13g2_decap_8
XFILLER_16_723 VPWR VGND sg13g2_decap_8
XFILLER_28_561 VPWR VGND sg13g2_decap_8
XFILLER_43_542 VPWR VGND sg13g2_decap_8
XFILLER_15_222 VPWR VGND sg13g2_fill_1
XFILLER_31_726 VPWR VGND sg13g2_decap_8
XFILLER_12_940 VPWR VGND sg13g2_decap_8
XFILLER_8_955 VPWR VGND sg13g2_decap_8
XFILLER_7_421 VPWR VGND sg13g2_fill_2
X_2300_ VGND VPWR _1620_ _1716_ _1717_ _1622_ sg13g2_a21oi_1
X_3280_ _0751_ _0707_ _0748_ VPWR VGND sg13g2_nand2_1
X_2231_ _1638_ _1639_ _1643_ _1645_ _1648_ VPWR VGND sg13g2_or4_1
XFILLER_3_693 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_fill_2
X_2162_ VPWR _1579_ _1578_ VGND sg13g2_inv_1
XFILLER_39_837 VPWR VGND sg13g2_decap_8
X_2093_ VPWR _1511_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[1\]
+ VGND sg13g2_inv_1
XFILLER_26_509 VPWR VGND sg13g2_decap_8
XFILLER_0_1015 VPWR VGND sg13g2_decap_8
XFILLER_46_391 VPWR VGND sg13g2_decap_8
XFILLER_34_542 VPWR VGND sg13g2_decap_8
XFILLER_22_704 VPWR VGND sg13g2_decap_8
X_2995_ _0484_ _0486_ _0488_ _0494_ _0495_ VPWR VGND sg13g2_nor4_1
XFILLER_30_770 VPWR VGND sg13g2_decap_8
X_3616_ _0866_ _0981_ net611 _1075_ VPWR VGND sg13g2_nand3_1
X_3547_ _1010_ _1011_ net661 _1012_ VPWR VGND sg13g2_nand3_1
X_3478_ _0946_ _0813_ _0930_ VPWR VGND sg13g2_xnor2_1
X_2429_ _1846_ _1545_ net631 VPWR VGND sg13g2_nand2_1
XFILLER_44_328 VPWR VGND sg13g2_fill_1
XFILLER_38_881 VPWR VGND sg13g2_decap_8
XFILLER_25_520 VPWR VGND sg13g2_decap_8
XFILLER_13_704 VPWR VGND sg13g2_decap_8
XFILLER_40_534 VPWR VGND sg13g2_decap_8
XFILLER_25_597 VPWR VGND sg13g2_decap_8
XFILLER_5_947 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_48_612 VPWR VGND sg13g2_decap_8
XFILLER_48_689 VPWR VGND sg13g2_decap_8
XFILLER_16_520 VPWR VGND sg13g2_decap_8
XFILLER_44_862 VPWR VGND sg13g2_decap_8
XFILLER_16_597 VPWR VGND sg13g2_decap_8
XFILLER_31_523 VPWR VGND sg13g2_decap_8
XFILLER_15_1001 VPWR VGND sg13g2_decap_8
X_2780_ _0302_ net576 _2035_ VPWR VGND sg13g2_nand2_2
XFILLER_8_752 VPWR VGND sg13g2_decap_8
X_3401_ _0872_ _0679_ _0682_ _0871_ VPWR VGND sg13g2_and3_1
X_3332_ _0800_ _0801_ _0799_ _0803_ VPWR VGND sg13g2_nand3_1
Xfanout709 _2014_ net709 VPWR VGND sg13g2_buf_8
XFILLER_4_991 VPWR VGND sg13g2_decap_8
XFILLER_3_490 VPWR VGND sg13g2_decap_8
X_3263_ VGND VPWR _1681_ net721 _0734_ _1653_ sg13g2_a21oi_1
X_2214_ _1631_ net737 net736 _1580_ net743 VPWR VGND sg13g2_a22oi_1
X_3194_ _0665_ _0662_ _0663_ VPWR VGND sg13g2_nand2_2
XFILLER_22_1005 VPWR VGND sg13g2_decap_8
XFILLER_39_634 VPWR VGND sg13g2_decap_8
X_2145_ _1562_ net768 VPWR VGND net770 sg13g2_nand2b_2
XFILLER_15_0 VPWR VGND sg13g2_fill_1
X_2076_ _1494_ net766 VPWR VGND sg13g2_inv_2
XFILLER_22_501 VPWR VGND sg13g2_decap_8
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_35_862 VPWR VGND sg13g2_decap_8
XFILLER_22_578 VPWR VGND sg13g2_decap_8
X_2978_ _0443_ _0474_ _0476_ _0478_ VPWR VGND sg13g2_or3_1
XFILLER_2_939 VPWR VGND sg13g2_decap_8
XFILLER_45_659 VPWR VGND sg13g2_decap_8
XFILLER_41_810 VPWR VGND sg13g2_decap_8
XFILLER_13_501 VPWR VGND sg13g2_decap_8
XFILLER_26_873 VPWR VGND sg13g2_decap_8
XFILLER_41_887 VPWR VGND sg13g2_decap_8
XFILLER_40_386 VPWR VGND sg13g2_fill_1
XFILLER_13_578 VPWR VGND sg13g2_decap_8
XFILLER_5_744 VPWR VGND sg13g2_decap_8
XFILLER_45_1016 VPWR VGND sg13g2_decap_8
XFILLER_45_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_961 VPWR VGND sg13g2_decap_8
XFILLER_49_965 VPWR VGND sg13g2_decap_8
XFILLER_48_486 VPWR VGND sg13g2_decap_8
XFILLER_36_659 VPWR VGND sg13g2_decap_8
XFILLER_17_884 VPWR VGND sg13g2_decap_8
X_3950_ net803 sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[1\] _1327_
+ VPWR VGND sg13g2_nor2b_1
X_2901_ VPWR _0034_ _0403_ VGND sg13g2_inv_1
X_3881_ _1279_ net671 _1151_ VPWR VGND sg13g2_nand2_1
XFILLER_32_854 VPWR VGND sg13g2_decap_8
X_2832_ _2009_ _0333_ _2004_ _0336_ VPWR VGND sg13g2_nand3_1
X_2763_ net716 net725 _0290_ VPWR VGND sg13g2_nor2_1
X_2694_ VGND VPWR _0222_ _0225_ _0226_ _1720_ sg13g2_a21oi_1
XFILLER_6_72 VPWR VGND sg13g2_decap_4
X_4295_ net812 VGND VPWR _0152_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[6\]
+ clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3315_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[6\] _0785_
+ net651 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[6\] _0786_ net671
+ sg13g2_a221oi_1
X_3246_ VGND VPWR net764 _0644_ _0717_ _0716_ sg13g2_a21oi_1
X_3177_ _0648_ net740 _0647_ VPWR VGND sg13g2_nand2_1
XFILLER_27_637 VPWR VGND sg13g2_decap_8
X_2128_ VPWR _1546_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[7\]
+ VGND sg13g2_inv_1
XFILLER_42_618 VPWR VGND sg13g2_decap_8
XFILLER_23_865 VPWR VGND sg13g2_decap_8
XFILLER_10_548 VPWR VGND sg13g2_decap_8
XFILLER_6_519 VPWR VGND sg13g2_decap_8
XFILLER_2_736 VPWR VGND sg13g2_decap_8
XFILLER_46_902 VPWR VGND sg13g2_decap_8
XFILLER_18_648 VPWR VGND sg13g2_decap_8
XFILLER_46_979 VPWR VGND sg13g2_decap_8
XFILLER_45_456 VPWR VGND sg13g2_decap_8
XFILLER_14_821 VPWR VGND sg13g2_decap_8
XFILLER_26_670 VPWR VGND sg13g2_decap_8
XFILLER_32_106 VPWR VGND sg13g2_fill_2
XFILLER_41_684 VPWR VGND sg13g2_decap_8
XFILLER_9_324 VPWR VGND sg13g2_fill_1
XFILLER_14_898 VPWR VGND sg13g2_decap_8
XFILLER_40_183 VPWR VGND sg13g2_fill_2
XFILLER_5_541 VPWR VGND sg13g2_decap_8
X_3100_ _0596_ sap_3_inst.out\[0\] net705 VPWR VGND sg13g2_nand2_1
X_4080_ _2013_ _2054_ _1440_ VPWR VGND sg13g2_nor2_1
XFILLER_49_762 VPWR VGND sg13g2_decap_8
X_3031_ VGND VPWR _0353_ _0519_ _0530_ net702 sg13g2_a21oi_1
XFILLER_36_412 VPWR VGND sg13g2_fill_1
XFILLER_37_957 VPWR VGND sg13g2_decap_8
XFILLER_36_456 VPWR VGND sg13g2_fill_2
XFILLER_17_681 VPWR VGND sg13g2_decap_8
X_3933_ net78 sap_3_inst.reg_file_inst.array_serializer_inst.state\[1\] _1315_ VPWR
+ VGND sg13g2_nor2b_2
XFILLER_32_651 VPWR VGND sg13g2_decap_8
X_3864_ VGND VPWR _1263_ _1264_ _1266_ _1265_ sg13g2_a21oi_1
X_2815_ _1759_ VPWR _0319_ VGND net716 _1886_ sg13g2_o21ai_1
XFILLER_20_868 VPWR VGND sg13g2_decap_8
X_3795_ net24 _1087_ net581 _1219_ VPWR VGND sg13g2_nor3_1
X_2746_ _1579_ _0273_ mem_ram_we VPWR VGND sg13g2_nor2_1
X_2677_ _0209_ net615 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[2\]
+ net625 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[2\] VPWR VGND sg13g2_a22oi_1
X_4278_ net810 VGND VPWR _0135_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[5\]
+ clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3229_ VGND VPWR _1627_ _1633_ _0700_ _1657_ sg13g2_a21oi_1
XFILLER_27_434 VPWR VGND sg13g2_decap_8
XFILLER_28_946 VPWR VGND sg13g2_decap_8
XFILLER_43_927 VPWR VGND sg13g2_decap_8
XFILLER_42_426 VPWR VGND sg13g2_decap_8
XFILLER_11_824 VPWR VGND sg13g2_decap_8
XFILLER_23_662 VPWR VGND sg13g2_decap_8
XFILLER_7_828 VPWR VGND sg13g2_decap_8
XFILLER_2_533 VPWR VGND sg13g2_decap_8
XFILLER_19_924 VPWR VGND sg13g2_decap_8
XFILLER_46_776 VPWR VGND sg13g2_decap_8
XFILLER_34_927 VPWR VGND sg13g2_decap_8
XFILLER_42_982 VPWR VGND sg13g2_decap_8
XFILLER_41_481 VPWR VGND sg13g2_decap_8
XFILLER_14_695 VPWR VGND sg13g2_decap_8
XFILLER_9_187 VPWR VGND sg13g2_fill_1
X_2600_ _1571_ net728 _1617_ _2009_ VPWR VGND sg13g2_nor3_1
X_3580_ VGND VPWR net660 _1043_ _1044_ net612 sg13g2_a21oi_1
X_2531_ net667 net626 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[5\]
+ _1944_ VPWR VGND sg13g2_nand3_1
XFILLER_6_883 VPWR VGND sg13g2_decap_8
X_2462_ _1878_ VPWR _1879_ VGND _1634_ _1871_ sg13g2_o21ai_1
X_4201_ net804 VGND VPWR _0058_ sap_3_inst.controller_inst.opcode\[0\] clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_2393_ VGND VPWR _1810_ _1807_ net696 sg13g2_or2_1
XFILLER_3_73 VPWR VGND sg13g2_decap_4
X_4132_ _1480_ _1479_ _1336_ VPWR VGND sg13g2_nand2b_1
X_4063_ net645 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[0\] _1430_
+ _0169_ VPWR VGND sg13g2_a21o_1
X_3014_ _0477_ _0512_ _0513_ VPWR VGND sg13g2_and2_1
XFILLER_25_905 VPWR VGND sg13g2_decap_8
XFILLER_37_754 VPWR VGND sg13g2_decap_8
XFILLER_40_919 VPWR VGND sg13g2_decap_8
XFILLER_24_437 VPWR VGND sg13g2_decap_8
XFILLER_33_960 VPWR VGND sg13g2_decap_8
X_3916_ net594 VPWR _1302_ VGND net647 _0995_ sg13g2_o21ai_1
XFILLER_20_665 VPWR VGND sg13g2_decap_8
X_3847_ VGND VPWR _0897_ _0914_ _1252_ _0881_ sg13g2_a21oi_1
X_3778_ _1145_ _1207_ net675 _1210_ VPWR VGND _1209_ sg13g2_nand4_1
XFILLER_4_809 VPWR VGND sg13g2_decap_8
X_2729_ _0259_ net600 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[0\]
+ net630 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[0\] VPWR VGND sg13g2_a22oi_1
Xclkbuf_5_26__f_sap_3_inst.alu_inst.clk_regs clknet_4_13_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_47_529 VPWR VGND sg13g2_decap_8
XFILLER_28_743 VPWR VGND sg13g2_decap_8
XFILLER_16_905 VPWR VGND sg13g2_decap_8
XFILLER_43_724 VPWR VGND sg13g2_decap_8
XFILLER_42_212 VPWR VGND sg13g2_fill_1
XFILLER_31_908 VPWR VGND sg13g2_decap_8
XFILLER_42_289 VPWR VGND sg13g2_fill_1
XFILLER_11_621 VPWR VGND sg13g2_decap_8
XFILLER_7_625 VPWR VGND sg13g2_decap_8
XFILLER_11_698 VPWR VGND sg13g2_decap_8
Xclkbuf_5_15__f_sap_3_inst.alu_inst.clk_regs clknet_4_7_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_3_875 VPWR VGND sg13g2_decap_8
XFILLER_19_721 VPWR VGND sg13g2_decap_8
XFILLER_46_573 VPWR VGND sg13g2_decap_8
XFILLER_19_798 VPWR VGND sg13g2_decap_8
XFILLER_34_724 VPWR VGND sg13g2_decap_8
XFILLER_14_492 VPWR VGND sg13g2_decap_8
XFILLER_33_289 VPWR VGND sg13g2_fill_2
XFILLER_30_952 VPWR VGND sg13g2_decap_8
X_3701_ _1057_ _1058_ net582 _1148_ VPWR VGND sg13g2_or3_1
X_3632_ _1088_ _0779_ _0864_ VPWR VGND sg13g2_xnor2_1
X_3563_ _0851_ _0786_ _1028_ VPWR VGND sg13g2_xor2_1
XFILLER_6_680 VPWR VGND sg13g2_decap_8
X_3494_ _0961_ net682 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[4\]
+ net685 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[4\] VPWR VGND sg13g2_a22oi_1
X_2514_ VGND VPWR _1929_ _1928_ _1768_ sg13g2_or2_1
X_2445_ net667 net627 _1862_ VPWR VGND sg13g2_and2_1
XFILLER_25_1003 VPWR VGND sg13g2_decap_8
X_4115_ _1467_ _1465_ _1466_ VPWR VGND sg13g2_nand2_1
X_2376_ VPWR _1793_ net696 VGND sg13g2_inv_1
X_4046_ _1416_ _1351_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[6\]
+ _1346_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_37_551 VPWR VGND sg13g2_decap_8
XFILLER_25_702 VPWR VGND sg13g2_decap_8
XFILLER_40_716 VPWR VGND sg13g2_decap_8
XFILLER_25_779 VPWR VGND sg13g2_decap_8
XFILLER_21_930 VPWR VGND sg13g2_decap_8
XFILLER_4_606 VPWR VGND sg13g2_decap_8
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_47_326 VPWR VGND sg13g2_decap_8
XFILLER_28_540 VPWR VGND sg13g2_decap_8
XFILLER_16_702 VPWR VGND sg13g2_decap_8
XFILLER_43_521 VPWR VGND sg13g2_decap_8
XFILLER_16_779 VPWR VGND sg13g2_decap_8
XFILLER_31_705 VPWR VGND sg13g2_decap_8
XFILLER_43_598 VPWR VGND sg13g2_decap_8
XFILLER_8_934 VPWR VGND sg13g2_decap_8
XFILLER_12_996 VPWR VGND sg13g2_decap_8
XFILLER_11_495 VPWR VGND sg13g2_decap_8
XFILLER_7_499 VPWR VGND sg13g2_decap_8
XFILLER_48_1025 VPWR VGND sg13g2_decap_4
XFILLER_3_672 VPWR VGND sg13g2_decap_8
X_2230_ _1643_ _1645_ _1647_ VPWR VGND sg13g2_nor2_1
XFILLER_2_182 VPWR VGND sg13g2_fill_1
XFILLER_39_816 VPWR VGND sg13g2_decap_8
X_2161_ _1578_ _1574_ _1577_ net742 _1559_ VPWR VGND sg13g2_a22oi_1
X_2092_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[1\] _1510_ VPWR
+ VGND sg13g2_inv_4
XFILLER_47_893 VPWR VGND sg13g2_decap_8
XFILLER_46_370 VPWR VGND sg13g2_decap_8
XFILLER_0_85 VPWR VGND sg13g2_fill_1
XFILLER_0_74 VPWR VGND sg13g2_decap_8
XFILLER_19_595 VPWR VGND sg13g2_decap_8
XFILLER_34_521 VPWR VGND sg13g2_decap_8
X_2994_ _0493_ VPWR _0494_ VGND _0355_ _0474_ sg13g2_o21ai_1
XFILLER_34_598 VPWR VGND sg13g2_decap_8
X_3615_ VGND VPWR _1074_ _1073_ net21 sg13g2_or2_1
X_3546_ _1011_ net675 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[6\]
+ net686 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_0_108 VPWR VGND sg13g2_fill_2
X_3477_ _0942_ VPWR _0945_ VGND _0825_ net572 sg13g2_o21ai_1
X_2428_ VPWR VGND _1842_ _1810_ _1832_ net666 _1845_ net707 sg13g2_a221oi_1
X_2359_ _1639_ _1690_ _1776_ VPWR VGND sg13g2_nor2_1
XFILLER_28_48 VPWR VGND sg13g2_fill_2
X_4029_ _0154_ VPWR _1401_ VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[4\]
+ _1344_ sg13g2_o21ai_1
XFILLER_38_860 VPWR VGND sg13g2_decap_8
XFILLER_25_576 VPWR VGND sg13g2_decap_8
XFILLER_40_513 VPWR VGND sg13g2_decap_8
XFILLER_20_270 VPWR VGND sg13g2_fill_1
XFILLER_5_926 VPWR VGND sg13g2_decap_8
XFILLER_4_403 VPWR VGND sg13g2_fill_2
XFILLER_0_686 VPWR VGND sg13g2_decap_8
XFILLER_48_668 VPWR VGND sg13g2_decap_8
XFILLER_35_329 VPWR VGND sg13g2_fill_1
XFILLER_44_841 VPWR VGND sg13g2_decap_8
XFILLER_16_576 VPWR VGND sg13g2_decap_8
XFILLER_31_502 VPWR VGND sg13g2_decap_8
XFILLER_34_80 VPWR VGND sg13g2_fill_1
XFILLER_8_731 VPWR VGND sg13g2_decap_8
XFILLER_31_579 VPWR VGND sg13g2_decap_8
XFILLER_11_292 VPWR VGND sg13g2_fill_1
XFILLER_12_793 VPWR VGND sg13g2_decap_8
X_3400_ VPWR VGND _1645_ _0723_ _0672_ net734 _0871_ _1705_ sg13g2_a221oi_1
X_3331_ _0802_ _0799_ _0800_ _0801_ VPWR VGND sg13g2_and3_2
XFILLER_4_970 VPWR VGND sg13g2_decap_8
X_3262_ _0733_ _0654_ _0691_ _1783_ _1634_ VPWR VGND sg13g2_a22oi_1
X_2213_ _1630_ net737 net736 VPWR VGND sg13g2_nand2_2
X_3193_ _0662_ _0663_ _0664_ VPWR VGND sg13g2_and2_1
XFILLER_39_613 VPWR VGND sg13g2_decap_8
X_2144_ net770 net767 _1561_ VPWR VGND sg13g2_nor2b_2
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_819 VPWR VGND sg13g2_decap_8
XFILLER_47_690 VPWR VGND sg13g2_decap_8
X_2075_ net764 _1493_ VPWR VGND sg13g2_inv_4
XFILLER_35_841 VPWR VGND sg13g2_decap_8
XFILLER_34_373 VPWR VGND sg13g2_fill_2
XFILLER_22_557 VPWR VGND sg13g2_decap_8
X_2977_ _0474_ VPWR _0477_ VGND _0443_ _0476_ sg13g2_o21ai_1
XFILLER_30_38 VPWR VGND sg13g2_fill_2
XFILLER_2_918 VPWR VGND sg13g2_decap_8
X_3529_ _0995_ _0851_ _0994_ VPWR VGND sg13g2_nand2_2
XFILLER_45_638 VPWR VGND sg13g2_decap_8
XFILLER_26_852 VPWR VGND sg13g2_decap_8
XFILLER_41_866 VPWR VGND sg13g2_decap_8
XFILLER_13_557 VPWR VGND sg13g2_decap_8
XFILLER_5_723 VPWR VGND sg13g2_decap_8
XFILLER_1_940 VPWR VGND sg13g2_decap_8
XFILLER_49_944 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_48_465 VPWR VGND sg13g2_decap_8
XFILLER_36_638 VPWR VGND sg13g2_decap_8
XFILLER_17_863 VPWR VGND sg13g2_decap_8
X_2900_ _0403_ _0401_ _0402_ net599 net790 VPWR VGND sg13g2_a22oi_1
XFILLER_32_833 VPWR VGND sg13g2_decap_8
XFILLER_43_181 VPWR VGND sg13g2_fill_1
X_3880_ _1278_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[1\] net652
+ VPWR VGND sg13g2_nand2_1
X_2831_ _2008_ _0333_ _2004_ _0335_ VPWR VGND sg13g2_nand3_1
X_2762_ VPWR VGND _1995_ _1602_ _0287_ _0278_ _0289_ _0286_ sg13g2_a221oi_1
XFILLER_12_590 VPWR VGND sg13g2_decap_8
XFILLER_6_40 VPWR VGND sg13g2_fill_1
X_2693_ _0220_ _0221_ _0223_ _0224_ _0225_ VPWR VGND sg13g2_and4_1
X_4294_ net814 VGND VPWR _0151_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[5\]
+ clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3314_ _0782_ _0783_ _0781_ _0785_ VPWR VGND _0784_ sg13g2_nand4_1
X_3245_ _1651_ _0631_ _0716_ VPWR VGND sg13g2_nor2_1
X_3176_ _0642_ _0641_ _0646_ _0647_ VPWR VGND sg13g2_a21o_2
XFILLER_27_616 VPWR VGND sg13g2_decap_8
XFILLER_39_487 VPWR VGND sg13g2_decap_8
X_2127_ _1545_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[7\] VPWR
+ VGND sg13g2_inv_2
XFILLER_22_343 VPWR VGND sg13g2_fill_2
XFILLER_23_844 VPWR VGND sg13g2_decap_8
XFILLER_10_527 VPWR VGND sg13g2_decap_8
XFILLER_2_715 VPWR VGND sg13g2_decap_8
XFILLER_49_218 VPWR VGND sg13g2_fill_2
XFILLER_18_627 VPWR VGND sg13g2_decap_8
XFILLER_46_958 VPWR VGND sg13g2_decap_8
XFILLER_45_435 VPWR VGND sg13g2_decap_8
XFILLER_14_800 VPWR VGND sg13g2_decap_8
XFILLER_41_663 VPWR VGND sg13g2_decap_8
XFILLER_14_877 VPWR VGND sg13g2_decap_8
XFILLER_5_520 VPWR VGND sg13g2_decap_8
XFILLER_5_597 VPWR VGND sg13g2_decap_8
XFILLER_49_741 VPWR VGND sg13g2_decap_8
X_3030_ _0511_ _0517_ _0354_ _0529_ VPWR VGND _0528_ sg13g2_nand4_1
XFILLER_37_936 VPWR VGND sg13g2_decap_8
XFILLER_24_619 VPWR VGND sg13g2_decap_8
XFILLER_17_660 VPWR VGND sg13g2_decap_8
XFILLER_32_630 VPWR VGND sg13g2_decap_8
X_3932_ _1314_ net78 VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.state\[1\]
+ sg13g2_nand2b_2
X_3863_ _1265_ _0304_ net674 VPWR VGND sg13g2_nand2_1
X_2814_ net57 sap_3_inst.out\[7\] net799 _0024_ VPWR VGND sg13g2_mux2_1
XFILLER_20_847 VPWR VGND sg13g2_decap_8
X_3794_ net607 VPWR _1218_ VGND net683 _1047_ sg13g2_o21ai_1
XFILLER_11_29 VPWR VGND sg13g2_fill_1
X_2745_ _0273_ _1896_ _0272_ net722 net739 VPWR VGND sg13g2_a22oi_1
X_2676_ _2058_ VPWR _0027_ VGND _2057_ _0208_ sg13g2_o21ai_1
XFILLER_28_1023 VPWR VGND sg13g2_decap_4
X_4346_ regFile_serial_start net30 VPWR VGND sg13g2_buf_8
X_4277_ net811 VGND VPWR _0134_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[4\]
+ clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3228_ _0695_ _0696_ _0694_ _0699_ VPWR VGND _0698_ sg13g2_nand4_1
XFILLER_28_925 VPWR VGND sg13g2_decap_8
X_3159_ _0630_ _1627_ net720 VPWR VGND sg13g2_nand2b_1
XFILLER_43_906 VPWR VGND sg13g2_decap_8
XFILLER_23_641 VPWR VGND sg13g2_decap_8
XFILLER_11_803 VPWR VGND sg13g2_decap_8
XFILLER_35_1016 VPWR VGND sg13g2_decap_8
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_7_807 VPWR VGND sg13g2_decap_8
XFILLER_2_512 VPWR VGND sg13g2_decap_8
XFILLER_2_589 VPWR VGND sg13g2_decap_8
XFILLER_19_903 VPWR VGND sg13g2_decap_8
XFILLER_46_755 VPWR VGND sg13g2_decap_8
XFILLER_34_906 VPWR VGND sg13g2_decap_8
XFILLER_27_980 VPWR VGND sg13g2_decap_8
XFILLER_42_961 VPWR VGND sg13g2_decap_8
XFILLER_41_460 VPWR VGND sg13g2_decap_8
XFILLER_14_674 VPWR VGND sg13g2_decap_8
XFILLER_9_177 VPWR VGND sg13g2_fill_1
X_2530_ _1943_ net632 sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[5\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_6_862 VPWR VGND sg13g2_decap_8
XFILLER_10_891 VPWR VGND sg13g2_decap_8
X_2461_ _1873_ _1874_ _1875_ _1877_ _1878_ VPWR VGND sg13g2_nor4_1
X_4200_ net817 VGND VPWR _0057_ sap_3_inst.alu_inst.tmp\[7\] clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_2
X_2392_ net696 _1807_ _1809_ VPWR VGND sg13g2_nor2_2
X_4131_ _1479_ net77 _0189_ VPWR VGND sg13g2_xor2_1
XFILLER_3_63 VPWR VGND sg13g2_decap_4
X_4062_ net645 _1057_ _1058_ _1430_ VPWR VGND sg13g2_nor3_1
X_3013_ _0512_ net781 sap_3_inst.alu_inst.tmp\[4\] VPWR VGND sg13g2_nand2b_1
XFILLER_37_733 VPWR VGND sg13g2_decap_8
XFILLER_18_991 VPWR VGND sg13g2_decap_8
XFILLER_24_416 VPWR VGND sg13g2_decap_8
X_3915_ net643 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[4\] _1301_
+ _0150_ VPWR VGND sg13g2_a21o_1
XFILLER_20_644 VPWR VGND sg13g2_decap_8
X_3846_ _0131_ _1251_ _0302_ net652 _1513_ VPWR VGND sg13g2_a22oi_1
X_3777_ _1209_ _1208_ _1041_ VPWR VGND sg13g2_nand2b_1
X_2728_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[0\] net620
+ _1850_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[0\] _0258_ net712
+ sg13g2_a221oi_1
X_2659_ _2066_ net622 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[3\]
+ _1847_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[3\] VPWR VGND sg13g2_a22oi_1
X_4329_ net817 VGND VPWR _0186_ u_ser.state\[1\] clknet_3_1__leaf_clk sg13g2_dfrbpq_2
XFILLER_47_508 VPWR VGND sg13g2_decap_8
XFILLER_41_1020 VPWR VGND sg13g2_decap_8
XFILLER_47_69 VPWR VGND sg13g2_fill_1
XFILLER_28_722 VPWR VGND sg13g2_decap_8
XFILLER_43_703 VPWR VGND sg13g2_decap_8
XFILLER_28_799 VPWR VGND sg13g2_decap_8
XFILLER_27_287 VPWR VGND sg13g2_fill_1
XFILLER_11_600 VPWR VGND sg13g2_decap_8
XFILLER_24_983 VPWR VGND sg13g2_decap_8
XFILLER_7_604 VPWR VGND sg13g2_decap_8
XFILLER_10_176 VPWR VGND sg13g2_fill_2
XFILLER_10_154 VPWR VGND sg13g2_fill_2
XFILLER_6_125 VPWR VGND sg13g2_fill_1
XFILLER_11_677 VPWR VGND sg13g2_decap_8
XFILLER_3_854 VPWR VGND sg13g2_decap_8
XFILLER_19_700 VPWR VGND sg13g2_decap_8
Xfanout690 _0709_ net690 VPWR VGND sg13g2_buf_1
XFILLER_46_552 VPWR VGND sg13g2_decap_8
XFILLER_19_777 VPWR VGND sg13g2_decap_8
XFILLER_34_703 VPWR VGND sg13g2_decap_8
XFILLER_37_80 VPWR VGND sg13g2_fill_1
XFILLER_15_994 VPWR VGND sg13g2_decap_8
XFILLER_30_931 VPWR VGND sg13g2_decap_8
X_3700_ VGND VPWR _1147_ net604 net669 sg13g2_or2_1
X_3631_ net612 _1043_ _1087_ VPWR VGND sg13g2_nor2_1
X_3562_ _1025_ _1026_ _1027_ VPWR VGND sg13g2_and2_1
X_2513_ _1918_ VPWR _1928_ VGND _1925_ _1927_ sg13g2_o21ai_1
X_3493_ _0960_ net678 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[4\]
+ net686 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[4\] VPWR VGND sg13g2_a22oi_1
X_2444_ _1861_ net616 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[7\]
+ net619 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[7\] VPWR VGND
+ sg13g2_a22oi_1
X_2375_ _1555_ _1578_ _1790_ _1791_ _1792_ VPWR VGND sg13g2_and4_1
XFILLER_38_0 VPWR VGND sg13g2_fill_2
X_4114_ _1466_ u_ser.bit_pos\[1\] net800 VPWR VGND sg13g2_nand2_1
X_4045_ _1415_ _1347_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[6\]
+ _1340_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_37_530 VPWR VGND sg13g2_decap_8
XFILLER_25_758 VPWR VGND sg13g2_decap_8
XFILLER_12_419 VPWR VGND sg13g2_fill_1
XFILLER_32_1008 VPWR VGND sg13g2_decap_8
X_3829_ _1238_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[6\] net634
+ VPWR VGND sg13g2_nand2_1
XFILLER_21_986 VPWR VGND sg13g2_decap_8
XFILLER_3_139 VPWR VGND sg13g2_fill_2
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_47_305 VPWR VGND sg13g2_fill_2
XFILLER_43_500 VPWR VGND sg13g2_decap_8
XFILLER_16_758 VPWR VGND sg13g2_decap_8
XFILLER_28_596 VPWR VGND sg13g2_decap_8
XFILLER_43_577 VPWR VGND sg13g2_decap_8
XFILLER_24_780 VPWR VGND sg13g2_decap_8
XFILLER_8_913 VPWR VGND sg13g2_decap_8
XFILLER_12_975 VPWR VGND sg13g2_decap_8
XFILLER_7_478 VPWR VGND sg13g2_decap_8
XFILLER_48_1004 VPWR VGND sg13g2_decap_8
XFILLER_3_651 VPWR VGND sg13g2_decap_8
X_2160_ _1575_ _1576_ _1577_ VPWR VGND sg13g2_nor2_1
X_2091_ net781 _1509_ VPWR VGND sg13g2_inv_4
XFILLER_47_872 VPWR VGND sg13g2_decap_8
XFILLER_0_53 VPWR VGND sg13g2_fill_2
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_574 VPWR VGND sg13g2_decap_8
XFILLER_34_500 VPWR VGND sg13g2_decap_8
XFILLER_0_97 VPWR VGND sg13g2_decap_8
XFILLER_34_577 VPWR VGND sg13g2_decap_8
X_2993_ _0491_ _0492_ _0344_ _0493_ VPWR VGND sg13g2_nand3_1
XFILLER_15_791 VPWR VGND sg13g2_decap_8
XFILLER_22_739 VPWR VGND sg13g2_decap_8
XFILLER_21_249 VPWR VGND sg13g2_fill_1
XFILLER_9_95 VPWR VGND sg13g2_decap_4
X_3614_ net592 _0969_ _1073_ VPWR VGND sg13g2_and2_1
X_3545_ _1010_ net680 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[6\]
+ net683 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[6\] VPWR VGND sg13g2_a22oi_1
X_3476_ net590 net571 _0944_ VPWR VGND sg13g2_nor2_1
X_2427_ VPWR _1844_ _1843_ VGND sg13g2_inv_1
X_2358_ VGND VPWR net764 net761 _1775_ _1495_ sg13g2_a21oi_1
X_2289_ _1706_ _1580_ net732 VPWR VGND sg13g2_nand2_1
X_4028_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[4\] _1399_
+ _1352_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[4\] _1400_ _1348_
+ sg13g2_a221oi_1
XFILLER_44_48 VPWR VGND sg13g2_fill_1
XFILLER_25_555 VPWR VGND sg13g2_decap_8
XFILLER_13_739 VPWR VGND sg13g2_decap_8
XFILLER_40_569 VPWR VGND sg13g2_decap_8
XFILLER_21_783 VPWR VGND sg13g2_decap_8
XFILLER_5_905 VPWR VGND sg13g2_decap_8
XFILLER_4_459 VPWR VGND sg13g2_decap_8
XFILLER_0_665 VPWR VGND sg13g2_decap_8
XFILLER_48_647 VPWR VGND sg13g2_decap_8
XFILLER_44_820 VPWR VGND sg13g2_decap_8
XFILLER_29_894 VPWR VGND sg13g2_decap_8
XFILLER_16_555 VPWR VGND sg13g2_decap_8
XFILLER_44_897 VPWR VGND sg13g2_decap_8
XFILLER_31_558 VPWR VGND sg13g2_decap_8
XFILLER_8_710 VPWR VGND sg13g2_decap_8
XFILLER_12_772 VPWR VGND sg13g2_decap_8
XFILLER_8_787 VPWR VGND sg13g2_decap_8
X_3330_ _0801_ net669 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[4\]
+ net665 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[4\] VPWR VGND sg13g2_a22oi_1
X_3261_ _0732_ _0719_ net659 VPWR VGND sg13g2_nand2_2
X_2212_ net737 _1610_ _1629_ VPWR VGND sg13g2_and2_1
X_3192_ net754 _1563_ net721 _1837_ _0663_ VPWR VGND sg13g2_or4_1
X_2143_ net760 net757 _1560_ VPWR VGND net762 sg13g2_nand3b_1
XFILLER_39_669 VPWR VGND sg13g2_decap_8
X_2074_ VPWR _1492_ net767 VGND sg13g2_inv_1
XFILLER_35_820 VPWR VGND sg13g2_decap_8
XFILLER_35_897 VPWR VGND sg13g2_decap_8
XFILLER_10_709 VPWR VGND sg13g2_decap_8
XFILLER_22_536 VPWR VGND sg13g2_decap_8
X_2976_ sap_3_inst.alu_inst.tmp\[3\] net784 _0476_ VPWR VGND sg13g2_nor2b_1
X_3528_ _0850_ _0802_ _0793_ _0994_ VPWR VGND sg13g2_a21o_1
X_3459_ _0928_ _0898_ _0914_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_809 VPWR VGND sg13g2_decap_8
XFILLER_45_617 VPWR VGND sg13g2_decap_8
XFILLER_17_308 VPWR VGND sg13g2_fill_1
XFILLER_26_831 VPWR VGND sg13g2_decap_8
XFILLER_38_1014 VPWR VGND sg13g2_decap_8
XFILLER_41_845 VPWR VGND sg13g2_decap_8
XFILLER_13_536 VPWR VGND sg13g2_decap_8
XFILLER_9_529 VPWR VGND sg13g2_decap_8
XFILLER_21_580 VPWR VGND sg13g2_decap_8
XFILLER_5_702 VPWR VGND sg13g2_decap_8
XFILLER_4_212 VPWR VGND sg13g2_fill_2
XFILLER_5_779 VPWR VGND sg13g2_decap_8
XFILLER_49_923 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_1_996 VPWR VGND sg13g2_decap_8
XFILLER_48_444 VPWR VGND sg13g2_decap_8
XFILLER_36_617 VPWR VGND sg13g2_decap_8
XFILLER_29_691 VPWR VGND sg13g2_decap_8
XFILLER_17_842 VPWR VGND sg13g2_decap_8
XFILLER_44_694 VPWR VGND sg13g2_decap_8
XFILLER_32_812 VPWR VGND sg13g2_decap_8
X_2830_ _2006_ _0333_ _2004_ _0334_ VPWR VGND sg13g2_nand3_1
XFILLER_32_889 VPWR VGND sg13g2_decap_8
X_2761_ _0288_ _0287_ VPWR VGND _1994_ sg13g2_nand2b_2
X_2692_ _0224_ net623 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[2\]
+ net630 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_8_584 VPWR VGND sg13g2_decap_8
X_4293_ net810 VGND VPWR _0150_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[4\]
+ clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3313_ _0784_ net675 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[6\]
+ net664 sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[6\] VPWR VGND sg13g2_a22oi_1
X_3244_ VGND VPWR _0715_ _1744_ _1691_ sg13g2_or2_1
XFILLER_6_1023 VPWR VGND sg13g2_decap_4
X_3175_ _0645_ net719 net739 _0646_ VPWR VGND sg13g2_a21o_1
XFILLER_39_466 VPWR VGND sg13g2_decap_8
X_2126_ VPWR _1544_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[6\]
+ VGND sg13g2_inv_1
XFILLER_23_823 VPWR VGND sg13g2_decap_8
XFILLER_35_694 VPWR VGND sg13g2_decap_8
XFILLER_10_506 VPWR VGND sg13g2_decap_8
X_2959_ _0460_ _0418_ _0458_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_606 VPWR VGND sg13g2_decap_8
XFILLER_46_937 VPWR VGND sg13g2_decap_8
XFILLER_45_414 VPWR VGND sg13g2_decap_8
XFILLER_17_149 VPWR VGND sg13g2_fill_1
XFILLER_41_642 VPWR VGND sg13g2_decap_8
XFILLER_14_856 VPWR VGND sg13g2_decap_8
XFILLER_40_185 VPWR VGND sg13g2_fill_1
XFILLER_12_1017 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_576 VPWR VGND sg13g2_decap_8
XFILLER_49_720 VPWR VGND sg13g2_decap_8
XFILLER_1_793 VPWR VGND sg13g2_decap_8
XFILLER_37_915 VPWR VGND sg13g2_decap_8
XFILLER_49_797 VPWR VGND sg13g2_decap_8
XFILLER_45_981 VPWR VGND sg13g2_decap_8
XFILLER_44_491 VPWR VGND sg13g2_decap_8
X_3931_ net798 _0154_ VPWR VGND sg13g2_inv_4
X_3862_ net585 _1004_ _1264_ VPWR VGND sg13g2_nor2_1
X_2813_ net72 sap_3_inst.out\[6\] _0185_ _0023_ VPWR VGND sg13g2_mux2_1
XFILLER_20_826 VPWR VGND sg13g2_decap_8
XFILLER_32_686 VPWR VGND sg13g2_decap_8
X_3793_ _1162_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[6\] net581
+ _0112_ VPWR VGND sg13g2_mux2_1
X_2744_ _1887_ _0271_ _1798_ _0272_ VPWR VGND sg13g2_nand3_1
XFILLER_9_893 VPWR VGND sg13g2_decap_8
X_2675_ _0207_ VPWR _0208_ VGND _1916_ net32 sg13g2_o21ai_1
XFILLER_28_1002 VPWR VGND sg13g2_decap_8
X_4345_ regFile_serial net29 VPWR VGND sg13g2_buf_8
X_4276_ net828 VGND VPWR _0133_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[3\]
+ clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3227_ _0698_ _0697_ _1645_ _1875_ _1775_ VPWR VGND sg13g2_a22oi_1
XFILLER_28_904 VPWR VGND sg13g2_decap_8
X_3158_ _1633_ _1667_ _1627_ _0629_ VPWR VGND sg13g2_nand3_1
X_2109_ VPWR _1527_ sap_3_inst.alu_inst.tmp\[5\] VGND sg13g2_inv_1
XFILLER_15_609 VPWR VGND sg13g2_decap_8
XFILLER_27_469 VPWR VGND sg13g2_decap_8
X_3089_ _0542_ _0573_ _0586_ VPWR VGND sg13g2_nor2_1
XFILLER_36_981 VPWR VGND sg13g2_decap_8
XFILLER_23_620 VPWR VGND sg13g2_decap_8
XFILLER_35_491 VPWR VGND sg13g2_decap_8
XFILLER_23_697 VPWR VGND sg13g2_decap_8
XFILLER_11_859 VPWR VGND sg13g2_decap_8
XFILLER_2_568 VPWR VGND sg13g2_decap_8
XFILLER_46_734 VPWR VGND sg13g2_decap_8
XFILLER_19_959 VPWR VGND sg13g2_decap_8
XFILLER_42_940 VPWR VGND sg13g2_decap_8
XFILLER_14_653 VPWR VGND sg13g2_decap_8
XFILLER_13_185 VPWR VGND sg13g2_fill_2
XFILLER_10_870 VPWR VGND sg13g2_decap_8
XFILLER_6_841 VPWR VGND sg13g2_decap_8
X_2460_ _1493_ _1876_ _1877_ VPWR VGND sg13g2_nor2_1
X_2391_ VPWR _1808_ _1807_ VGND sg13g2_inv_1
X_4130_ _1479_ sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos\[2\] _1315_
+ _1316_ VPWR VGND sg13g2_and3_2
XFILLER_1_590 VPWR VGND sg13g2_decap_8
X_4061_ _1313_ net53 _1429_ _0168_ VPWR VGND sg13g2_a21o_1
XFILLER_49_594 VPWR VGND sg13g2_decap_8
X_3012_ VGND VPWR _0511_ _0510_ _0506_ sg13g2_or2_1
XFILLER_3_1015 VPWR VGND sg13g2_decap_8
XFILLER_37_712 VPWR VGND sg13g2_decap_8
XFILLER_18_970 VPWR VGND sg13g2_decap_8
XFILLER_37_789 VPWR VGND sg13g2_decap_8
X_3914_ _1297_ _1300_ _1301_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_623 VPWR VGND sg13g2_decap_8
XFILLER_33_995 VPWR VGND sg13g2_decap_8
X_3845_ net652 _1222_ _1250_ _1251_ VPWR VGND sg13g2_nor3_1
X_3776_ VGND VPWR net655 _1043_ _1208_ net612 sg13g2_a21oi_1
XFILLER_9_690 VPWR VGND sg13g2_decap_8
X_2727_ _0257_ _0255_ _0256_ VPWR VGND sg13g2_nand2_1
X_2658_ _2065_ net618 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[3\]
+ net621 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[3\] VPWR VGND
+ sg13g2_a22oi_1
X_2589_ _1723_ VPWR _1998_ VGND net728 _1762_ sg13g2_o21ai_1
X_4328_ net817 VGND VPWR net799 u_ser.state\[0\] clknet_3_0__leaf_clk sg13g2_dfrbpq_2
X_4259_ net827 VGND VPWR _0116_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[2\]
+ clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_28_701 VPWR VGND sg13g2_decap_8
XFILLER_28_778 VPWR VGND sg13g2_decap_8
XFILLER_43_759 VPWR VGND sg13g2_decap_8
XFILLER_24_962 VPWR VGND sg13g2_decap_8
XFILLER_11_656 VPWR VGND sg13g2_decap_8
XFILLER_23_494 VPWR VGND sg13g2_decap_8
XFILLER_3_833 VPWR VGND sg13g2_decap_8
Xclkbuf_5_6__f_sap_3_inst.alu_inst.clk_regs clknet_4_3_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
Xfanout680 net682 net680 VPWR VGND sg13g2_buf_8
Xfanout691 _0359_ net691 VPWR VGND sg13g2_buf_8
XFILLER_46_531 VPWR VGND sg13g2_decap_8
XFILLER_19_756 VPWR VGND sg13g2_decap_8
XFILLER_33_203 VPWR VGND sg13g2_fill_1
XFILLER_34_759 VPWR VGND sg13g2_decap_8
XFILLER_15_973 VPWR VGND sg13g2_decap_8
XFILLER_18_1012 VPWR VGND sg13g2_decap_8
XFILLER_30_910 VPWR VGND sg13g2_decap_8
X_3630_ _0080_ _1085_ _1086_ net584 _1544_ VPWR VGND sg13g2_a22oi_1
XFILLER_30_987 VPWR VGND sg13g2_decap_8
X_3561_ _0991_ _0950_ _1017_ _1026_ VPWR VGND sg13g2_a21o_1
X_2512_ _1924_ _1926_ _1923_ _1927_ VPWR VGND sg13g2_nand3_1
X_3492_ _0959_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[4\] net596
+ VPWR VGND sg13g2_nand2_1
X_2443_ net696 net666 net707 _1844_ _1860_ VPWR VGND sg13g2_and4_1
X_2374_ _1591_ VPWR _1791_ VGND net721 _1769_ sg13g2_o21ai_1
X_4113_ u_ser.state\[0\] _1489_ _1465_ VPWR VGND sg13g2_nor2_2
XFILLER_29_509 VPWR VGND sg13g2_decap_8
XFILLER_49_391 VPWR VGND sg13g2_decap_8
X_4044_ VGND VPWR sap_3_inst.reg_file_inst.array_serializer_inst.data\[1\]\[6\] _1348_
+ _1414_ net794 sg13g2_a21oi_1
XFILLER_25_737 VPWR VGND sg13g2_decap_8
XFILLER_37_586 VPWR VGND sg13g2_decap_8
XFILLER_33_792 VPWR VGND sg13g2_decap_8
XFILLER_21_965 VPWR VGND sg13g2_decap_8
XFILLER_32_280 VPWR VGND sg13g2_fill_2
X_3828_ _1237_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[5\] net634
+ _0127_ VPWR VGND sg13g2_mux2_1
XFILLER_20_497 VPWR VGND sg13g2_decap_8
X_3759_ net594 VPWR _1193_ VGND net676 _0995_ sg13g2_o21ai_1
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_48_829 VPWR VGND sg13g2_decap_8
XFILLER_28_575 VPWR VGND sg13g2_decap_8
XFILLER_16_737 VPWR VGND sg13g2_decap_8
XFILLER_43_556 VPWR VGND sg13g2_decap_8
XFILLER_30_217 VPWR VGND sg13g2_fill_2
XFILLER_12_954 VPWR VGND sg13g2_decap_8
XFILLER_8_969 VPWR VGND sg13g2_decap_8
XFILLER_23_94 VPWR VGND sg13g2_fill_2
XFILLER_3_630 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_fill_1
XFILLER_47_851 VPWR VGND sg13g2_decap_8
X_2090_ VPWR _1508_ net793 VGND sg13g2_inv_1
XFILLER_19_553 VPWR VGND sg13g2_decap_8
XFILLER_22_718 VPWR VGND sg13g2_decap_8
XFILLER_34_556 VPWR VGND sg13g2_decap_8
X_2992_ VGND VPWR _0492_ _0490_ _0459_ sg13g2_or2_1
XFILLER_15_770 VPWR VGND sg13g2_decap_8
XFILLER_30_784 VPWR VGND sg13g2_decap_8
XFILLER_31_1020 VPWR VGND sg13g2_decap_8
X_3613_ _0077_ _1070_ _1072_ net583 _1499_ VPWR VGND sg13g2_a22oi_1
X_3544_ _0982_ VPWR _0071_ VGND _1003_ _1008_ sg13g2_o21ai_1
X_3475_ _0891_ _0915_ _0865_ _0943_ VPWR VGND _0941_ sg13g2_nand4_1
X_2426_ _1832_ _1842_ _1843_ VPWR VGND sg13g2_and2_1
X_2357_ VPWR VGND _1595_ net719 _1770_ net730 _1774_ net734 sg13g2_a221oi_1
X_2288_ _1491_ _1683_ _1705_ VPWR VGND sg13g2_nor2_2
X_4027_ _1395_ _1397_ _1394_ _1399_ VPWR VGND _1398_ sg13g2_nand4_1
XFILLER_25_534 VPWR VGND sg13g2_decap_8
XFILLER_38_895 VPWR VGND sg13g2_decap_8
XFILLER_13_718 VPWR VGND sg13g2_decap_8
XFILLER_40_548 VPWR VGND sg13g2_decap_8
XFILLER_12_228 VPWR VGND sg13g2_fill_2
XFILLER_21_762 VPWR VGND sg13g2_decap_8
XFILLER_20_283 VPWR VGND sg13g2_fill_2
XFILLER_4_405 VPWR VGND sg13g2_fill_1
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_48_626 VPWR VGND sg13g2_decap_8
XFILLER_29_873 VPWR VGND sg13g2_decap_8
XFILLER_16_534 VPWR VGND sg13g2_decap_8
XFILLER_44_876 VPWR VGND sg13g2_decap_8
XFILLER_31_537 VPWR VGND sg13g2_decap_8
XFILLER_12_751 VPWR VGND sg13g2_decap_8
XFILLER_15_1015 VPWR VGND sg13g2_decap_8
XFILLER_11_272 VPWR VGND sg13g2_fill_2
XFILLER_8_766 VPWR VGND sg13g2_decap_8
X_3260_ _0731_ net659 VPWR VGND sg13g2_inv_2
X_2211_ _1493_ _1623_ _1628_ VPWR VGND net749 sg13g2_nand3b_1
X_3191_ net740 VPWR _0662_ VGND _0655_ _0661_ sg13g2_o21ai_1
XFILLER_22_4 VPWR VGND sg13g2_fill_1
X_2142_ net763 net752 _1559_ VPWR VGND sg13g2_nor2_1
XFILLER_22_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_648 VPWR VGND sg13g2_decap_8
X_2073_ _1491_ net747 VPWR VGND sg13g2_inv_2
XFILLER_26_309 VPWR VGND sg13g2_fill_1
XFILLER_35_876 VPWR VGND sg13g2_decap_8
XFILLER_22_515 VPWR VGND sg13g2_decap_8
X_2975_ VPWR _0475_ _0474_ VGND sg13g2_inv_1
XFILLER_30_581 VPWR VGND sg13g2_decap_8
X_3527_ VGND VPWR _0992_ _0993_ _0991_ _0950_ sg13g2_a21oi_2
X_3458_ _0891_ _0915_ _0865_ _0927_ VPWR VGND sg13g2_nand3_1
X_2409_ VGND VPWR _1820_ _1821_ _1826_ _1602_ sg13g2_a21oi_1
X_3389_ VGND VPWR _0860_ _0847_ _0836_ sg13g2_or2_1
XFILLER_39_49 VPWR VGND sg13g2_fill_1
XFILLER_26_810 VPWR VGND sg13g2_decap_8
XFILLER_38_692 VPWR VGND sg13g2_decap_8
XFILLER_41_824 VPWR VGND sg13g2_decap_8
XFILLER_13_515 VPWR VGND sg13g2_decap_8
XFILLER_26_887 VPWR VGND sg13g2_decap_8
XFILLER_9_508 VPWR VGND sg13g2_decap_8
XFILLER_25_386 VPWR VGND sg13g2_fill_1
XFILLER_5_758 VPWR VGND sg13g2_decap_8
XFILLER_49_902 VPWR VGND sg13g2_decap_8
XFILLER_1_975 VPWR VGND sg13g2_decap_8
XFILLER_48_423 VPWR VGND sg13g2_decap_8
XFILLER_49_979 VPWR VGND sg13g2_decap_8
XFILLER_17_821 VPWR VGND sg13g2_decap_8
XFILLER_29_670 VPWR VGND sg13g2_decap_8
XFILLER_44_673 VPWR VGND sg13g2_decap_8
XFILLER_17_898 VPWR VGND sg13g2_decap_8
XFILLER_32_868 VPWR VGND sg13g2_decap_8
X_2760_ VGND VPWR _1608_ _1731_ _0287_ _1620_ sg13g2_a21oi_1
XFILLER_8_563 VPWR VGND sg13g2_decap_8
X_2691_ _0223_ net617 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[2\]
+ net711 sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[2\] VPWR VGND
+ sg13g2_a22oi_1
X_3312_ _0783_ net669 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[6\]
+ net680 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[6\] VPWR VGND sg13g2_a22oi_1
X_4292_ net831 VGND VPWR _0149_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[3\]
+ clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_6_1002 VPWR VGND sg13g2_decap_8
X_3243_ _0670_ net735 _1709_ _0714_ VPWR VGND sg13g2_a21o_1
X_3174_ net759 VPWR _0645_ VGND _0643_ _0644_ sg13g2_o21ai_1
XFILLER_48_990 VPWR VGND sg13g2_decap_8
X_2125_ VPWR _1543_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[6\]
+ VGND sg13g2_inv_1
XFILLER_26_117 VPWR VGND sg13g2_fill_2
XFILLER_23_802 VPWR VGND sg13g2_decap_8
XFILLER_35_673 VPWR VGND sg13g2_decap_8
XFILLER_23_879 VPWR VGND sg13g2_decap_8
X_2958_ _0419_ _0458_ _0459_ VPWR VGND sg13g2_nor2_1
X_2889_ _0361_ VPWR _0392_ VGND net790 sap_3_inst.alu_inst.tmp\[1\] sg13g2_o21ai_1
XFILLER_46_916 VPWR VGND sg13g2_decap_8
XFILLER_26_684 VPWR VGND sg13g2_decap_8
XFILLER_41_621 VPWR VGND sg13g2_decap_8
XFILLER_14_835 VPWR VGND sg13g2_decap_8
XFILLER_41_698 VPWR VGND sg13g2_decap_8
XFILLER_5_555 VPWR VGND sg13g2_decap_8
XFILLER_1_772 VPWR VGND sg13g2_decap_8
XFILLER_0_260 VPWR VGND sg13g2_fill_1
XFILLER_49_776 VPWR VGND sg13g2_decap_8
XFILLER_48_297 VPWR VGND sg13g2_decap_8
XFILLER_45_960 VPWR VGND sg13g2_decap_8
X_3930_ VGND VPWR _1313_ sap_3_inst.reg_file_inst.array_serializer_inst.state\[1\]
+ sap_3_inst.reg_file_inst.array_serializer_inst.state\[0\] sg13g2_or2_1
XFILLER_44_470 VPWR VGND sg13g2_decap_8
XFILLER_17_695 VPWR VGND sg13g2_decap_8
XFILLER_20_805 VPWR VGND sg13g2_decap_8
XFILLER_32_665 VPWR VGND sg13g2_decap_8
X_3861_ _0990_ VPWR _1263_ VGND net571 net573 sg13g2_o21ai_1
X_3792_ _1217_ VPWR _0111_ VGND _1081_ net580 sg13g2_o21ai_1
X_2812_ net76 sap_3_inst.out\[5\] _0185_ _0022_ VPWR VGND sg13g2_mux2_1
XFILLER_31_175 VPWR VGND sg13g2_fill_1
X_2743_ _1730_ _1748_ _1754_ net719 _0271_ VPWR VGND sg13g2_nor4_1
XFILLER_9_872 VPWR VGND sg13g2_decap_8
X_2674_ _0207_ _1916_ net774 VPWR VGND sg13g2_nand2b_1
X_4344_ sap_3_outputReg_start_sync net28 VPWR VGND sg13g2_buf_1
X_4275_ net827 VGND VPWR _0132_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[2\]
+ clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3226_ _1634_ VPWR _0697_ VGND _1656_ _1693_ sg13g2_o21ai_1
X_3157_ VGND VPWR _1585_ _1914_ _0065_ _0628_ sg13g2_a21oi_1
X_2108_ VPWR _1526_ sap_3_inst.alu_inst.act\[7\] VGND sg13g2_inv_1
XFILLER_27_448 VPWR VGND sg13g2_decap_8
X_3088_ _0579_ _0580_ _0581_ _0584_ _0585_ VPWR VGND sg13g2_and4_1
XFILLER_36_960 VPWR VGND sg13g2_decap_8
XFILLER_23_676 VPWR VGND sg13g2_decap_8
XFILLER_11_838 VPWR VGND sg13g2_decap_8
XFILLER_2_547 VPWR VGND sg13g2_decap_8
XFILLER_46_713 VPWR VGND sg13g2_decap_8
XFILLER_19_938 VPWR VGND sg13g2_decap_8
XFILLER_45_223 VPWR VGND sg13g2_fill_2
XFILLER_18_459 VPWR VGND sg13g2_fill_1
XFILLER_14_632 VPWR VGND sg13g2_decap_8
XFILLER_26_481 VPWR VGND sg13g2_decap_8
XFILLER_42_996 VPWR VGND sg13g2_decap_8
XFILLER_41_495 VPWR VGND sg13g2_decap_8
XFILLER_9_168 VPWR VGND sg13g2_fill_2
XFILLER_6_820 VPWR VGND sg13g2_decap_8
XFILLER_5_330 VPWR VGND sg13g2_fill_1
XFILLER_6_897 VPWR VGND sg13g2_decap_8
XFILLER_3_10 VPWR VGND sg13g2_fill_1
X_2390_ _1556_ _1606_ _1806_ _1807_ VPWR VGND sg13g2_or3_1
X_4060_ VPWR VGND _1428_ net798 _1422_ _1545_ _1429_ net794 sg13g2_a221oi_1
XFILLER_49_573 VPWR VGND sg13g2_decap_8
X_3011_ _0361_ _0509_ _0510_ VPWR VGND sg13g2_nor2_1
XFILLER_36_223 VPWR VGND sg13g2_decap_4
XFILLER_37_768 VPWR VGND sg13g2_decap_8
XFILLER_25_919 VPWR VGND sg13g2_decap_8
XFILLER_17_492 VPWR VGND sg13g2_decap_8
X_3913_ _1299_ VPWR _1300_ VGND _0968_ _1298_ sg13g2_o21ai_1
XFILLER_33_974 VPWR VGND sg13g2_decap_8
XFILLER_20_602 VPWR VGND sg13g2_decap_8
X_3844_ net585 _1249_ _1250_ VPWR VGND sg13g2_nor2_1
XFILLER_20_679 VPWR VGND sg13g2_decap_8
X_3775_ _1206_ VPWR _1207_ VGND net24 net602 sg13g2_o21ai_1
X_2726_ _0256_ net625 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[0\]
+ net629 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2657_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[3\] net632
+ net616 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[3\] _2064_ net712
+ sg13g2_a221oi_1
X_2588_ _1997_ _1592_ _1612_ VPWR VGND sg13g2_nand2_1
X_4327_ net824 VGND VPWR _0184_ sap_3_inst.alu_inst.act\[7\] clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4258_ net804 VGND VPWR _0115_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[1\]
+ clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3209_ _1639_ _1699_ _0680_ VPWR VGND sg13g2_nor2_1
X_4189_ net822 VGND VPWR _0046_ sap_3_inst.out\[5\] clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
XFILLER_28_757 VPWR VGND sg13g2_decap_8
XFILLER_16_919 VPWR VGND sg13g2_decap_8
XFILLER_43_738 VPWR VGND sg13g2_decap_8
XFILLER_42_259 VPWR VGND sg13g2_fill_2
XFILLER_24_941 VPWR VGND sg13g2_decap_8
XFILLER_23_473 VPWR VGND sg13g2_decap_8
XFILLER_11_635 VPWR VGND sg13g2_decap_8
XFILLER_10_156 VPWR VGND sg13g2_fill_1
XFILLER_7_639 VPWR VGND sg13g2_decap_8
XFILLER_6_105 VPWR VGND sg13g2_fill_1
XFILLER_3_812 VPWR VGND sg13g2_decap_8
XFILLER_3_889 VPWR VGND sg13g2_decap_8
XFILLER_46_510 VPWR VGND sg13g2_decap_8
Xfanout692 _0357_ net692 VPWR VGND sg13g2_buf_8
Xfanout670 _0763_ net670 VPWR VGND sg13g2_buf_8
Xfanout681 net682 net681 VPWR VGND sg13g2_buf_8
XFILLER_19_735 VPWR VGND sg13g2_decap_8
XFILLER_46_587 VPWR VGND sg13g2_decap_8
XFILLER_34_738 VPWR VGND sg13g2_decap_8
XFILLER_15_952 VPWR VGND sg13g2_decap_8
XFILLER_42_793 VPWR VGND sg13g2_decap_8
XFILLER_30_966 VPWR VGND sg13g2_decap_8
X_3560_ _0991_ _1017_ _0950_ _1025_ VPWR VGND sg13g2_nand3_1
X_2511_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[6\] net631
+ net621 sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[6\] _1926_ net624
+ sg13g2_a221oi_1
XFILLER_6_694 VPWR VGND sg13g2_decap_8
XFILLER_5_160 VPWR VGND sg13g2_fill_1
X_3491_ VGND VPWR _1497_ net597 _0069_ _0958_ sg13g2_a21oi_1
X_2442_ _1807_ net666 net707 _1844_ _1859_ VPWR VGND sg13g2_and4_1
X_2373_ _1569_ VPWR _1790_ VGND _1771_ _1789_ sg13g2_o21ai_1
XFILLER_38_2 VPWR VGND sg13g2_fill_1
X_4112_ _0184_ _1463_ _1464_ net579 _1526_ VPWR VGND sg13g2_a22oi_1
XFILLER_25_1017 VPWR VGND sg13g2_decap_8
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
X_4043_ _1413_ _1353_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[6\]
+ _1352_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_49_370 VPWR VGND sg13g2_decap_8
XFILLER_25_716 VPWR VGND sg13g2_decap_8
XFILLER_37_565 VPWR VGND sg13g2_decap_8
XFILLER_33_771 VPWR VGND sg13g2_decap_8
XFILLER_21_944 VPWR VGND sg13g2_decap_8
X_3827_ _1078_ VPWR _1237_ VGND net588 _1009_ sg13g2_o21ai_1
XFILLER_20_476 VPWR VGND sg13g2_decap_8
X_3758_ _1192_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[4\]\[5\] net656
+ VPWR VGND sg13g2_nand2_1
X_2709_ _0239_ net633 sap_3_inst.reg_file_inst.array_serializer_inst.data\[0\]\[0\]
+ VPWR VGND sg13g2_nand2b_1
X_3689_ _1138_ _0786_ _0863_ VPWR VGND sg13g2_nand2_1
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_48_808 VPWR VGND sg13g2_decap_8
XFILLER_47_307 VPWR VGND sg13g2_fill_1
Xclkbuf_5_19__f_sap_3_inst.alu_inst.clk_regs clknet_4_9_0_sap_3_inst.alu_inst.clk_regs
+ clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs VPWR VGND sg13g2_buf_8
XFILLER_16_716 VPWR VGND sg13g2_decap_8
XFILLER_28_554 VPWR VGND sg13g2_decap_8
XFILLER_43_535 VPWR VGND sg13g2_decap_8
XFILLER_31_719 VPWR VGND sg13g2_decap_8
XFILLER_12_933 VPWR VGND sg13g2_decap_8
XFILLER_23_270 VPWR VGND sg13g2_fill_1
XFILLER_8_948 VPWR VGND sg13g2_decap_8
XFILLER_3_686 VPWR VGND sg13g2_decap_8
XFILLER_47_830 VPWR VGND sg13g2_decap_8
XFILLER_19_532 VPWR VGND sg13g2_decap_8
XFILLER_0_1008 VPWR VGND sg13g2_decap_8
XFILLER_46_384 VPWR VGND sg13g2_decap_8
XFILLER_34_535 VPWR VGND sg13g2_decap_8
X_2991_ _0491_ _0459_ _0490_ VPWR VGND sg13g2_nand2_1
XFILLER_42_590 VPWR VGND sg13g2_decap_8
XFILLER_9_64 VPWR VGND sg13g2_fill_1
XFILLER_30_763 VPWR VGND sg13g2_decap_8
X_3612_ net583 _1071_ _1072_ VPWR VGND sg13g2_nor2_1
X_3543_ _1009_ _0793_ _0866_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_0 VPWR VGND sg13g2_fill_2
XFILLER_6_491 VPWR VGND sg13g2_decap_8
X_3474_ _0940_ VPWR _0942_ VGND _0825_ _0927_ sg13g2_o21ai_1
X_2425_ _1840_ _1841_ _1569_ _1842_ VPWR VGND sg13g2_nand3_1
X_2356_ net729 _1662_ _1773_ VPWR VGND sg13g2_nor2_1
X_2287_ _1612_ _1703_ _1704_ VPWR VGND sg13g2_and2_1
X_4026_ _1398_ _1351_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[4\]
+ _1350_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[4\] VPWR VGND sg13g2_a22oi_1
XFILLER_38_874 VPWR VGND sg13g2_decap_8
XFILLER_25_513 VPWR VGND sg13g2_decap_8
XFILLER_40_527 VPWR VGND sg13g2_decap_8
XFILLER_21_741 VPWR VGND sg13g2_decap_8
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_20_295 VPWR VGND sg13g2_fill_2
XFILLER_0_623 VPWR VGND sg13g2_decap_8
XFILLER_48_605 VPWR VGND sg13g2_decap_8
XFILLER_29_852 VPWR VGND sg13g2_decap_8
XFILLER_16_513 VPWR VGND sg13g2_decap_8
XFILLER_28_373 VPWR VGND sg13g2_fill_2
XFILLER_44_855 VPWR VGND sg13g2_decap_8
XFILLER_31_516 VPWR VGND sg13g2_decap_8
XFILLER_12_730 VPWR VGND sg13g2_decap_8
XFILLER_34_94 VPWR VGND sg13g2_fill_2
XFILLER_8_745 VPWR VGND sg13g2_decap_8
XFILLER_11_262 VPWR VGND sg13g2_fill_1
XFILLER_7_266 VPWR VGND sg13g2_fill_1
XFILLER_4_984 VPWR VGND sg13g2_decap_8
XFILLER_3_483 VPWR VGND sg13g2_decap_8
X_2210_ net762 _1624_ _1625_ _1627_ VPWR VGND sg13g2_nor3_2
X_3190_ _0658_ _0660_ _0656_ _0661_ VPWR VGND sg13g2_nand3_1
XFILLER_39_627 VPWR VGND sg13g2_decap_8
X_2141_ _1558_ net759 net758 VPWR VGND sg13g2_nand2_2
X_2072_ VPWR _1490_ u_ser.bit_pos\[2\] VGND sg13g2_inv_1
XFILLER_38_148 VPWR VGND sg13g2_fill_2
XFILLER_35_855 VPWR VGND sg13g2_decap_8
X_2974_ _0474_ net781 sap_3_inst.alu_inst.tmp\[4\] VPWR VGND sg13g2_xnor2_1
XFILLER_30_560 VPWR VGND sg13g2_decap_8
X_3526_ VGND VPWR _0950_ net574 _0992_ _0990_ sg13g2_a21oi_1
X_3457_ VPWR VGND _0922_ _0925_ _0921_ net594 _0926_ _0920_ sg13g2_a221oi_1
X_2408_ _1825_ _1820_ _1821_ _1824_ VPWR VGND sg13g2_and3_1
X_3388_ _0859_ _0841_ _0846_ _0835_ _0830_ VPWR VGND sg13g2_a22oi_1
X_2339_ _1747_ _1751_ _1695_ _1756_ VPWR VGND _1755_ sg13g2_nand4_1
XFILLER_29_148 VPWR VGND sg13g2_fill_1
X_4009_ _1382_ VPWR _0163_ VGND _1549_ _0154_ sg13g2_o21ai_1
XFILLER_38_671 VPWR VGND sg13g2_decap_8
XFILLER_26_866 VPWR VGND sg13g2_decap_8
XFILLER_41_803 VPWR VGND sg13g2_decap_8
XFILLER_5_737 VPWR VGND sg13g2_decap_8
XFILLER_45_1009 VPWR VGND sg13g2_decap_8
XFILLER_1_954 VPWR VGND sg13g2_decap_8
XFILLER_48_402 VPWR VGND sg13g2_decap_8
XFILLER_49_958 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_48_479 VPWR VGND sg13g2_decap_8
XFILLER_17_800 VPWR VGND sg13g2_decap_8
XFILLER_44_652 VPWR VGND sg13g2_decap_8
XFILLER_17_877 VPWR VGND sg13g2_decap_8
XFILLER_32_847 VPWR VGND sg13g2_decap_8
XFILLER_40_891 VPWR VGND sg13g2_decap_8
XFILLER_8_542 VPWR VGND sg13g2_decap_8
X_2690_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[2\] net620
+ net615 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[2\] _0222_ net625
+ sg13g2_a221oi_1
XFILLER_6_10 VPWR VGND sg13g2_fill_1
XFILLER_6_76 VPWR VGND sg13g2_fill_2
XFILLER_6_65 VPWR VGND sg13g2_decap_8
XFILLER_6_54 VPWR VGND sg13g2_fill_1
X_3311_ _0782_ net638 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[6\]
+ net641 sap_3_inst.reg_file_inst.array_serializer_inst.data\[2\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_4_781 VPWR VGND sg13g2_decap_8
X_4291_ net819 VGND VPWR _0148_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[2\]
+ clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3242_ VGND VPWR _0713_ net689 _0667_ sg13g2_or2_1
XFILLER_39_402 VPWR VGND sg13g2_fill_1
X_3173_ _1573_ net729 _1616_ _0644_ VPWR VGND sg13g2_nor3_2
X_2124_ VPWR _1542_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[6\]
+ VGND sg13g2_inv_1
XFILLER_35_652 VPWR VGND sg13g2_decap_8
XFILLER_23_858 VPWR VGND sg13g2_decap_8
X_2957_ _0458_ _0439_ _0457_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_880 VPWR VGND sg13g2_decap_8
X_2888_ VGND VPWR _0391_ _0379_ _0346_ sg13g2_or2_1
XFILLER_2_729 VPWR VGND sg13g2_decap_8
X_3509_ _0971_ _0972_ _0975_ _0976_ VPWR VGND sg13g2_nor3_1
XFILLER_39_991 VPWR VGND sg13g2_decap_8
XFILLER_45_449 VPWR VGND sg13g2_decap_8
XFILLER_41_600 VPWR VGND sg13g2_decap_8
XFILLER_14_814 VPWR VGND sg13g2_decap_8
XFILLER_26_663 VPWR VGND sg13g2_decap_8
XFILLER_41_677 VPWR VGND sg13g2_decap_8
XFILLER_5_534 VPWR VGND sg13g2_decap_8
XFILLER_1_751 VPWR VGND sg13g2_decap_8
XFILLER_49_755 VPWR VGND sg13g2_decap_8
XFILLER_17_674 VPWR VGND sg13g2_decap_8
XFILLER_31_110 VPWR VGND sg13g2_fill_1
X_3860_ _0134_ _1259_ _1262_ net652 _1531_ VPWR VGND sg13g2_a22oi_1
XFILLER_32_644 VPWR VGND sg13g2_decap_8
X_3791_ _1217_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[5\] net581
+ VPWR VGND sg13g2_nand2_1
X_2811_ net67 sap_3_inst.out\[4\] net799 _0021_ VPWR VGND sg13g2_mux2_1
XFILLER_9_851 VPWR VGND sg13g2_decap_8
X_2742_ _0270_ sap_3_inst.alu_flags\[0\] _0238_ _0025_ VPWR VGND sg13g2_mux2_1
XFILLER_8_350 VPWR VGND sg13g2_fill_2
X_2673_ _0204_ _0205_ _0196_ net20 VPWR VGND _0206_ sg13g2_nand4_1
X_4343_ sap_3_outputReg_serial net27 VPWR VGND sg13g2_buf_1
X_4274_ net805 VGND VPWR _0131_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3225_ _0696_ net758 _1886_ VPWR VGND sg13g2_nand2_1
X_3156_ net754 net718 _0628_ VPWR VGND sg13g2_nor2_1
XFILLER_28_939 VPWR VGND sg13g2_decap_8
X_3087_ _0582_ _0583_ _0584_ VPWR VGND sg13g2_nor2_1
X_2107_ VPWR _1525_ sap_3_inst.alu_inst.act\[0\] VGND sg13g2_inv_1
XFILLER_23_655 VPWR VGND sg13g2_decap_8
XFILLER_11_817 VPWR VGND sg13g2_decap_8
X_3989_ _1364_ VPWR _0161_ VGND _1362_ _1363_ sg13g2_o21ai_1
XFILLER_2_526 VPWR VGND sg13g2_decap_8
Xfanout830 net832 net830 VPWR VGND sg13g2_buf_8
XFILLER_45_202 VPWR VGND sg13g2_fill_2
XFILLER_18_416 VPWR VGND sg13g2_fill_1
XFILLER_19_917 VPWR VGND sg13g2_decap_8
XFILLER_46_769 VPWR VGND sg13g2_decap_8
XFILLER_14_611 VPWR VGND sg13g2_decap_8
XFILLER_26_460 VPWR VGND sg13g2_decap_8
XFILLER_27_994 VPWR VGND sg13g2_decap_8
XFILLER_42_975 VPWR VGND sg13g2_decap_8
XFILLER_41_474 VPWR VGND sg13g2_decap_8
XFILLER_14_688 VPWR VGND sg13g2_decap_8
XFILLER_13_187 VPWR VGND sg13g2_fill_1
XFILLER_6_876 VPWR VGND sg13g2_decap_8
XFILLER_3_77 VPWR VGND sg13g2_fill_1
XFILLER_49_552 VPWR VGND sg13g2_decap_8
X_3010_ _0355_ _0507_ _0509_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_747 VPWR VGND sg13g2_decap_8
X_3912_ VGND VPWR net13 _1286_ _1299_ _0975_ sg13g2_a21oi_1
XFILLER_33_953 VPWR VGND sg13g2_decap_8
X_3843_ _1249_ _0865_ _0891_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_658 VPWR VGND sg13g2_decap_8
X_3774_ _1206_ _0306_ net602 VPWR VGND sg13g2_nand2_1
X_2725_ _0255_ net619 sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[0\]
+ net623 sap_3_inst.reg_file_inst.array_serializer_inst.data\[3\]\[0\] VPWR VGND sg13g2_a22oi_1
X_2656_ _2061_ _2062_ _2060_ _2063_ VPWR VGND sg13g2_nand3_1
X_2587_ _1993_ VPWR _1996_ VGND _1602_ _1995_ sg13g2_o21ai_1
X_4326_ net823 VGND VPWR _0183_ sap_3_inst.alu_inst.act\[6\] clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_4257_ net827 VGND VPWR _0114_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[0\]
+ clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3208_ _0679_ _0673_ _0675_ _0678_ VPWR VGND sg13g2_and3_1
X_4188_ net822 VGND VPWR _0045_ sap_3_inst.out\[4\] clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs
+ sg13g2_dfrbpq_1
X_3139_ _0620_ sap_3_inst.alu_inst.tmp\[6\] net700 VPWR VGND sg13g2_nand2_1
XFILLER_28_736 VPWR VGND sg13g2_decap_8
XFILLER_43_717 VPWR VGND sg13g2_decap_8
XFILLER_24_920 VPWR VGND sg13g2_decap_8
XFILLER_11_614 VPWR VGND sg13g2_decap_8
XFILLER_23_452 VPWR VGND sg13g2_decap_8
XFILLER_24_997 VPWR VGND sg13g2_decap_8
XFILLER_7_618 VPWR VGND sg13g2_decap_8
XFILLER_6_117 VPWR VGND sg13g2_fill_2
XFILLER_3_868 VPWR VGND sg13g2_decap_8
Xfanout660 net661 net660 VPWR VGND sg13g2_buf_8
Xfanout693 _0330_ net693 VPWR VGND sg13g2_buf_2
XFILLER_19_714 VPWR VGND sg13g2_decap_8
Xfanout682 _0750_ net682 VPWR VGND sg13g2_buf_8
Xfanout671 net674 net671 VPWR VGND sg13g2_buf_8
XFILLER_46_566 VPWR VGND sg13g2_decap_8
XFILLER_34_717 VPWR VGND sg13g2_decap_8
XFILLER_15_931 VPWR VGND sg13g2_decap_8
XFILLER_18_279 VPWR VGND sg13g2_fill_2
XFILLER_27_791 VPWR VGND sg13g2_decap_8
XFILLER_14_441 VPWR VGND sg13g2_fill_1
XFILLER_42_772 VPWR VGND sg13g2_decap_8
XFILLER_30_945 VPWR VGND sg13g2_decap_8
X_2510_ _1920_ _1921_ _1919_ _1925_ VPWR VGND _1922_ sg13g2_nand4_1
X_3490_ net597 _0948_ _0954_ _0956_ _0958_ VPWR VGND sg13g2_nor4_1
XFILLER_6_673 VPWR VGND sg13g2_decap_8
X_2441_ VPWR VGND sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[7\] net631
+ net621 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[7\] _1858_ net711
+ sg13g2_a221oi_1
X_2372_ _1778_ _1781_ _1785_ _1788_ _1789_ VPWR VGND sg13g2_nor4_1
XFILLER_2_890 VPWR VGND sg13g2_decap_8
X_4111_ VGND VPWR net773 _1439_ _1464_ net579 sg13g2_a21oi_1
X_4042_ _1412_ _1350_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[6\]
+ net797 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_37_544 VPWR VGND sg13g2_decap_8
XFILLER_40_709 VPWR VGND sg13g2_decap_8
XFILLER_21_923 VPWR VGND sg13g2_decap_8
XFILLER_33_750 VPWR VGND sg13g2_decap_8
XFILLER_32_282 VPWR VGND sg13g2_fill_1
X_3826_ _1160_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[4\] net634
+ _0126_ VPWR VGND sg13g2_mux2_1
X_3757_ _0102_ _1120_ _1191_ net656 _1533_ VPWR VGND sg13g2_a22oi_1
X_2708_ _2003_ VPWR _0238_ VGND _1492_ net754 sg13g2_o21ai_1
X_3688_ VGND VPWR net570 _1097_ _1137_ _1136_ sg13g2_a21oi_1
XFILLER_0_805 VPWR VGND sg13g2_decap_8
X_2639_ _2048_ net615 sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[1\]
+ net624 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[1\] VPWR VGND sg13g2_a22oi_1
X_4309_ net835 VGND VPWR _0166_ sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg\[5\]
+ clknet_3_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_47_319 VPWR VGND sg13g2_decap_8
XFILLER_28_533 VPWR VGND sg13g2_decap_8
XFILLER_43_514 VPWR VGND sg13g2_decap_8
XFILLER_12_912 VPWR VGND sg13g2_decap_8
XFILLER_30_219 VPWR VGND sg13g2_fill_1
XFILLER_24_794 VPWR VGND sg13g2_decap_8
XFILLER_8_927 VPWR VGND sg13g2_decap_8
XFILLER_7_415 VPWR VGND sg13g2_fill_1
XFILLER_12_989 VPWR VGND sg13g2_decap_8
XFILLER_7_437 VPWR VGND sg13g2_fill_1
XFILLER_11_488 VPWR VGND sg13g2_decap_8
XFILLER_48_1018 VPWR VGND sg13g2_decap_8
XFILLER_3_665 VPWR VGND sg13g2_decap_8
XFILLER_39_809 VPWR VGND sg13g2_decap_8
XFILLER_19_511 VPWR VGND sg13g2_decap_8
XFILLER_47_886 VPWR VGND sg13g2_decap_8
XFILLER_46_363 VPWR VGND sg13g2_decap_8
XFILLER_0_67 VPWR VGND sg13g2_decap_8
XFILLER_19_588 VPWR VGND sg13g2_decap_8
XFILLER_34_514 VPWR VGND sg13g2_decap_8
X_2990_ _0490_ _0474_ _0489_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_742 VPWR VGND sg13g2_decap_8
X_3611_ net611 _0946_ _1071_ VPWR VGND sg13g2_and2_1
XFILLER_7_982 VPWR VGND sg13g2_decap_8
XFILLER_6_470 VPWR VGND sg13g2_decap_8
X_3542_ _0742_ VPWR _1008_ VGND net586 _1006_ sg13g2_o21ai_1
X_3473_ VPWR _0941_ _0940_ VGND sg13g2_inv_1
XFILLER_9_1012 VPWR VGND sg13g2_decap_8
X_2424_ VGND VPWR net771 _1834_ _1841_ _1838_ sg13g2_a21oi_1
X_2355_ _1636_ _1656_ net720 _1772_ VPWR VGND sg13g2_nor3_1
XFILLER_36_0 VPWR VGND sg13g2_fill_2
X_2286_ net758 _1562_ _1573_ _1703_ VPWR VGND sg13g2_nor3_2
XFILLER_38_853 VPWR VGND sg13g2_decap_8
X_4025_ _1397_ _1353_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[11\]\[4\]
+ net797 sap_3_inst.reg_file_inst.array_serializer_inst.data\[7\]\[4\] VPWR VGND sg13g2_a22oi_1
Xheichips25_sap3_33 VPWR VGND uo_out[6] sg13g2_tielo
XFILLER_40_506 VPWR VGND sg13g2_decap_8
XFILLER_25_569 VPWR VGND sg13g2_decap_8
XFILLER_21_720 VPWR VGND sg13g2_decap_8
X_3809_ _0118_ _1120_ _1227_ net657 _1532_ VPWR VGND sg13g2_a22oi_1
XFILLER_21_797 VPWR VGND sg13g2_decap_8
XFILLER_5_919 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_29_831 VPWR VGND sg13g2_decap_8
XFILLER_44_834 VPWR VGND sg13g2_decap_8
XFILLER_16_569 VPWR VGND sg13g2_decap_8
XFILLER_24_591 VPWR VGND sg13g2_decap_8
XFILLER_8_724 VPWR VGND sg13g2_decap_8
XFILLER_12_786 VPWR VGND sg13g2_decap_8
XFILLER_4_963 VPWR VGND sg13g2_decap_8
XFILLER_3_462 VPWR VGND sg13g2_decap_8
XFILLER_39_606 VPWR VGND sg13g2_decap_8
X_2140_ net760 net757 _1557_ VPWR VGND sg13g2_and2_1
X_2071_ VPWR _1489_ u_ser.state\[1\] VGND sg13g2_inv_1
XFILLER_47_683 VPWR VGND sg13g2_decap_8
XFILLER_35_834 VPWR VGND sg13g2_decap_8
X_2973_ net782 sap_3_inst.alu_inst.tmp\[4\] _0473_ VPWR VGND sg13g2_and2_1
X_3525_ net573 _0990_ _0991_ VPWR VGND sg13g2_and2_1
X_3456_ VGND VPWR net659 _0925_ _0924_ _0923_ sg13g2_a21oi_2
X_2407_ net727 net716 _1823_ _1824_ VPWR VGND sg13g2_nor3_1
X_3387_ _0858_ _0719_ _0731_ VPWR VGND sg13g2_nand2_1
X_2338_ VPWR VGND net752 _1606_ _1754_ _1608_ _1755_ _1614_ sg13g2_a221oi_1
XFILLER_29_105 VPWR VGND sg13g2_fill_2
X_2269_ _1679_ net738 _1684_ _1686_ VPWR VGND sg13g2_a21o_1
XFILLER_38_650 VPWR VGND sg13g2_decap_8
X_4008_ _1381_ VPWR _1382_ VGND _1377_ _1380_ sg13g2_o21ai_1
XFILLER_26_845 VPWR VGND sg13g2_decap_8
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_859 VPWR VGND sg13g2_decap_8
XFILLER_21_594 VPWR VGND sg13g2_decap_8
XFILLER_5_716 VPWR VGND sg13g2_decap_8
XFILLER_0_410 VPWR VGND sg13g2_fill_2
XFILLER_1_933 VPWR VGND sg13g2_decap_8
XFILLER_49_937 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_48_458 VPWR VGND sg13g2_decap_8
XFILLER_29_73 VPWR VGND sg13g2_fill_1
XFILLER_21_1021 VPWR VGND sg13g2_decap_8
XFILLER_44_631 VPWR VGND sg13g2_decap_8
XFILLER_17_856 VPWR VGND sg13g2_decap_8
XFILLER_32_826 VPWR VGND sg13g2_decap_8
XFILLER_40_870 VPWR VGND sg13g2_decap_8
XFILLER_8_521 VPWR VGND sg13g2_decap_8
XFILLER_12_583 VPWR VGND sg13g2_decap_8
XFILLER_8_598 VPWR VGND sg13g2_decap_8
X_3310_ _0781_ net683 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[6\]
+ net686 sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_4_760 VPWR VGND sg13g2_decap_8
X_4290_ net809 VGND VPWR _0147_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[10\]\[1\]
+ clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
X_3241_ _0667_ net689 _0712_ VPWR VGND sg13g2_nor2_1
X_3172_ net750 net728 _1761_ _0643_ VPWR VGND sg13g2_nor3_1
X_2123_ VPWR _1541_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[9\]\[6\]
+ VGND sg13g2_inv_1
XFILLER_27_609 VPWR VGND sg13g2_decap_8
XFILLER_47_480 VPWR VGND sg13g2_decap_8
XFILLER_35_631 VPWR VGND sg13g2_decap_8
XFILLER_22_314 VPWR VGND sg13g2_fill_1
XFILLER_23_837 VPWR VGND sg13g2_decap_8
XFILLER_34_196 VPWR VGND sg13g2_fill_2
X_2956_ VGND VPWR net787 sap_3_inst.alu_inst.tmp\[2\] _0457_ _0415_ sg13g2_a21oi_1
X_2887_ VPWR VGND _0389_ net703 _0387_ net786 _0390_ net691 sg13g2_a221oi_1
XFILLER_2_708 VPWR VGND sg13g2_decap_8
X_3508_ _0975_ net588 _0974_ VPWR VGND sg13g2_nand2_1
X_3439_ _0908_ net681 sap_3_inst.reg_file_inst.array_serializer_inst.data\[6\]\[2\]
+ net684 sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_970 VPWR VGND sg13g2_decap_8
XFILLER_45_428 VPWR VGND sg13g2_decap_8
XFILLER_17_119 VPWR VGND sg13g2_fill_1
XFILLER_26_642 VPWR VGND sg13g2_decap_8
XFILLER_41_656 VPWR VGND sg13g2_decap_8
XFILLER_40_155 VPWR VGND sg13g2_fill_1
XFILLER_40_199 VPWR VGND sg13g2_fill_2
XFILLER_5_513 VPWR VGND sg13g2_decap_8
Xoutput30 net30 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_730 VPWR VGND sg13g2_decap_8
XFILLER_49_734 VPWR VGND sg13g2_decap_8
XFILLER_37_929 VPWR VGND sg13g2_decap_8
XFILLER_17_653 VPWR VGND sg13g2_decap_8
XFILLER_45_995 VPWR VGND sg13g2_decap_8
XFILLER_16_174 VPWR VGND sg13g2_fill_2
XFILLER_32_623 VPWR VGND sg13g2_decap_8
XFILLER_31_133 VPWR VGND sg13g2_fill_1
X_3790_ _1160_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[5\]\[4\] net581
+ _0110_ VPWR VGND sg13g2_mux2_1
X_2810_ net59 sap_3_inst.out\[3\] net799 _0020_ VPWR VGND sg13g2_mux2_1
XFILLER_9_830 VPWR VGND sg13g2_decap_8
X_2741_ net31 _0269_ _1916_ _0270_ VPWR VGND sg13g2_mux2_1
X_2672_ _0206_ _1900_ net785 _1884_ net4 VPWR VGND sg13g2_a22oi_1
X_4342_ mem_mar_we net26 VPWR VGND sg13g2_buf_1
XFILLER_28_1016 VPWR VGND sg13g2_decap_8
X_4273_ net827 VGND VPWR _0130_ sap_3_inst.reg_file_inst.array_serializer_inst.data\[8\]\[0\]
+ clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs sg13g2_dfrbpq_2
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
X_3224_ VGND VPWR net734 _1735_ _0695_ _1815_ sg13g2_a21oi_1
.ends

