module heichips25_sap3 (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire \sap_3_inst.alu_inst.clk_regs ;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire clk_div_out;
 wire mem_mar_we;
 wire mem_ram_we;
 wire regFile_serial;
 wire regFile_serial_start;
 wire \sap_3_inst.alu_flags[0] ;
 wire \sap_3_inst.alu_flags[1] ;
 wire \sap_3_inst.alu_flags[2] ;
 wire \sap_3_inst.alu_flags[3] ;
 wire \sap_3_inst.alu_flags[4] ;
 wire \sap_3_inst.alu_flags[5] ;
 wire \sap_3_inst.alu_flags[6] ;
 wire \sap_3_inst.alu_flags[7] ;
 wire \sap_3_inst.alu_inst.acc[0] ;
 wire \sap_3_inst.alu_inst.acc[1] ;
 wire \sap_3_inst.alu_inst.acc[2] ;
 wire \sap_3_inst.alu_inst.acc[3] ;
 wire \sap_3_inst.alu_inst.acc[4] ;
 wire \sap_3_inst.alu_inst.acc[5] ;
 wire \sap_3_inst.alu_inst.acc[6] ;
 wire \sap_3_inst.alu_inst.acc[7] ;
 wire \sap_3_inst.alu_inst.act[0] ;
 wire \sap_3_inst.alu_inst.act[1] ;
 wire \sap_3_inst.alu_inst.act[2] ;
 wire \sap_3_inst.alu_inst.act[3] ;
 wire \sap_3_inst.alu_inst.act[4] ;
 wire \sap_3_inst.alu_inst.act[5] ;
 wire \sap_3_inst.alu_inst.act[6] ;
 wire \sap_3_inst.alu_inst.act[7] ;
 wire \sap_3_inst.alu_inst.carry ;
 wire \sap_3_inst.alu_inst.clk ;
 wire \sap_3_inst.alu_inst.tmp[0] ;
 wire \sap_3_inst.alu_inst.tmp[1] ;
 wire \sap_3_inst.alu_inst.tmp[2] ;
 wire \sap_3_inst.alu_inst.tmp[3] ;
 wire \sap_3_inst.alu_inst.tmp[4] ;
 wire \sap_3_inst.alu_inst.tmp[5] ;
 wire \sap_3_inst.alu_inst.tmp[6] ;
 wire \sap_3_inst.alu_inst.tmp[7] ;
 wire \sap_3_inst.controller_inst.opcode[0] ;
 wire \sap_3_inst.controller_inst.opcode[1] ;
 wire \sap_3_inst.controller_inst.opcode[2] ;
 wire \sap_3_inst.controller_inst.opcode[3] ;
 wire \sap_3_inst.controller_inst.opcode[4] ;
 wire \sap_3_inst.controller_inst.opcode[5] ;
 wire \sap_3_inst.controller_inst.opcode[6] ;
 wire \sap_3_inst.controller_inst.opcode[7] ;
 wire \sap_3_inst.controller_inst.stage[0] ;
 wire \sap_3_inst.controller_inst.stage[1] ;
 wire \sap_3_inst.controller_inst.stage[2] ;
 wire \sap_3_inst.controller_inst.stage[3] ;
 wire \sap_3_inst.out[0] ;
 wire \sap_3_inst.out[1] ;
 wire \sap_3_inst.out[2] ;
 wire \sap_3_inst.out[3] ;
 wire \sap_3_inst.out[4] ;
 wire \sap_3_inst.out[5] ;
 wire \sap_3_inst.out[6] ;
 wire \sap_3_inst.out[7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[0][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[0][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[0][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[0][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[0][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[0][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[0][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[0][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[3] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[4] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[5] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[6] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[7] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.state[0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.state[1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ;
 wire \sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ;
 wire sap_3_outputReg_serial;
 wire sap_3_outputReg_start_sync;
 wire \u_ser.bit_pos[0] ;
 wire \u_ser.bit_pos[1] ;
 wire \u_ser.bit_pos[2] ;
 wire \u_ser.shadow_reg[0] ;
 wire \u_ser.shadow_reg[1] ;
 wire \u_ser.shadow_reg[2] ;
 wire \u_ser.shadow_reg[3] ;
 wire \u_ser.shadow_reg[4] ;
 wire \u_ser.shadow_reg[5] ;
 wire \u_ser.shadow_reg[6] ;
 wire \u_ser.shadow_reg[7] ;
 wire \u_ser.state[0] ;
 wire \u_ser.state[1] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net34;
 wire net35;
 wire net36;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net31;
 wire net32;
 wire net33;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_0_clk_div_out;
 wire clknet_1_0__leaf_clk_div_out;
 wire clknet_1_1__leaf_clk_div_out;
 wire \clknet_leaf_0_sap_3_inst.alu_inst.clk ;
 wire \clknet_leaf_1_sap_3_inst.alu_inst.clk ;
 wire \clknet_leaf_2_sap_3_inst.alu_inst.clk ;
 wire \clknet_0_sap_3_inst.alu_inst.clk ;
 wire \clknet_1_0__leaf_sap_3_inst.alu_inst.clk ;
 wire \clknet_1_1__leaf_sap_3_inst.alu_inst.clk ;
 wire \clknet_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_0_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_1_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_2_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_3_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_4_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_5_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_6_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_7_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_8_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_9_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_10_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_11_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_12_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_13_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_14_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_4_15_0_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire \clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs ;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;

 sg13g2_inv_2 _2069_ (.Y(_1487_),
    .A(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2070_ (.VDD(VPWR),
    .Y(_1488_),
    .A(\u_ser.state[0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2071_ (.VDD(VPWR),
    .Y(_1489_),
    .A(\u_ser.state[1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2072_ (.VDD(VPWR),
    .Y(_1490_),
    .A(\u_ser.bit_pos[2] ),
    .VSS(VGND));
 sg13g2_inv_2 _2073_ (.Y(_1491_),
    .A(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2074_ (.VDD(VPWR),
    .Y(_1492_),
    .A(net767),
    .VSS(VGND));
 sg13g2_inv_4 _2075_ (.A(net764),
    .Y(_1493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2076_ (.Y(_1494_),
    .A(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2077_ (.VDD(VPWR),
    .Y(_1495_),
    .A(net758),
    .VSS(VGND));
 sg13g2_inv_1 _2078_ (.VDD(VPWR),
    .Y(_1496_),
    .A(net756),
    .VSS(VGND));
 sg13g2_inv_1 _2079_ (.VDD(VPWR),
    .Y(_1497_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2080_ (.VDD(VPWR),
    .Y(_1498_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2081_ (.VDD(VPWR),
    .Y(_1499_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2082_ (.VDD(VPWR),
    .Y(_1500_),
    .A(net788),
    .VSS(VGND));
 sg13g2_inv_2 _2083_ (.Y(_1501_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2084_ (.VDD(VPWR),
    .Y(_1502_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2085_ (.VDD(VPWR),
    .Y(_1503_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2086_ (.VDD(VPWR),
    .Y(_1504_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2087_ (.VDD(VPWR),
    .Y(_1505_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2088_ (.VDD(VPWR),
    .Y(_1506_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2089_ (.VDD(VPWR),
    .Y(_1507_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2090_ (.VDD(VPWR),
    .Y(_1508_),
    .A(net793),
    .VSS(VGND));
 sg13g2_inv_4 _2091_ (.A(net781),
    .Y(_1509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2092_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][1] ),
    .Y(_1510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2093_ (.VDD(VPWR),
    .Y(_1511_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2094_ (.VDD(VPWR),
    .Y(_1512_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2095_ (.VDD(VPWR),
    .Y(_1513_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2096_ (.VDD(VPWR),
    .Y(_1514_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2097_ (.VDD(VPWR),
    .Y(_1515_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2098_ (.VDD(VPWR),
    .Y(_1516_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2099_ (.VDD(VPWR),
    .Y(_1517_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2100_ (.VDD(VPWR),
    .Y(_1518_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2101_ (.VDD(VPWR),
    .Y(_1519_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2102_ (.VDD(VPWR),
    .Y(_1520_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2103_ (.VDD(VPWR),
    .Y(_1521_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2104_ (.VDD(VPWR),
    .Y(_1522_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2105_ (.VDD(VPWR),
    .Y(_1523_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2106_ (.VDD(VPWR),
    .Y(_1524_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2107_ (.VDD(VPWR),
    .Y(_1525_),
    .A(\sap_3_inst.alu_inst.act[0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2108_ (.VDD(VPWR),
    .Y(_1526_),
    .A(\sap_3_inst.alu_inst.act[7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2109_ (.VDD(VPWR),
    .Y(_1527_),
    .A(\sap_3_inst.alu_inst.tmp[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2110_ (.VDD(VPWR),
    .Y(_1528_),
    .A(\sap_3_inst.alu_inst.tmp[6] ),
    .VSS(VGND));
 sg13g2_inv_2 _2111_ (.Y(_1529_),
    .A(\sap_3_inst.alu_inst.tmp[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2112_ (.VDD(VPWR),
    .Y(_1530_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2113_ (.VDD(VPWR),
    .Y(_1531_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2114_ (.VDD(VPWR),
    .Y(_1532_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2115_ (.VDD(VPWR),
    .Y(_1533_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2116_ (.VDD(VPWR),
    .Y(_1534_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2117_ (.VDD(VPWR),
    .Y(_1535_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .VSS(VGND));
 sg13g2_inv_1 _2118_ (.VDD(VPWR),
    .Y(_1536_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2119_ (.VDD(VPWR),
    .Y(_1537_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2120_ (.VDD(VPWR),
    .Y(_1538_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .VSS(VGND));
 sg13g2_inv_2 _2121_ (.Y(_1539_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2122_ (.VDD(VPWR),
    .Y(_1540_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2123_ (.VDD(VPWR),
    .Y(_1541_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2124_ (.VDD(VPWR),
    .Y(_1542_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2125_ (.VDD(VPWR),
    .Y(_1543_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2126_ (.VDD(VPWR),
    .Y(_1544_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ),
    .VSS(VGND));
 sg13g2_inv_2 _2127_ (.Y(_1545_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2128_ (.VDD(VPWR),
    .Y(_1546_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2129_ (.VDD(VPWR),
    .Y(_1547_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2130_ (.VDD(VPWR),
    .Y(_1548_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2131_ (.VDD(VPWR),
    .Y(_1549_),
    .A(net50),
    .VSS(VGND));
 sg13g2_inv_1 _2132_ (.VDD(VPWR),
    .Y(_1550_),
    .A(net52),
    .VSS(VGND));
 sg13g2_inv_1 _4145__3 (.VDD(VPWR),
    .Y(net37),
    .A(\clknet_leaf_1_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_nor2_2 _2134_ (.A(net745),
    .B(net744),
    .Y(_1551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2135_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1552_),
    .B(net744),
    .A(net745));
 sg13g2_nor2_2 _2136_ (.A(net747),
    .B(net746),
    .Y(_1553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2137_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1554_),
    .B(net746),
    .A(net747));
 sg13g2_nand2b_2 _2138_ (.Y(_1555_),
    .B(net743),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\sap_3_inst.controller_inst.stage[1] ));
 sg13g2_nor2_2 _2139_ (.A(_1552_),
    .B(_1554_),
    .Y(_1556_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2140_ (.A(net760),
    .B(net757),
    .X(_1557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2141_ (.Y(_1558_),
    .A(net759),
    .B(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2142_ (.A(net763),
    .B(net752),
    .Y(_1559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2143_ (.B(net760),
    .C(net757),
    .Y(_1560_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net762));
 sg13g2_nor2b_2 _2144_ (.A(net770),
    .B_N(net767),
    .Y(_1561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2145_ (.Y(_1562_),
    .B(net768),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net770));
 sg13g2_nand3b_1 _2146_ (.B(net765),
    .C(net768),
    .Y(_1563_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net771));
 sg13g2_nor2_1 _2147_ (.A(net753),
    .B(_1496_),
    .Y(_1564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2148_ (.Y(_1565_),
    .B(net756),
    .A_N(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2149_ (.A(net751),
    .B(net750),
    .Y(_1566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2150_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1567_),
    .B(net750),
    .A(net751));
 sg13g2_nor2_1 _2151_ (.A(_1560_),
    .B(net750),
    .Y(_1568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2152_ (.Y(_1569_),
    .A(_1559_),
    .B(_1564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2153_ (.A(net753),
    .B(net755),
    .Y(_1570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2154_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1571_),
    .B(net755),
    .A(net753));
 sg13g2_nor3_1 _2155_ (.A(net766),
    .B(net754),
    .C(net755),
    .Y(_1572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2156_ (.A(net766),
    .B(net754),
    .C(net755),
    .X(_1573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2157_ (.A(net763),
    .B(net765),
    .C(net753),
    .Y(_1574_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net755));
 sg13g2_or2_1 _2158_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1575_),
    .B(net757),
    .A(net760));
 sg13g2_or2_1 _2159_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1576_),
    .B(net770),
    .A(net767));
 sg13g2_nor2_1 _2160_ (.A(_1575_),
    .B(_1576_),
    .Y(_1577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2161_ (.Y(_1578_),
    .B1(_1574_),
    .B2(_1577_),
    .A2(net742),
    .A1(_1559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2162_ (.VDD(VPWR),
    .Y(_1579_),
    .A(_1578_),
    .VSS(VGND));
 sg13g2_and2_1 _2163_ (.A(net747),
    .B(net746),
    .X(_1580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2164_ (.Y(_1581_),
    .A(net747),
    .B(\sap_3_inst.controller_inst.stage[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2165_ (.A(_1552_),
    .B(_1581_),
    .Y(_1582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2166_ (.Y(_1583_),
    .A(net743),
    .B(_1580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2167_ (.A(net746),
    .B_N(net747),
    .Y(_1584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2168_ (.A(_1491_),
    .B(_1555_),
    .Y(_1585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2169_ (.A(net747),
    .B_N(net746),
    .Y(_1586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2170_ (.Y(_1587_),
    .A(net747),
    .B(net746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2171_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net743),
    .C1(net718),
    .B1(net737),
    .A1(net741),
    .Y(_1588_),
    .A2(net727));
 sg13g2_nand2_1 _2172_ (.Y(_1589_),
    .A(_1578_),
    .B(_1588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2173_ (.Y(_1590_),
    .A(net739),
    .B(net727),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2174_ (.VDD(VPWR),
    .Y(_1591_),
    .A(_1590_),
    .VSS(VGND));
 sg13g2_nor4_2 _2175_ (.A(_1494_),
    .B(_1560_),
    .C(_1571_),
    .Y(_1592_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1576_));
 sg13g2_and2_1 _2176_ (.A(net730),
    .B(_1592_),
    .X(_1593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2177_ (.A(net739),
    .B(_1593_),
    .Y(_1594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2178_ (.A(net755),
    .B_N(net753),
    .Y(_1595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2179_ (.Y(_1596_),
    .A(net753),
    .B(_1496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2180_ (.B(_1561_),
    .C(net731),
    .A(net765),
    .Y(_1597_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1595_));
 sg13g2_nor2_1 _2181_ (.A(net751),
    .B(_1596_),
    .Y(_1598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2182_ (.Y(_1599_),
    .A(_1594_),
    .B(_1597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2183_ (.B(net765),
    .C(_1570_),
    .A(_1492_),
    .Y(_1600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2184_ (.A(_1598_),
    .B_N(_1600_),
    .Y(_1601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2185_ (.B1(_1600_),
    .VDD(VPWR),
    .Y(_1602_),
    .VSS(VGND),
    .A1(net751),
    .A2(_1596_));
 sg13g2_and3_2 _2186_ (.X(_1603_),
    .A(net765),
    .B(net753),
    .C(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2187_ (.B(net753),
    .C(net755),
    .A(net766),
    .Y(_1604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2188_ (.Y(_1605_),
    .A(_1561_),
    .B(_1603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2189_ (.A(net728),
    .B(_1605_),
    .Y(_1606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2190_ (.Y(_1607_),
    .B(_1570_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net751));
 sg13g2_nor2_1 _2191_ (.A(_1560_),
    .B(_1607_),
    .Y(_1608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2192_ (.A(_1560_),
    .B(net751),
    .C(_1571_),
    .X(_1609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2193_ (.A(net744),
    .B_N(net745),
    .Y(_1610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2194_ (.Y(_1611_),
    .B(net745),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net744));
 sg13g2_and2_1 _2195_ (.A(net738),
    .B(net736),
    .X(_1612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2196_ (.Y(_1613_),
    .A(net738),
    .B(_1610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2197_ (.Y(_1614_),
    .A(net729),
    .B(net725),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2198_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1608_),
    .A2(_1614_),
    .Y(_1615_),
    .B1(_1606_));
 sg13g2_nand2_2 _2199_ (.Y(_1616_),
    .A(net767),
    .B(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2200_ (.B(net771),
    .C(net765),
    .A(net767),
    .Y(_1617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2201_ (.A(_1571_),
    .B(_1617_),
    .Y(_1618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2202_ (.B(_1605_),
    .C(_1609_),
    .A(_1596_),
    .Y(_1619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2203_ (.A(_1618_),
    .B(_1619_),
    .Y(_1620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2204_ (.VDD(VPWR),
    .Y(_1621_),
    .A(_1620_),
    .VSS(VGND));
 sg13g2_a21o_1 _2205_ (.A2(_1621_),
    .A1(_1615_),
    .B1(_1602_),
    .X(_1622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2206_ (.A(net767),
    .B_N(net770),
    .Y(_1623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2207_ (.Y(_1624_),
    .B(net770),
    .A_N(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2208_ (.B(net754),
    .C(net756),
    .Y(_1625_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net766));
 sg13g2_nor2_1 _2209_ (.A(net762),
    .B(_1625_),
    .Y(_1626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2210_ (.A(net762),
    .B(_1624_),
    .C(_1625_),
    .Y(_1627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2211_ (.B(_1493_),
    .C(_1623_),
    .Y(_1628_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net749));
 sg13g2_and2_1 _2212_ (.A(net737),
    .B(_1610_),
    .X(_1629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2213_ (.Y(_1630_),
    .A(net737),
    .B(net736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2214_ (.Y(_1631_),
    .B1(net737),
    .B2(net736),
    .A2(_1580_),
    .A1(net743),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2215_ (.A(_1628_),
    .B(net724),
    .Y(_1632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2216_ (.A(_1587_),
    .B(net736),
    .X(_1633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2217_ (.Y(_1634_),
    .A(_1587_),
    .B(net736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2218_ (.A(_1604_),
    .B(_1624_),
    .Y(_1635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2219_ (.Y(_1636_),
    .A(_1603_),
    .B(_1623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2220_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1632_),
    .Y(_1637_),
    .A2(_1635_),
    .A1(_1633_));
 sg13g2_nor2_1 _2221_ (.A(net770),
    .B(net749),
    .Y(_1638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2222_ (.A(net762),
    .B(_1575_),
    .C(_1616_),
    .Y(_1639_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1625_));
 sg13g2_or4_1 _2223_ (.A(net763),
    .B(_1575_),
    .C(_1616_),
    .D(net749),
    .X(_1640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2224_ (.B(net770),
    .C(net762),
    .Y(_1641_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net767));
 sg13g2_nor2_1 _2225_ (.A(_1575_),
    .B(_1641_),
    .Y(_1642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2226_ (.A(_1575_),
    .B(net749),
    .C(_1641_),
    .Y(_1643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2227_ (.A(_1575_),
    .B(net749),
    .C(_1641_),
    .X(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2228_ (.A(_1574_),
    .B(_1623_),
    .X(_1645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2229_ (.Y(_1646_),
    .A(_1574_),
    .B(_1623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2230_ (.A(_1643_),
    .B(_1645_),
    .Y(_1647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _2231_ (.A(_1638_),
    .B(_1639_),
    .C(_1643_),
    .D(_1645_),
    .X(_1648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2232_ (.A(_1576_),
    .B(_1604_),
    .Y(_1649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2233_ (.Y(_1650_),
    .B(_1603_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1576_));
 sg13g2_nor3_2 _2234_ (.A(_1575_),
    .B(_1604_),
    .C(_1641_),
    .Y(_1651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2235_ (.A(_1575_),
    .B(_1604_),
    .C(_1641_),
    .X(_1652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2236_ (.A(_1649_),
    .B(_1651_),
    .Y(_1653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2237_ (.Y(_1654_),
    .A(_1650_),
    .B(net735),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2238_ (.A(net761),
    .B_N(net757),
    .Y(_1655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2239_ (.Y(_1656_),
    .B(net758),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net759));
 sg13g2_nor2_2 _2240_ (.A(_1562_),
    .B(_1573_),
    .Y(_1657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2241_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1656_),
    .A2(_1657_),
    .Y(_1658_),
    .B1(_1654_));
 sg13g2_nor3_2 _2242_ (.A(_1562_),
    .B(_1573_),
    .C(_1656_),
    .Y(_1659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2243_ (.B(_1572_),
    .C(_1655_),
    .A(_1561_),
    .Y(_1660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2244_ (.A(_1573_),
    .B(_1641_),
    .Y(_1661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2245_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1662_),
    .B(_1641_),
    .A(_1573_));
 sg13g2_nand2_1 _2246_ (.Y(_1663_),
    .A(_1607_),
    .B(net733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2247_ (.A(_1648_),
    .B(_1654_),
    .C(_1657_),
    .D(_1663_),
    .Y(_1664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2248_ (.Y(_1665_),
    .A(_1637_),
    .B(net714),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2249_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1666_),
    .B(net749),
    .A(_1576_));
 sg13g2_nor2b_2 _2250_ (.A(\sap_3_inst.controller_inst.opcode[5] ),
    .B_N(net760),
    .Y(_1667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _2251_ (.S0(net757),
    .A0(\sap_3_inst.alu_flags[0] ),
    .A1(\sap_3_inst.alu_flags[2] ),
    .A2(net748),
    .A3(\sap_3_inst.alu_flags[3] ),
    .S1(net760),
    .X(_1668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2252_ (.Y(_1669_),
    .A(net762),
    .B(_1668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2253_ (.Y(_1670_),
    .A(net730),
    .B(_1669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2254_ (.A(\sap_3_inst.controller_inst.stage[2] ),
    .B_N(net744),
    .Y(_1671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2255_ (.A(net738),
    .B(net732),
    .X(_1672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2256_ (.Y(_1673_),
    .A(_1584_),
    .B(net732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2257_ (.A(_1629_),
    .B(_1672_),
    .Y(_1674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2258_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1670_),
    .A2(_1674_),
    .Y(_1675_),
    .B1(_1666_));
 sg13g2_nor2_1 _2259_ (.A(net731),
    .B(_1672_),
    .Y(_1676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2260_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net724),
    .A2(_1673_),
    .Y(_1677_),
    .B1(_1644_));
 sg13g2_or3_1 _2261_ (.A(net714),
    .B(_1675_),
    .C(_1677_),
    .X(_1678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2262_ (.A(net745),
    .B(net744),
    .X(_1679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2263_ (.Y(_1680_),
    .A(\sap_3_inst.controller_inst.stage[2] ),
    .B(net744),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2264_ (.Y(_1681_),
    .A(net745),
    .B(_1580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2265_ (.Y(_1682_),
    .A(_1580_),
    .B(_1679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2266_ (.B(\sap_3_inst.controller_inst.stage[3] ),
    .C(net746),
    .Y(_1683_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net745));
 sg13g2_nor2_2 _2267_ (.A(\sap_3_inst.controller_inst.stage[0] ),
    .B(_1683_),
    .Y(_1684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2268_ (.Y(_1685_),
    .B1(_1679_),
    .B2(net738),
    .A2(net732),
    .A1(net737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2269_ (.A2(_1679_),
    .A1(net738),
    .B1(_1684_),
    .X(_1686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2270_ (.Y(_1687_),
    .A(_1630_),
    .B(_1670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2271_ (.Y(_1688_),
    .A(_1682_),
    .B(_1685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2272_ (.B1(_1649_),
    .VDD(VPWR),
    .Y(_1689_),
    .VSS(VGND),
    .A1(_1687_),
    .A2(_1688_));
 sg13g2_nor2_1 _2273_ (.A(_1562_),
    .B(net749),
    .Y(_1690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2274_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1691_),
    .B(net749),
    .A(_1562_));
 sg13g2_and2_1 _2275_ (.A(_1553_),
    .B(net732),
    .X(_1692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2276_ (.Y(_1693_),
    .A(_1553_),
    .B(_1671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2277_ (.A(_1629_),
    .B(_1692_),
    .Y(_1694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2278_ (.A2(_1694_),
    .A1(_1670_),
    .B1(_1691_),
    .X(_1695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2279_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net724),
    .A2(_1693_),
    .Y(_1696_),
    .B1(_1646_));
 sg13g2_nor2_2 _2280_ (.A(net726),
    .B(_1607_),
    .Y(_1697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2281_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net726),
    .A2(_1682_),
    .Y(_1698_),
    .B1(net735));
 sg13g2_nor3_2 _2282_ (.A(_1558_),
    .B(_1562_),
    .C(_1573_),
    .Y(_1699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2283_ (.B(_1561_),
    .C(_1572_),
    .A(_1557_),
    .Y(_1700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2284_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net724),
    .A2(_1673_),
    .Y(_1701_),
    .B1(_1700_));
 sg13g2_a21oi_1 _2285_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1630_),
    .A2(_1685_),
    .Y(_1702_),
    .B1(net735));
 sg13g2_nor3_2 _2286_ (.A(net758),
    .B(_1562_),
    .C(_1573_),
    .Y(_1703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2287_ (.A(_1612_),
    .B(_1703_),
    .X(_1704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2288_ (.A(_1491_),
    .B(_1683_),
    .Y(_1705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2289_ (.Y(_1706_),
    .A(_1580_),
    .B(net732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2290_ (.A(net733),
    .B(_1706_),
    .Y(_1707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2291_ (.A(_1704_),
    .B(_1707_),
    .Y(_1708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2292_ (.Y(_1709_),
    .B1(_1679_),
    .B2(_1553_),
    .A2(net732),
    .A1(net738),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2293_ (.A(_1660_),
    .B(_1709_),
    .Y(_1710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2294_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net724),
    .A2(_1709_),
    .Y(_1711_),
    .B1(_1660_));
 sg13g2_a22oi_1 _2295_ (.Y(_1712_),
    .B1(_1693_),
    .B2(_1631_),
    .A2(_1646_),
    .A1(_1640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2296_ (.A(_1698_),
    .B(_1702_),
    .C(_1711_),
    .D(_1712_),
    .Y(_1713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2297_ (.A(_1697_),
    .B(_1701_),
    .C(_1704_),
    .D(_1707_),
    .Y(_1714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2298_ (.B(_1695_),
    .C(_1713_),
    .A(_1689_),
    .Y(_1715_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1714_));
 sg13g2_o21ai_1 _2299_ (.B1(_1665_),
    .VDD(VPWR),
    .Y(_1716_),
    .VSS(VGND),
    .A1(_1678_),
    .A2(_1715_));
 sg13g2_a21oi_1 _2300_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1620_),
    .A2(_1716_),
    .Y(_1717_),
    .B1(_1622_));
 sg13g2_o21ai_1 _2301_ (.B1(_1590_),
    .VDD(VPWR),
    .Y(_1718_),
    .VSS(VGND),
    .A1(_1599_),
    .A2(_1717_));
 sg13g2_a21oi_1 _2302_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net740),
    .A2(_1718_),
    .Y(_1719_),
    .B1(_1589_));
 sg13g2_nor2_2 _2303_ (.A(_1556_),
    .B(_1719_),
    .Y(_1720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2304_ (.VDD(VPWR),
    .Y(_1721_),
    .A(_1720_),
    .VSS(VGND));
 sg13g2_nor2_1 _2305_ (.A(_1554_),
    .B(_1611_),
    .Y(_1722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2306_ (.Y(_1723_),
    .A(_1553_),
    .B(net736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2307_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1617_),
    .A2(net722),
    .Y(_1724_),
    .B1(_1590_));
 sg13g2_a21oi_1 _2308_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net758),
    .A2(_1657_),
    .Y(_1725_),
    .B1(_1651_));
 sg13g2_nor4_1 _2309_ (.A(_1643_),
    .B(_1651_),
    .C(_1657_),
    .D(_1661_),
    .Y(_1726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2310_ (.Y(_1727_),
    .B(_1726_),
    .A_N(_1694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2311_ (.VDD(VPWR),
    .Y(_1728_),
    .A(_1727_),
    .VSS(VGND));
 sg13g2_o21ai_1 _2312_ (.B1(net722),
    .VDD(VPWR),
    .Y(_1729_),
    .VSS(VGND),
    .A1(net734),
    .A2(_1703_));
 sg13g2_nor3_2 _2313_ (.A(net764),
    .B(_1660_),
    .C(_1685_),
    .Y(_1730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2314_ (.A(_1581_),
    .B(_1611_),
    .Y(_1731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2315_ (.VDD(VPWR),
    .Y(_1732_),
    .A(_1731_),
    .VSS(VGND));
 sg13g2_nand2_1 _2316_ (.Y(_1733_),
    .A(_1587_),
    .B(net732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2317_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1732_),
    .A2(_1733_),
    .Y(_1734_),
    .B1(net733));
 sg13g2_nand2_1 _2318_ (.Y(_1735_),
    .A(_1630_),
    .B(_1683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2319_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1554_),
    .A2(_1679_),
    .Y(_1736_),
    .B1(_1735_));
 sg13g2_nor2_1 _2320_ (.A(net735),
    .B(_1736_),
    .Y(_1737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2321_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1629_),
    .A2(_1659_),
    .Y(_1738_),
    .B1(net730));
 sg13g2_nor4_1 _2322_ (.A(_1677_),
    .B(_1701_),
    .C(_1734_),
    .D(_1737_),
    .Y(_1739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2323_ (.A(_1704_),
    .B(_1710_),
    .C(_1728_),
    .D(_1730_),
    .Y(_1740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2324_ (.B(_1738_),
    .C(_1739_),
    .A(_1729_),
    .Y(_1741_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1740_));
 sg13g2_nand2_1 _2325_ (.Y(_1742_),
    .A(_1640_),
    .B(_1726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2326_ (.B1(_1741_),
    .VDD(VPWR),
    .Y(_1743_),
    .VSS(VGND),
    .A1(_1696_),
    .A2(_1742_));
 sg13g2_nand2b_2 _2327_ (.Y(_1744_),
    .B(net730),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1669_));
 sg13g2_nand2_1 _2328_ (.Y(_1745_),
    .A(_1649_),
    .B(_1744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2329_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net726),
    .A2(_1736_),
    .Y(_1746_),
    .B1(_1745_));
 sg13g2_nand2b_1 _2330_ (.Y(_1747_),
    .B(net735),
    .A_N(_1637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2331_ (.A(_1609_),
    .B(_1630_),
    .Y(_1748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2332_ (.Y(_1749_),
    .A(net731),
    .B(_1617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2333_ (.A(_1596_),
    .B(_1749_),
    .Y(_1750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2334_ (.A(_1602_),
    .B(_1697_),
    .C(_1748_),
    .D(_1750_),
    .Y(_1751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2335_ (.Y(_1752_),
    .B1(net732),
    .B2(_1553_),
    .A2(net736),
    .A1(net738),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2336_ (.Y(_1753_),
    .A(net725),
    .B(_1693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2337_ (.A(_1636_),
    .B(_1642_),
    .C(net720),
    .Y(_1754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2338_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net752),
    .C1(_1606_),
    .B1(_1754_),
    .A1(_1608_),
    .Y(_1755_),
    .A2(_1614_));
 sg13g2_nand4_1 _2339_ (.B(_1747_),
    .C(_1751_),
    .A(_1695_),
    .Y(_1756_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1755_));
 sg13g2_nor3_1 _2340_ (.A(_1675_),
    .B(_1746_),
    .C(_1756_),
    .Y(_1757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2341_ (.B1(net750),
    .VDD(VPWR),
    .Y(_1758_),
    .VSS(VGND),
    .A1(_1573_),
    .A2(_1616_));
 sg13g2_nor2_2 _2342_ (.A(_1592_),
    .B(_1758_),
    .Y(_1759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2343_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1760_),
    .B(_1758_),
    .A(_1592_));
 sg13g2_nor2_1 _2344_ (.A(_1493_),
    .B(net752),
    .Y(_1761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2345_ (.B(net760),
    .C(net757),
    .A(net763),
    .Y(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2346_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net731),
    .A2(_1762_),
    .Y(_1763_),
    .B1(net716));
 sg13g2_a221oi_1 _2347_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1597_),
    .C1(net719),
    .B1(_1763_),
    .A1(_1743_),
    .Y(_1764_),
    .A2(_1757_));
 sg13g2_nor2_1 _2348_ (.A(net750),
    .B(_1749_),
    .Y(_1765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2349_ (.A(net739),
    .B(_1593_),
    .C(_1764_),
    .D(_1765_),
    .Y(_1766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2350_ (.B1(_1567_),
    .VDD(VPWR),
    .Y(_1767_),
    .VSS(VGND),
    .A1(_1724_),
    .A2(_1766_));
 sg13g2_nand4_1 _2351_ (.B(_1588_),
    .C(_1720_),
    .A(_1578_),
    .Y(_1768_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1767_));
 sg13g2_nand2_1 _2352_ (.Y(_1769_),
    .A(net765),
    .B(_1616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2353_ (.A(net727),
    .B(_1769_),
    .Y(_1770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2354_ (.A(_1759_),
    .B(_1770_),
    .Y(_1771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2355_ (.A(_1636_),
    .B(_1656_),
    .C(net720),
    .Y(_1772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2356_ (.A(net729),
    .B(_1662_),
    .Y(_1773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2357_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1595_),
    .C1(net719),
    .B1(_1770_),
    .A1(net730),
    .Y(_1774_),
    .A2(net734));
 sg13g2_a21oi_1 _2358_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net764),
    .A2(net761),
    .Y(_1775_),
    .B1(_1495_));
 sg13g2_nor2_1 _2359_ (.A(_1639_),
    .B(_1690_),
    .Y(_1776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2360_ (.B(_1646_),
    .C(_1691_),
    .A(_1640_),
    .Y(_1777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2361_ (.A(_1653_),
    .B(_1682_),
    .Y(_1778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2362_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1693_),
    .A2(net721),
    .Y(_1779_),
    .B1(_1656_));
 sg13g2_nor3_1 _2363_ (.A(_1705_),
    .B(_1731_),
    .C(_1779_),
    .Y(_1780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2364_ (.A(net733),
    .B(_1780_),
    .Y(_1781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2365_ (.Y(_1782_),
    .A(_1644_),
    .B(_1666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2366_ (.Y(_1783_),
    .B1(_1782_),
    .B2(_1672_),
    .A2(_1777_),
    .A1(_1692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2367_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1672_),
    .A2(_1699_),
    .Y(_1784_),
    .B1(_1710_));
 sg13g2_and3_1 _2368_ (.X(_1785_),
    .A(net730),
    .B(_1602_),
    .C(_1775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2369_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net725),
    .A2(_1630_),
    .Y(_1786_),
    .B1(_1609_));
 sg13g2_nor4_1 _2370_ (.A(_1704_),
    .B(_1730_),
    .C(_1772_),
    .D(_1786_),
    .Y(_1787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2371_ (.B(_1783_),
    .C(_1784_),
    .A(_1774_),
    .Y(_1788_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1787_));
 sg13g2_nor4_1 _2372_ (.A(_1778_),
    .B(_1781_),
    .C(_1785_),
    .D(_1788_),
    .Y(_1789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2373_ (.B1(_1569_),
    .VDD(VPWR),
    .Y(_1790_),
    .VSS(VGND),
    .A1(_1771_),
    .A2(_1789_));
 sg13g2_o21ai_1 _2374_ (.B1(_1591_),
    .VDD(VPWR),
    .Y(_1791_),
    .VSS(VGND),
    .A1(net721),
    .A2(_1769_));
 sg13g2_and4_1 _2375_ (.A(_1555_),
    .B(_1578_),
    .C(_1790_),
    .D(_1791_),
    .X(_1792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2376_ (.VDD(VPWR),
    .Y(_1793_),
    .A(net696),
    .VSS(VGND));
 sg13g2_nor2_1 _2377_ (.A(_1638_),
    .B(_1649_),
    .Y(_1794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2378_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1630_),
    .A2(_1670_),
    .Y(_1795_),
    .B1(_1794_));
 sg13g2_nor2_1 _2379_ (.A(_1653_),
    .B(_1706_),
    .Y(_1796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2380_ (.A(net737),
    .B(_1679_),
    .X(_1797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2381_ (.B1(_1654_),
    .VDD(VPWR),
    .Y(_1798_),
    .VSS(VGND),
    .A1(_1705_),
    .A2(_1797_));
 sg13g2_nor2_1 _2382_ (.A(net724),
    .B(_1725_),
    .Y(_1799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2383_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net733),
    .Y(_1800_),
    .A2(net721),
    .A1(_1693_));
 sg13g2_a22oi_1 _2384_ (.Y(_1801_),
    .B1(_1800_),
    .B2(_1557_),
    .A2(_1686_),
    .A1(_1654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2385_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1640_),
    .A2(_1647_),
    .Y(_1802_),
    .B1(_1631_));
 sg13g2_nand2b_1 _2386_ (.Y(_1803_),
    .B(_1801_),
    .A_N(_1697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2387_ (.A(_1799_),
    .B_N(_1798_),
    .Y(_1804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2388_ (.A(net714),
    .B(_1795_),
    .C(_1802_),
    .D(_1803_),
    .Y(_1805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2389_ (.Y(_1806_),
    .B1(_1804_),
    .B2(_1805_),
    .A2(net714),
    .A1(_1637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2390_ (.A(_1556_),
    .B(_1606_),
    .C(_1806_),
    .X(_1807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2391_ (.VDD(VPWR),
    .Y(_1808_),
    .A(_1807_),
    .VSS(VGND));
 sg13g2_nor2_2 _2392_ (.A(net696),
    .B(_1807_),
    .Y(_1809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2393_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1810_),
    .B(_1807_),
    .A(net696));
 sg13g2_a21oi_1 _2394_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net768),
    .A2(_1765_),
    .Y(_1811_),
    .B1(_1759_));
 sg13g2_nand3_1 _2395_ (.B(_1667_),
    .C(_1753_),
    .A(_1635_),
    .Y(_1812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2396_ (.B(net714),
    .C(_1812_),
    .A(_1637_),
    .Y(_1813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2397_ (.Y(_1814_),
    .B1(net736),
    .B2(_1553_),
    .A2(_1580_),
    .A1(net743),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2398_ (.A(_1814_),
    .B_N(_1703_),
    .Y(_1815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2399_ (.Y(_1816_),
    .B(_1703_),
    .A_N(_1814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2400_ (.B1(net759),
    .VDD(VPWR),
    .Y(_1817_),
    .VSS(VGND),
    .A1(_1800_),
    .A2(_1815_));
 sg13g2_a22oi_1 _2401_ (.Y(_1818_),
    .B1(_1692_),
    .B2(_1777_),
    .A2(_1688_),
    .A1(_1654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2402_ (.B(_1784_),
    .C(_1817_),
    .A(_1708_),
    .Y(_1819_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1818_));
 sg13g2_o21ai_1 _2403_ (.B1(_1813_),
    .VDD(VPWR),
    .Y(_1820_),
    .VSS(VGND),
    .A1(_1678_),
    .A2(_1819_));
 sg13g2_a21oi_1 _2404_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net769),
    .A2(_1750_),
    .Y(_1821_),
    .B1(_1748_));
 sg13g2_and2_1 _2405_ (.A(net759),
    .B(_1762_),
    .X(_1822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2406_ (.Y(_1823_),
    .A(net759),
    .B(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2407_ (.A(net727),
    .B(net716),
    .C(_1823_),
    .Y(_1824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2408_ (.X(_1825_),
    .A(_1820_),
    .B(_1821_),
    .C(_1824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2409_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1820_),
    .A2(_1821_),
    .Y(_1826_),
    .B1(_1602_));
 sg13g2_nor3_1 _2410_ (.A(net719),
    .B(_1825_),
    .C(_1826_),
    .Y(_1827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2411_ (.B1(_1569_),
    .VDD(VPWR),
    .Y(_1828_),
    .VSS(VGND),
    .A1(_1811_),
    .A2(_1827_));
 sg13g2_nand3_1 _2412_ (.B(_1617_),
    .C(net722),
    .A(net769),
    .Y(_1829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2413_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net739),
    .C1(net741),
    .B1(_1829_),
    .A1(net743),
    .Y(_1830_),
    .A2(_1581_));
 sg13g2_nand4_1 _2414_ (.B(_1553_),
    .C(_1610_),
    .A(\sap_3_inst.controller_inst.opcode[0] ),
    .Y(_1831_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1617_));
 sg13g2_nand2_2 _2415_ (.Y(_1832_),
    .A(net739),
    .B(_1831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2416_ (.A(net752),
    .B(_1635_),
    .C(net715),
    .D(_1692_),
    .X(_1833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2417_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net750),
    .A2(_1620_),
    .Y(_1834_),
    .B1(_1749_));
 sg13g2_nand3_1 _2418_ (.B(_1659_),
    .C(_1679_),
    .A(net738),
    .Y(_1835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2419_ (.A(net764),
    .B(_1835_),
    .Y(_1836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2420_ (.Y(_1837_),
    .A(net763),
    .B(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2421_ (.A(net728),
    .B(_1600_),
    .C(_1837_),
    .Y(_1838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2422_ (.B1(_1729_),
    .VDD(VPWR),
    .Y(_1839_),
    .VSS(VGND),
    .A1(net726),
    .A2(net733));
 sg13g2_nor4_1 _2423_ (.A(net713),
    .B(_1833_),
    .C(_1836_),
    .D(_1839_),
    .Y(_1840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2424_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net771),
    .A2(_1834_),
    .Y(_1841_),
    .B1(_1838_));
 sg13g2_nand3_1 _2425_ (.B(_1840_),
    .C(_1841_),
    .A(_1569_),
    .Y(_1842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2426_ (.A(_1832_),
    .B(_1842_),
    .X(_1843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2427_ (.VDD(VPWR),
    .Y(_1844_),
    .A(_1843_),
    .VSS(VGND));
 sg13g2_a221oi_1 _2428_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1842_),
    .C1(_1810_),
    .B1(_1832_),
    .A1(net666),
    .Y(_1845_),
    .A2(net707));
 sg13g2_nand2_1 _2429_ (.Y(_1846_),
    .A(_1545_),
    .B(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2430_ (.A(net667),
    .B(net666),
    .C(net707),
    .D(_1843_),
    .X(_1847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2431_ (.Y(_1848_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2432_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net666),
    .A2(net707),
    .Y(_1849_),
    .B1(_1844_));
 sg13g2_and2_1 _2433_ (.A(net696),
    .B(_1849_),
    .X(_1850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2434_ (.B(net696),
    .C(net626),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .Y(_1851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2435_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1842_),
    .C1(_1793_),
    .B1(_1832_),
    .A1(net666),
    .Y(_1852_),
    .A2(net707));
 sg13g2_and4_1 _2436_ (.A(net667),
    .B(net666),
    .C(net707),
    .D(_1844_),
    .X(_1853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2437_ (.Y(_1854_),
    .B1(net623),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .A2(net624),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2438_ (.B(_1851_),
    .C(_1854_),
    .A(_1848_),
    .Y(_1855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2439_ (.A(_1807_),
    .B(_1828_),
    .C(_1830_),
    .D(_1843_),
    .X(_1856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2440_ (.VDD(VPWR),
    .Y(_1857_),
    .A(net621),
    .VSS(VGND));
 sg13g2_a221oi_1 _2441_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .C1(net631),
    .B1(net621),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .Y(_1858_),
    .A2(net711));
 sg13g2_and4_1 _2442_ (.A(_1807_),
    .B(net666),
    .C(net707),
    .D(_1844_),
    .X(_1859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2443_ (.A(net696),
    .B(net666),
    .C(net707),
    .D(_1844_),
    .X(_1860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2444_ (.Y(_1861_),
    .B1(net616),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .A2(net619),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2445_ (.A(net667),
    .B(net627),
    .X(_1862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2446_ (.B(net667),
    .C(net626),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .Y(_1863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2447_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1842_),
    .C1(_1808_),
    .B1(_1832_),
    .A1(net666),
    .Y(_1864_),
    .A2(net707));
 sg13g2_nand2_1 _2448_ (.Y(_1865_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .B(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2449_ (.B(_1861_),
    .C(_1863_),
    .A(_1858_),
    .Y(_1866_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1865_));
 sg13g2_o21ai_1 _2450_ (.B1(_1846_),
    .VDD(VPWR),
    .Y(_1867_),
    .VSS(VGND),
    .A1(_1855_),
    .A2(_1866_));
 sg13g2_or2_1 _2451_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1868_),
    .B(_1867_),
    .A(_1768_));
 sg13g2_a21oi_1 _2452_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net741),
    .A2(net721),
    .Y(_1869_),
    .B1(_1579_));
 sg13g2_o21ai_1 _2453_ (.B1(_1578_),
    .VDD(VPWR),
    .Y(_1870_),
    .VSS(VGND),
    .A1(net740),
    .A2(net722));
 sg13g2_nor4_1 _2454_ (.A(_1627_),
    .B(_1648_),
    .C(_1654_),
    .D(_1699_),
    .Y(_1871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2455_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net764),
    .A2(_1686_),
    .Y(_1872_),
    .B1(_1633_));
 sg13g2_o21ai_1 _2456_ (.B1(net716),
    .VDD(VPWR),
    .Y(_1873_),
    .VSS(VGND),
    .A1(_1660_),
    .A2(_1872_));
 sg13g2_nor2_1 _2457_ (.A(_1605_),
    .B(_1723_),
    .Y(_1874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2458_ (.A(_1554_),
    .B(net751),
    .C(_1571_),
    .Y(_1875_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1611_));
 sg13g2_a22oi_1 _2459_ (.Y(_1876_),
    .B1(_1703_),
    .B2(_1731_),
    .A2(_1699_),
    .A1(_1684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2460_ (.A(_1493_),
    .B(_1876_),
    .Y(_1877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2461_ (.A(_1873_),
    .B(_1874_),
    .C(_1875_),
    .D(_1877_),
    .Y(_1878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2462_ (.B1(_1878_),
    .VDD(VPWR),
    .Y(_1879_),
    .VSS(VGND),
    .A1(_1634_),
    .A2(_1871_));
 sg13g2_nand2_1 _2463_ (.Y(_1880_),
    .A(_1602_),
    .B(_1829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2464_ (.B(_1879_),
    .C(_1880_),
    .A(_1759_),
    .Y(_1881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2465_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1592_),
    .A2(net723),
    .Y(_1882_),
    .B1(net741));
 sg13g2_a21oi_1 _2466_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1881_),
    .A2(_1882_),
    .Y(_1883_),
    .B1(_1870_));
 sg13g2_or2_1 _2467_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1884_),
    .B(_1883_),
    .A(net718));
 sg13g2_nor3_1 _2468_ (.A(_1569_),
    .B(_1617_),
    .C(_1723_),
    .Y(_1885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2469_ (.A(_1600_),
    .B(net725),
    .Y(_1886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2470_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1887_),
    .B(_1876_),
    .A(net764));
 sg13g2_nand3_1 _2471_ (.B(_1612_),
    .C(_1635_),
    .A(_1557_),
    .Y(_1888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2472_ (.B1(net734),
    .VDD(VPWR),
    .Y(_1889_),
    .VSS(VGND),
    .A1(_1629_),
    .A2(_1684_));
 sg13g2_a21oi_1 _2473_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net734),
    .A2(_1684_),
    .Y(_1890_),
    .B1(_1602_));
 sg13g2_nand4_1 _2474_ (.B(_1887_),
    .C(_1888_),
    .A(net716),
    .Y(_1891_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1889_));
 sg13g2_o21ai_1 _2475_ (.B1(_1891_),
    .VDD(VPWR),
    .Y(_1892_),
    .VSS(VGND),
    .A1(_1601_),
    .A2(_1886_));
 sg13g2_nor2_1 _2476_ (.A(net729),
    .B(_1616_),
    .Y(_1893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2477_ (.A(net729),
    .B(_1617_),
    .Y(_1894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2478_ (.Y(_1895_),
    .A(_1592_),
    .B(_1629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2479_ (.Y(_1896_),
    .A(net719),
    .B(_1895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2480_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1564_),
    .A2(_1894_),
    .Y(_1897_),
    .B1(_1896_));
 sg13g2_a21oi_1 _2481_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1759_),
    .A2(_1892_),
    .Y(_1898_),
    .B1(_1897_));
 sg13g2_a21oi_2 _2482_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1885_),
    .Y(_1899_),
    .A2(_1898_),
    .A1(_1569_));
 sg13g2_inv_2 _2483_ (.Y(_1900_),
    .A(net695),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2484_ (.A(net774),
    .B(net695),
    .Y(_1901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2485_ (.A(net752),
    .B(_1636_),
    .C(_1693_),
    .Y(_1902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2486_ (.Y(_1903_),
    .A(\sap_3_inst.alu_flags[7] ),
    .B(_1902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2487_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net695),
    .A2(_1903_),
    .Y(_1904_),
    .B1(_1901_));
 sg13g2_a21oi_1 _2488_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net8),
    .A2(_1884_),
    .Y(_1905_),
    .B1(_1904_));
 sg13g2_a22oi_1 _2489_ (.Y(_1906_),
    .B1(net614),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .A2(net618),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2490_ (.Y(_1907_),
    .B1(net628),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .A2(net631),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2491_ (.Y(_1908_),
    .A(_1906_),
    .B(_1907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2492_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .C1(net620),
    .B1(net600),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .Y(_1909_),
    .A2(net711));
 sg13g2_a22oi_1 _2493_ (.Y(_1910_),
    .B1(net616),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .A2(net624),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2494_ (.Y(_1911_),
    .B1(net622),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .A2(net601),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2495_ (.B(_1910_),
    .C(_1911_),
    .A(_1909_),
    .Y(_1912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2496_ (.B1(net576),
    .VDD(VPWR),
    .Y(_1913_),
    .VSS(VGND),
    .A1(_1908_),
    .A2(_1912_));
 sg13g2_nand3_1 _2497_ (.B(_1905_),
    .C(_1913_),
    .A(_1868_),
    .Y(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2498_ (.A(net24),
    .Y(_1914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2499_ (.A(net752),
    .B(_1628_),
    .C(net721),
    .Y(_1915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2500_ (.B(_1627_),
    .C(net722),
    .A(_1557_),
    .Y(_1916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2501_ (.A(\sap_3_inst.alu_flags[7] ),
    .B(_1915_),
    .Y(_1917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2502_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1914_),
    .A2(_1915_),
    .Y(_0032_),
    .B1(_1917_));
 sg13g2_nand2_1 _2503_ (.Y(_1918_),
    .A(_1539_),
    .B(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2504_ (.B(net667),
    .C(net626),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ),
    .Y(_1919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2505_ (.Y(_1920_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .B(net711),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2506_ (.Y(_1921_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2507_ (.B(net697),
    .C(net626),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .Y(_1922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2508_ (.Y(_1923_),
    .B1(net614),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .A2(net618),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2509_ (.Y(_1924_),
    .B1(net616),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .A2(net622),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2510_ (.B(_1920_),
    .C(_1921_),
    .A(_1919_),
    .Y(_1925_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1922_));
 sg13g2_a221oi_1 _2511_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .C1(net631),
    .B1(net621),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .Y(_1926_),
    .A2(net624));
 sg13g2_nand3_1 _2512_ (.B(_1924_),
    .C(_1926_),
    .A(_1923_),
    .Y(_1927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2513_ (.B1(_1918_),
    .VDD(VPWR),
    .Y(_1928_),
    .VSS(VGND),
    .A1(_1925_),
    .A2(_1927_));
 sg13g2_or2_1 _2514_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1929_),
    .B(_1928_),
    .A(_1768_));
 sg13g2_or2_1 _2515_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1930_),
    .B(_1899_),
    .A(net777));
 sg13g2_a21o_1 _2516_ (.A2(_1902_),
    .A1(\sap_3_inst.alu_flags[6] ),
    .B1(_1900_),
    .X(_1931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2517_ (.Y(_1932_),
    .B1(_1930_),
    .B2(_1931_),
    .A2(_1884_),
    .A1(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2518_ (.Y(_1933_),
    .B1(net614),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .A2(net600),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2519_ (.Y(_1934_),
    .B1(net624),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .A2(net631),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2520_ (.Y(_1935_),
    .A(_1933_),
    .B(_1934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2521_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .C1(net621),
    .B1(net601),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ),
    .Y(_1936_),
    .A2(net711));
 sg13g2_a22oi_1 _2522_ (.Y(_1937_),
    .B1(net622),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .A2(net628),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2523_ (.Y(_1938_),
    .B1(net616),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .A2(net618),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2524_ (.B(_1937_),
    .C(_1938_),
    .A(_1936_),
    .Y(_1939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2525_ (.B1(net576),
    .VDD(VPWR),
    .Y(_1940_),
    .VSS(VGND),
    .A1(_1935_),
    .A2(_1939_));
 sg13g2_and3_2 _2526_ (.X(_1941_),
    .A(_1929_),
    .B(_1932_),
    .C(_1940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2527_ (.Y(net23),
    .A(net570),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2528_ (.A(\sap_3_inst.alu_flags[6] ),
    .B(net710),
    .Y(_1942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2529_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net710),
    .A2(net570),
    .Y(_0031_),
    .B1(_1942_));
 sg13g2_nand2b_1 _2530_ (.Y(_1943_),
    .B(net632),
    .A_N(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2531_ (.B(net667),
    .C(net626),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ),
    .Y(_1944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2532_ (.Y(_1945_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .B(net621),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2533_ (.Y(_1946_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .B(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2534_ (.B(net697),
    .C(net626),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .Y(_1947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2535_ (.Y(_1948_),
    .B1(net625),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .A2(net628),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2536_ (.B(_1947_),
    .C(_1948_),
    .A(_1945_),
    .Y(_1949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2537_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .C1(net632),
    .B1(_1860_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .Y(_1950_),
    .A2(_1859_));
 sg13g2_a22oi_1 _2538_ (.Y(_1951_),
    .B1(net615),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .A2(_1853_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2539_ (.B(_1946_),
    .C(_1950_),
    .A(_1944_),
    .Y(_1952_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1951_));
 sg13g2_o21ai_1 _2540_ (.B1(_1943_),
    .VDD(VPWR),
    .Y(_1953_),
    .VSS(VGND),
    .A1(_1949_),
    .A2(_1952_));
 sg13g2_nor2_1 _2541_ (.A(_1768_),
    .B(_1953_),
    .Y(_1954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2542_ (.A(net780),
    .B(net695),
    .Y(_1955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2543_ (.Y(_1956_),
    .A(\sap_3_inst.alu_flags[5] ),
    .B(_1902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2544_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net695),
    .A2(_1956_),
    .Y(_1957_),
    .B1(_1955_));
 sg13g2_and2_1 _2545_ (.A(net6),
    .B(_1884_),
    .X(_1958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2546_ (.Y(_1959_),
    .B1(net614),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .A2(net618),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2547_ (.Y(_1960_),
    .B1(_1862_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .A2(net617),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2548_ (.Y(_1961_),
    .B1(net625),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .A2(net712),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2549_ (.Y(_1962_),
    .B1(net622),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .A2(net632),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2550_ (.A(_1959_),
    .B(_1962_),
    .X(_1963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2551_ (.Y(_1964_),
    .B1(net601),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .A2(net628),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2552_ (.A(_1857_),
    .B(_1960_),
    .C(_1963_),
    .D(_1964_),
    .X(_1965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2553_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1961_),
    .A2(_1965_),
    .Y(_1966_),
    .B1(_1720_));
 sg13g2_nor4_2 _2554_ (.A(_1954_),
    .B(_1957_),
    .C(_1958_),
    .Y(_1967_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1966_));
 sg13g2_inv_2 _2555_ (.Y(net22),
    .A(net569),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2556_ (.A(\sap_3_inst.alu_flags[5] ),
    .B(net710),
    .Y(_1968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2557_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net710),
    .A2(net569),
    .Y(_0030_),
    .B1(_1968_));
 sg13g2_nand2b_1 _2558_ (.Y(_1969_),
    .B(net632),
    .A_N(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2559_ (.Y(_1970_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .B(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2560_ (.Y(_1971_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .B(net621),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2561_ (.Y(_1972_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .B(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2562_ (.Y(_1973_),
    .B1(net616),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .A2(net628),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2563_ (.Y(_1974_),
    .B1(net600),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .A2(net624),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2564_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .A2(net614),
    .Y(_1975_),
    .B1(net631));
 sg13g2_a22oi_1 _2565_ (.Y(_1976_),
    .B1(net618),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .A2(net711),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2566_ (.A(_1971_),
    .B(_1973_),
    .C(_1975_),
    .D(_1976_),
    .X(_1977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2567_ (.B(_1972_),
    .C(_1974_),
    .A(_1970_),
    .Y(_1978_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1977_));
 sg13g2_nand3b_1 _2568_ (.B(_1969_),
    .C(_1978_),
    .Y(_1979_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1768_));
 sg13g2_nand2_1 _2569_ (.Y(_1980_),
    .A(_1509_),
    .B(_1900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2570_ (.A2(_1902_),
    .A1(\sap_3_inst.alu_flags[4] ),
    .B1(_1900_),
    .X(_1981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2571_ (.Y(_1982_),
    .B1(_1980_),
    .B2(_1981_),
    .A2(_1884_),
    .A1(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2572_ (.Y(_1983_),
    .B1(net616),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .A2(net628),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2573_ (.Y(_1984_),
    .A(_1857_),
    .B(_1983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2574_ (.Y(_1985_),
    .B1(net614),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .A2(net624),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2575_ (.Y(_1986_),
    .B1(net600),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .A2(net622),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2576_ (.Y(_1987_),
    .B1(net618),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .A2(net631),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2577_ (.Y(_1988_),
    .B1(net601),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .A2(net711),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2578_ (.B(_1986_),
    .C(_1987_),
    .A(_1985_),
    .Y(_1989_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1988_));
 sg13g2_o21ai_1 _2579_ (.B1(net576),
    .VDD(VPWR),
    .Y(_1990_),
    .VSS(VGND),
    .A1(_1984_),
    .A2(_1989_));
 sg13g2_nand3_1 _2580_ (.B(_1982_),
    .C(_1990_),
    .A(_1979_),
    .Y(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2581_ (.A(net21),
    .Y(_1991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2582_ (.A(\sap_3_inst.alu_flags[4] ),
    .B(net710),
    .Y(_1992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2583_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net710),
    .A2(_1991_),
    .Y(_0029_),
    .B1(_1992_));
 sg13g2_nand2_1 _2584_ (.Y(_1993_),
    .A(_1598_),
    .B(_1612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2585_ (.A(_1605_),
    .B(net725),
    .Y(_1994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2586_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1496_),
    .C1(_1994_),
    .B1(_1894_),
    .A1(_1595_),
    .Y(_1995_),
    .A2(net722));
 sg13g2_o21ai_1 _2587_ (.B1(_1993_),
    .VDD(VPWR),
    .Y(_1996_),
    .VSS(VGND),
    .A1(_1602_),
    .A2(_1995_));
 sg13g2_nand2_1 _2588_ (.Y(_1997_),
    .A(_1592_),
    .B(_1612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2589_ (.B1(_1723_),
    .VDD(VPWR),
    .Y(_1998_),
    .VSS(VGND),
    .A1(net728),
    .A2(_1762_));
 sg13g2_nand2b_1 _2590_ (.Y(_1999_),
    .B(_1998_),
    .A_N(_1600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2591_ (.B1(_1997_),
    .VDD(VPWR),
    .Y(_2000_),
    .VSS(VGND),
    .A1(_1760_),
    .A2(_1999_));
 sg13g2_a21oi_1 _2592_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net725),
    .A2(_1673_),
    .Y(_2001_),
    .B1(net733));
 sg13g2_nor3_2 _2593_ (.A(_1996_),
    .B(net704),
    .C(_2001_),
    .Y(_2002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2594_ (.Y(_2003_),
    .A(_1916_),
    .B(_2002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2595_ (.A(net757),
    .B(_1996_),
    .X(_2004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2596_ (.Y(_2005_),
    .A(net757),
    .B(_1996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2597_ (.A(_1494_),
    .B(_1571_),
    .C(net728),
    .D(_1616_),
    .Y(_2006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2598_ (.B(_1570_),
    .C(_1893_),
    .A(net765),
    .Y(_2007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2599_ (.A(net731),
    .B(_1618_),
    .X(_2008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2600_ (.A(_1571_),
    .B(net728),
    .C(_1617_),
    .Y(_2009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2601_ (.Y(_2010_),
    .A(_2005_),
    .B(_2007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2602_ (.A(net704),
    .B(_2010_),
    .Y(_2011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2603_ (.A(_2005_),
    .B(_2009_),
    .Y(_2012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2604_ (.Y(_2013_),
    .A(_2004_),
    .B(_2007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2605_ (.A(_1600_),
    .B(_1831_),
    .Y(_2014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2606_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net762),
    .A2(_1996_),
    .Y(_2015_),
    .B1(_2014_));
 sg13g2_a221oi_1 _2607_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net762),
    .C1(_2014_),
    .B1(_1996_),
    .A1(net734),
    .Y(_2016_),
    .A2(_1672_));
 sg13g2_o21ai_1 _2608_ (.B1(_2015_),
    .VDD(VPWR),
    .Y(_2017_),
    .VSS(VGND),
    .A1(net733),
    .A2(_1673_));
 sg13g2_and2_1 _2609_ (.A(net760),
    .B(_1996_),
    .X(_2018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2610_ (.Y(_2019_),
    .A(_2016_),
    .B(_2018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2611_ (.Y(_2020_),
    .A(_1655_),
    .B(_1996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2612_ (.B1(_2019_),
    .VDD(VPWR),
    .Y(_2021_),
    .VSS(VGND),
    .A1(net760),
    .A2(_2013_));
 sg13g2_a21oi_1 _2613_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2008_),
    .A2(_2020_),
    .Y(_2022_),
    .B1(_2021_));
 sg13g2_nor2b_1 _2614_ (.A(_2011_),
    .B_N(_2022_),
    .Y(_2023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2615_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1916_),
    .A2(_2002_),
    .Y(_2024_),
    .B1(_2023_));
 sg13g2_nand2_1 _2616_ (.Y(_2025_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .B(net629),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2617_ (.Y(_2026_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .B(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2618_ (.B(net696),
    .C(net627),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .Y(_2027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2619_ (.B(net667),
    .C(net627),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .Y(_2028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2620_ (.Y(_2029_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .B(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2621_ (.Y(_2030_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ),
    .B(net619),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2622_ (.A(_2026_),
    .B(_2028_),
    .C(_2029_),
    .D(_2030_),
    .X(_2031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2623_ (.Y(_2032_),
    .B1(net615),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ),
    .A2(net617),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2624_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .C1(net630),
    .B1(net624),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .Y(_2033_),
    .A2(net713));
 sg13g2_and4_1 _2625_ (.A(_2025_),
    .B(_2027_),
    .C(_2032_),
    .D(_2033_),
    .X(_2034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2626_ (.Y(_2035_),
    .B1(_2031_),
    .B2(_2034_),
    .A2(net630),
    .A1(_1510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2627_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2034_),
    .C1(_1768_),
    .B1(_2031_),
    .A1(_1510_),
    .Y(_2036_),
    .A2(net630));
 sg13g2_nor2_1 _2628_ (.A(net791),
    .B(net695),
    .Y(_2037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2629_ (.Y(_2038_),
    .A(net748),
    .B(_1902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net695),
    .A2(_2038_),
    .Y(_2039_),
    .B1(_2037_));
 sg13g2_and2_1 _2631_ (.A(net2),
    .B(_1884_),
    .X(_2040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2632_ (.Y(_2041_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .B(net630),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2633_ (.B(net667),
    .C(net627),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .Y(_2042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2634_ (.Y(_2043_),
    .B1(net617),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .A2(net619),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2635_ (.X(_2044_),
    .A(_2041_),
    .B(_2042_),
    .C(_2043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2636_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .C1(net620),
    .B1(net629),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ),
    .Y(_2045_),
    .A2(net713));
 sg13g2_nand2_1 _2637_ (.Y(_2046_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .B(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2638_ (.B(net696),
    .C(net627),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .Y(_2047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2639_ (.Y(_2048_),
    .B1(net615),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .A2(net624),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2640_ (.A(_2045_),
    .B(_2046_),
    .C(_2047_),
    .D(_2048_),
    .X(_2049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2641_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2044_),
    .A2(_2049_),
    .Y(_2050_),
    .B1(_1720_));
 sg13g2_nor4_2 _2642_ (.A(_2036_),
    .B(_2039_),
    .C(_2040_),
    .Y(_2051_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_2050_));
 sg13g2_inv_2 _2643_ (.Y(net18),
    .A(_2051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2644_ (.B1(_2024_),
    .VDD(VPWR),
    .Y(_2052_),
    .VSS(VGND),
    .A1(\sap_3_inst.alu_inst.carry ),
    .A2(net710));
 sg13g2_a21o_1 _2645_ (.A2(_2051_),
    .A1(net710),
    .B1(_2052_),
    .X(_2053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2646_ (.B1(_2053_),
    .VDD(VPWR),
    .Y(_0028_),
    .VSS(VGND),
    .A1(_1487_),
    .A2(_2024_));
 sg13g2_nand2_2 _2647_ (.Y(_2054_),
    .A(_2017_),
    .B(_2018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2648_ (.Y(_2055_),
    .A(_2012_),
    .B(_2054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2649_ (.Y(_2056_),
    .A(_2010_),
    .B(_2055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2650_ (.Y(_2057_),
    .A(_2003_),
    .B(_2056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2651_ (.Y(_2058_),
    .A(\sap_3_inst.alu_flags[3] ),
    .B(_2057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2652_ (.Y(_2059_),
    .A(_1497_),
    .B(net632),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2653_ (.B(net697),
    .C(net626),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .Y(_2060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2654_ (.B(_1809_),
    .C(net626),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .Y(_2061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2655_ (.Y(_2062_),
    .B1(_1864_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .A2(net625),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2656_ (.B(_2061_),
    .C(_2062_),
    .A(_2060_),
    .Y(_2063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2657_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .C1(net632),
    .B1(net616),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .Y(_2064_),
    .A2(net712));
 sg13g2_a22oi_1 _2658_ (.Y(_2065_),
    .B1(net618),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ),
    .A2(net621),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2659_ (.Y(_2066_),
    .B1(net622),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .A2(_1847_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2660_ (.B(_2065_),
    .C(_2066_),
    .A(_2064_),
    .Y(_2067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2661_ (.B1(_2059_),
    .VDD(VPWR),
    .Y(_2068_),
    .VSS(VGND),
    .A1(_2063_),
    .A2(_2067_));
 sg13g2_or2_1 _2662_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0196_),
    .B(_2068_),
    .A(_1768_));
 sg13g2_a22oi_1 _2663_ (.Y(_0197_),
    .B1(net614),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .A2(net622),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2664_ (.Y(_0198_),
    .B1(net616),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .A2(net625),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2665_ (.Y(_0199_),
    .A(_0197_),
    .B(_0198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2666_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .C1(net620),
    .B1(net601),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ),
    .Y(_0200_),
    .A2(net712));
 sg13g2_a22oi_1 _2667_ (.Y(_0201_),
    .B1(net600),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .A2(net629),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2668_ (.Y(_0202_),
    .B1(net618),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .A2(net632),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2669_ (.B(_0201_),
    .C(_0202_),
    .A(_0200_),
    .Y(_0203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2670_ (.B1(net577),
    .VDD(VPWR),
    .Y(_0204_),
    .VSS(VGND),
    .A1(_0199_),
    .A2(_0203_));
 sg13g2_nand2_1 _2671_ (.Y(_0205_),
    .A(\sap_3_inst.alu_flags[3] ),
    .B(_1902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2672_ (.Y(_0206_),
    .B1(_1900_),
    .B2(net785),
    .A2(_1884_),
    .A1(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2673_ (.B(_0204_),
    .C(_0205_),
    .A(_0196_),
    .Y(net20),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0206_));
 sg13g2_nand2b_1 _2674_ (.Y(_0207_),
    .B(_1916_),
    .A_N(net774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2675_ (.B1(_0207_),
    .VDD(VPWR),
    .Y(_0208_),
    .VSS(VGND),
    .A1(_1916_),
    .A2(net32));
 sg13g2_o21ai_1 _2676_ (.B1(_2058_),
    .VDD(VPWR),
    .Y(_0027_),
    .VSS(VGND),
    .A1(_2057_),
    .A2(_0208_));
 sg13g2_a22oi_1 _2677_ (.Y(_0209_),
    .B1(net615),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .A2(net625),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2678_ (.Y(_0210_),
    .B1(net620),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .A2(net623),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2679_ (.A(_0209_),
    .B(_0210_),
    .X(_0211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2680_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .C1(net630),
    .B1(net629),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .Y(_0212_),
    .A2(net711));
 sg13g2_a22oi_1 _2681_ (.Y(_0213_),
    .B1(net600),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .A2(net619),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2682_ (.Y(_0214_),
    .B1(net617),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .A2(net601),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2683_ (.X(_0215_),
    .A(_0212_),
    .B(_0213_),
    .C(_0214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2684_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0215_),
    .C1(_1768_),
    .B1(_0211_),
    .A1(_1501_),
    .Y(_0216_),
    .A2(net633));
 sg13g2_a21oi_1 _2685_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu_flags[2] ),
    .A2(_1902_),
    .Y(_0217_),
    .B1(_1900_));
 sg13g2_a21oi_1 _2686_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1500_),
    .A2(_1900_),
    .Y(_0218_),
    .B1(_0217_));
 sg13g2_and2_1 _2687_ (.A(net3),
    .B(_1884_),
    .X(_0219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2688_ (.Y(_0220_),
    .B1(net601),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .A2(net629),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2689_ (.Y(_0221_),
    .B1(net600),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .A2(net619),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2690_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .C1(net620),
    .B1(net615),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .Y(_0222_),
    .A2(net625));
 sg13g2_a22oi_1 _2691_ (.Y(_0223_),
    .B1(net617),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .A2(net711),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2692_ (.Y(_0224_),
    .B1(net623),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .A2(net630),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2693_ (.A(_0220_),
    .B(_0221_),
    .C(_0223_),
    .D(_0224_),
    .X(_0225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2694_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0222_),
    .A2(_0225_),
    .Y(_0226_),
    .B1(_1720_));
 sg13g2_or4_1 _2695_ (.A(_0216_),
    .B(_0218_),
    .C(_0219_),
    .D(_0226_),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2696_ (.A(net19),
    .Y(_0227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2697_ (.Y(_0228_),
    .A(net774),
    .B(net777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2698_ (.B(net782),
    .A(net780),
    .X(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2699_ (.Y(_0230_),
    .A(_0228_),
    .B(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2700_ (.B(net793),
    .A(net791),
    .X(_0231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2701_ (.B(net788),
    .A(net785),
    .X(_0232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2702_ (.Y(_0233_),
    .A(_0231_),
    .B(_0232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2703_ (.Y(_0234_),
    .A(_0230_),
    .B(_0233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2704_ (.Y(_0235_),
    .A(_1916_),
    .B(_0234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2705_ (.B1(_0235_),
    .VDD(VPWR),
    .Y(_0236_),
    .VSS(VGND),
    .A1(_1916_),
    .A2(net19));
 sg13g2_nand2_1 _2706_ (.Y(_0237_),
    .A(\sap_3_inst.alu_flags[2] ),
    .B(_2057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2707_ (.B1(_0237_),
    .VDD(VPWR),
    .Y(_0026_),
    .VSS(VGND),
    .A1(_2057_),
    .A2(_0236_));
 sg13g2_o21ai_1 _2708_ (.B1(_2003_),
    .VDD(VPWR),
    .Y(_0238_),
    .VSS(VGND),
    .A1(_1492_),
    .A2(net754));
 sg13g2_nand2b_1 _2709_ (.Y(_0239_),
    .B(net633),
    .A_N(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2710_ (.Y(_0240_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .B(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2711_ (.B(_1809_),
    .C(net627),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ),
    .Y(_0241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2712_ (.Y(_0242_),
    .B1(net617),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .A2(net625),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2713_ (.B(_0241_),
    .C(_0242_),
    .A(_0240_),
    .Y(_0243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2714_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .C1(net630),
    .B1(net629),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ),
    .Y(_0244_),
    .A2(net712));
 sg13g2_a22oi_1 _2715_ (.Y(_0245_),
    .B1(net619),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ),
    .A2(net620),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2716_ (.Y(_0246_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .B(net615),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2717_ (.B(net697),
    .C(net627),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .Y(_0247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2718_ (.B(_0245_),
    .C(_0246_),
    .A(_0244_),
    .Y(_0248_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0247_));
 sg13g2_o21ai_1 _2719_ (.B1(_0239_),
    .VDD(VPWR),
    .Y(_0249_),
    .VSS(VGND),
    .A1(_0243_),
    .A2(_0248_));
 sg13g2_or2_1 _2720_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0250_),
    .B(_0249_),
    .A(_1768_));
 sg13g2_nor2_1 _2721_ (.A(net793),
    .B(net695),
    .Y(_0251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2722_ (.Y(_0252_),
    .A(\sap_3_inst.alu_flags[0] ),
    .B(_1902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2723_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1899_),
    .A2(_0252_),
    .Y(_0253_),
    .B1(_0251_));
 sg13g2_a21oi_1 _2724_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1),
    .A2(_1884_),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_a22oi_1 _2725_ (.Y(_0255_),
    .B1(net619),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .A2(net623),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2726_ (.Y(_0256_),
    .B1(net625),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .A2(net629),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2727_ (.Y(_0257_),
    .A(_0255_),
    .B(_0256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2728_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .C1(net620),
    .B1(_1850_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ),
    .Y(_0258_),
    .A2(net712));
 sg13g2_a22oi_1 _2729_ (.Y(_0259_),
    .B1(net600),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .A2(net630),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2730_ (.Y(_0260_),
    .B1(net615),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ),
    .A2(net617),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2731_ (.B(_0259_),
    .C(_0260_),
    .A(_0258_),
    .Y(_0261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2732_ (.B1(net577),
    .VDD(VPWR),
    .Y(_0262_),
    .VSS(VGND),
    .A1(_0257_),
    .A2(_0261_));
 sg13g2_nand3_1 _2733_ (.B(_0254_),
    .C(_0262_),
    .A(_0250_),
    .Y(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2734_ (.A(net774),
    .B(net780),
    .C(net782),
    .D(net777),
    .Y(_0263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2735_ (.A(net785),
    .B(net788),
    .C(net791),
    .D(net793),
    .Y(_0264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2736_ (.B(_0263_),
    .C(_0264_),
    .A(_2056_),
    .Y(_0265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2737_ (.A(\sap_3_inst.alu_inst.act[5] ),
    .B(\sap_3_inst.alu_inst.act[4] ),
    .C(\sap_3_inst.alu_inst.act[7] ),
    .D(\sap_3_inst.alu_inst.act[6] ),
    .Y(_0266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2738_ (.A(\sap_3_inst.alu_inst.act[1] ),
    .B(\sap_3_inst.alu_inst.act[0] ),
    .C(\sap_3_inst.alu_inst.act[3] ),
    .D(\sap_3_inst.alu_inst.act[2] ),
    .Y(_0267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2739_ (.Y(_0268_),
    .A(_0266_),
    .B(_0267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2740_ (.B1(_0265_),
    .VDD(VPWR),
    .Y(_0269_),
    .VSS(VGND),
    .A1(_2056_),
    .A2(_0268_));
 sg13g2_mux2_1 _2741_ (.A0(net31),
    .A1(_0269_),
    .S(_1916_),
    .X(_0270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2742_ (.A0(_0270_),
    .A1(\sap_3_inst.alu_flags[0] ),
    .S(_0238_),
    .X(_0025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2743_ (.A(_1730_),
    .B(_1748_),
    .C(_1754_),
    .D(net719),
    .Y(_0271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2744_ (.B(_1887_),
    .C(_0271_),
    .A(_1798_),
    .Y(_0272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2745_ (.Y(_0273_),
    .B1(_1896_),
    .B2(_0272_),
    .A2(net722),
    .A1(net739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2746_ (.A(_1579_),
    .B(_0273_),
    .Y(mem_ram_we),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2747_ (.B(_1667_),
    .C(_1893_),
    .A(_1626_),
    .Y(_0274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2748_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net726),
    .A2(_1682_),
    .Y(_0275_),
    .B1(_1650_));
 sg13g2_o21ai_1 _2749_ (.B1(_1690_),
    .VDD(VPWR),
    .Y(_0276_),
    .VSS(VGND),
    .A1(net731),
    .A2(_1692_));
 sg13g2_o21ai_1 _2750_ (.B1(_0276_),
    .VDD(VPWR),
    .Y(_0277_),
    .VSS(VGND),
    .A1(_1666_),
    .A2(_1676_));
 sg13g2_o21ai_1 _2751_ (.B1(_1670_),
    .VDD(VPWR),
    .Y(_0278_),
    .VSS(VGND),
    .A1(_0275_),
    .A2(_0277_));
 sg13g2_nand2b_1 _2752_ (.Y(_0279_),
    .B(_1612_),
    .A_N(_1607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2753_ (.B1(_1692_),
    .VDD(VPWR),
    .Y(_0280_),
    .VSS(VGND),
    .A1(_1627_),
    .A2(_1635_));
 sg13g2_a21oi_1 _2754_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net705),
    .A2(_0280_),
    .Y(_0281_),
    .B1(_1651_));
 sg13g2_nand2_1 _2755_ (.Y(_0282_),
    .A(_1639_),
    .B(_1692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2756_ (.A(_1620_),
    .B(_1876_),
    .C(_0279_),
    .D(_0282_),
    .X(_0283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2757_ (.B1(_0283_),
    .VDD(VPWR),
    .Y(_0284_),
    .VSS(VGND),
    .A1(_1647_),
    .A2(_1673_));
 sg13g2_o21ai_1 _2758_ (.B1(_1835_),
    .VDD(VPWR),
    .Y(_0285_),
    .VSS(VGND),
    .A1(net735),
    .A2(_1682_));
 sg13g2_nor4_1 _2759_ (.A(_1707_),
    .B(_0281_),
    .C(_0284_),
    .D(_0285_),
    .Y(_0286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2760_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1608_),
    .A2(_1731_),
    .Y(_0287_),
    .B1(_1620_));
 sg13g2_nand2b_2 _2761_ (.Y(_0288_),
    .B(_0287_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1994_));
 sg13g2_a221oi_1 _2762_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1995_),
    .C1(_1602_),
    .B1(_0287_),
    .A1(_0278_),
    .Y(_0289_),
    .A2(_0286_));
 sg13g2_nor2_1 _2763_ (.A(net716),
    .B(net725),
    .Y(_0290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2764_ (.A(net728),
    .B(_1600_),
    .C(_1762_),
    .Y(_0291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2765_ (.A(_1760_),
    .B(_0289_),
    .C(_0290_),
    .D(_0291_),
    .Y(_0292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2766_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net731),
    .A2(_1758_),
    .Y(_0293_),
    .B1(_1896_));
 sg13g2_nor4_1 _2767_ (.A(net742),
    .B(net739),
    .C(_0292_),
    .D(_0293_),
    .Y(_0294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2768_ (.B1(net723),
    .VDD(VPWR),
    .Y(_0295_),
    .VSS(VGND),
    .A1(net742),
    .A2(_1568_));
 sg13g2_nand3b_1 _2769_ (.B(_0295_),
    .C(_1578_),
    .Y(_0296_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0294_));
 sg13g2_o21ai_1 _2770_ (.B1(_0296_),
    .VDD(VPWR),
    .Y(_0297_),
    .VSS(VGND),
    .A1(net751),
    .A2(_1569_));
 sg13g2_a21o_1 _2771_ (.A2(_1581_),
    .A1(net743),
    .B1(_0297_),
    .X(_0298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2772_ (.A(_1491_),
    .B(_0298_),
    .X(_0001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2773_ (.A(_1587_),
    .B_N(_0298_),
    .Y(_0002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2774_ (.B1(_0297_),
    .VDD(VPWR),
    .Y(_0299_),
    .VSS(VGND),
    .A1(net745),
    .A2(_1580_));
 sg13g2_nor2b_1 _2775_ (.A(_0299_),
    .B_N(_1681_),
    .Y(_0003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2776_ (.Y(_0300_),
    .B(_1681_),
    .A_N(net744),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2777_ (.X(_0004_),
    .A(_1682_),
    .B(_0297_),
    .C(_0300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2778_ (.Y(_0301_),
    .B(net577),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0249_));
 sg13g2_inv_1 _2779_ (.VDD(VPWR),
    .Y(net9),
    .A(_0301_),
    .VSS(VGND));
 sg13g2_nand2_2 _2780_ (.Y(_0302_),
    .A(net576),
    .B(_2035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2781_ (.VDD(VPWR),
    .Y(net10),
    .A(_0302_),
    .VSS(VGND));
 sg13g2_a221oi_1 _2782_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0215_),
    .C1(_1720_),
    .B1(_0211_),
    .A1(_1501_),
    .Y(net11),
    .A2(net633));
 sg13g2_nand2b_2 _2783_ (.Y(_0303_),
    .B(net577),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2068_));
 sg13g2_inv_1 _2784_ (.VDD(VPWR),
    .Y(net12),
    .A(_0303_),
    .VSS(VGND));
 sg13g2_and3_2 _2785_ (.X(net13),
    .A(net576),
    .B(_1969_),
    .C(_1978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2786_ (.Y(_0304_),
    .B(net576),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1953_));
 sg13g2_inv_2 _2787_ (.Y(net14),
    .A(_0304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2788_ (.Y(_0305_),
    .B(net576),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1928_));
 sg13g2_inv_4 _2789_ (.A(_0305_),
    .Y(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2790_ (.Y(_0306_),
    .B(net576),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1867_));
 sg13g2_inv_2 _2791_ (.Y(net16),
    .A(_0306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2792_ (.B(net741),
    .C(net731),
    .A(_1559_),
    .Y(_0000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2793_ (.A(_1651_),
    .B(_1659_),
    .C(_1674_),
    .Y(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2794_ (.A(_1702_),
    .B(_1711_),
    .C(_0307_),
    .Y(_0308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2795_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net726),
    .A2(_0308_),
    .Y(_0309_),
    .B1(_1725_));
 sg13g2_o21ai_1 _2796_ (.B1(net724),
    .VDD(VPWR),
    .Y(_0310_),
    .VSS(VGND),
    .A1(_1650_),
    .A2(_1685_));
 sg13g2_nor2b_1 _2797_ (.A(_1794_),
    .B_N(_0310_),
    .Y(_0311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2798_ (.Y(_0312_),
    .A(_1744_),
    .B(_0311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2799_ (.A(net714),
    .B(_1697_),
    .C(_1704_),
    .D(_1802_),
    .Y(_0313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2800_ (.Y(_0314_),
    .A(_0312_),
    .B(_0313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2801_ (.B1(_1665_),
    .VDD(VPWR),
    .Y(_0315_),
    .VSS(VGND),
    .A1(_0309_),
    .A2(_0314_));
 sg13g2_a21oi_1 _2802_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1620_),
    .A2(_0315_),
    .Y(_0316_),
    .B1(_1622_));
 sg13g2_o21ai_1 _2803_ (.B1(_1590_),
    .VDD(VPWR),
    .Y(_0317_),
    .VSS(VGND),
    .A1(_1599_),
    .A2(_0316_));
 sg13g2_a21oi_1 _2804_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net740),
    .A2(_0317_),
    .Y(_0318_),
    .B1(_1589_));
 sg13g2_or2_1 _2805_ (.VSS(VGND),
    .VDD(VPWR),
    .X(mem_mar_we),
    .B(_0318_),
    .A(_1556_));
 sg13g2_nor2_2 _2806_ (.A(\u_ser.state[0] ),
    .B(\u_ser.state[1] ),
    .Y(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2807_ (.A0(net58),
    .A1(\sap_3_inst.out[0] ),
    .S(net799),
    .X(_0017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2808_ (.A0(net60),
    .A1(\sap_3_inst.out[1] ),
    .S(net799),
    .X(_0018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2809_ (.A0(net56),
    .A1(\sap_3_inst.out[2] ),
    .S(net799),
    .X(_0019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2810_ (.A0(net59),
    .A1(\sap_3_inst.out[3] ),
    .S(net799),
    .X(_0020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2811_ (.A0(net67),
    .A1(\sap_3_inst.out[4] ),
    .S(net799),
    .X(_0021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2812_ (.A0(net76),
    .A1(\sap_3_inst.out[5] ),
    .S(_0185_),
    .X(_0022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2813_ (.A0(net72),
    .A1(\sap_3_inst.out[6] ),
    .S(_0185_),
    .X(_0023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2814_ (.A0(net57),
    .A1(\sap_3_inst.out[7] ),
    .S(net799),
    .X(_0024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2815_ (.B1(_1759_),
    .VDD(VPWR),
    .Y(_0319_),
    .VSS(VGND),
    .A1(net716),
    .A2(_1886_));
 sg13g2_o21ai_1 _2816_ (.B1(_1895_),
    .VDD(VPWR),
    .Y(_0320_),
    .VSS(VGND),
    .A1(_1890_),
    .A2(_0319_));
 sg13g2_nor3_1 _2817_ (.A(_1598_),
    .B(_1760_),
    .C(_1763_),
    .Y(_0321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2818_ (.Y(_0322_),
    .B(net716),
    .A_N(_1773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2819_ (.B1(_1662_),
    .VDD(VPWR),
    .Y(_0323_),
    .VSS(VGND),
    .A1(_1558_),
    .A2(_1628_));
 sg13g2_a221oi_1 _2820_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1731_),
    .C1(_0322_),
    .B1(_0323_),
    .A1(_1761_),
    .Y(_0324_),
    .A2(_1875_));
 sg13g2_nand2b_1 _2821_ (.Y(_0325_),
    .B(_0324_),
    .A_N(_1877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2822_ (.A(_1565_),
    .B(net728),
    .C(_1762_),
    .Y(_0326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2823_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0325_),
    .C1(_0326_),
    .B1(_0321_),
    .A1(_1592_),
    .Y(_0327_),
    .A2(net723));
 sg13g2_nor2_1 _2824_ (.A(net740),
    .B(_1762_),
    .Y(_0328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2825_ (.B(net723),
    .C(_1761_),
    .A(net742),
    .Y(_0329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2826_ (.B1(_0329_),
    .VDD(VPWR),
    .Y(_0330_),
    .VSS(VGND),
    .A1(net742),
    .A2(_0327_));
 sg13g2_nor2_1 _2827_ (.A(net703),
    .B(net694),
    .Y(_0331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2828_ (.Y(_0332_),
    .A(_2002_),
    .B(_0331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2829_ (.A(_2016_),
    .B(_2018_),
    .Y(_0333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2830_ (.B(_2006_),
    .C(_0333_),
    .A(_2004_),
    .Y(_0334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2831_ (.B(_2008_),
    .C(_0333_),
    .A(_2004_),
    .Y(_0335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2832_ (.B(_2009_),
    .C(_0333_),
    .A(_2004_),
    .Y(_0336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2833_ (.A(net704),
    .B_N(_0336_),
    .Y(_0337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2834_ (.B(_2055_),
    .C(_0337_),
    .A(_2004_),
    .Y(_0338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2835_ (.Y(_0339_),
    .A(_2005_),
    .B(_2006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2836_ (.Y(_0340_),
    .A(_0332_),
    .B(_0338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2837_ (.Y(_0341_),
    .A(net792),
    .B(\sap_3_inst.alu_inst.tmp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2838_ (.B(\sap_3_inst.alu_inst.tmp[0] ),
    .A(net792),
    .X(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2839_ (.Y(_0343_),
    .A(net792),
    .B(\sap_3_inst.alu_inst.tmp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2840_ (.A(_2011_),
    .B(_0333_),
    .X(_0344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2841_ (.Y(_0345_),
    .A(_2011_),
    .B(_0333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2842_ (.B(_2016_),
    .C(_2018_),
    .A(_2011_),
    .Y(_0346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2843_ (.VDD(VPWR),
    .Y(_0347_),
    .A(_0346_),
    .VSS(VGND));
 sg13g2_nor2_2 _2844_ (.A(_2010_),
    .B(_2054_),
    .Y(_0348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2845_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0349_),
    .B(_2054_),
    .A(_2010_));
 sg13g2_nand2_1 _2846_ (.Y(_0350_),
    .A(_0346_),
    .B(_0349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2847_ (.A(_0344_),
    .B(_0350_),
    .Y(_0351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2848_ (.Y(_0352_),
    .A(_2005_),
    .B(_2008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2849_ (.A(_2055_),
    .B(_0337_),
    .C(_0351_),
    .D(_0352_),
    .X(_0353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2850_ (.B(_0337_),
    .C(_0351_),
    .A(_2055_),
    .Y(_0354_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0352_));
 sg13g2_nand2_2 _2851_ (.Y(_0355_),
    .A(_2012_),
    .B(_0333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2852_ (.B(net575),
    .C(_0355_),
    .A(_0346_),
    .Y(_0356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2853_ (.A(_2017_),
    .B(_0339_),
    .Y(_0357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2854_ (.A(net748),
    .B(_2018_),
    .X(_0358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2855_ (.A(_2016_),
    .B(_0339_),
    .Y(_0359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2856_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net789),
    .C1(net703),
    .B1(net691),
    .A1(net692),
    .Y(_0360_),
    .A2(_0358_));
 sg13g2_nor2_2 _2857_ (.A(_2013_),
    .B(_2019_),
    .Y(_0361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2858_ (.B1(_0361_),
    .VDD(VPWR),
    .Y(_0362_),
    .VSS(VGND),
    .A1(net793),
    .A2(\sap_3_inst.alu_inst.tmp[0] ));
 sg13g2_nor3_2 _2859_ (.A(net761),
    .B(_2013_),
    .C(_2017_),
    .Y(_0363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2860_ (.Y(_0364_),
    .B(_0363_),
    .A_N(_0341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2861_ (.B(_0362_),
    .C(_0364_),
    .A(_0360_),
    .Y(_0365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2862_ (.Y(_0366_),
    .A(net748),
    .B(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2863_ (.Y(_0367_),
    .B1(_0345_),
    .B2(_0349_),
    .A2(_0343_),
    .A1(_1487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2864_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0367_),
    .C1(_0365_),
    .B1(_0366_),
    .A1(_0342_),
    .Y(_0368_),
    .A2(_0356_));
 sg13g2_o21ai_1 _2865_ (.B1(_0368_),
    .VDD(VPWR),
    .Y(_0369_),
    .VSS(VGND),
    .A1(net792),
    .A2(_0337_));
 sg13g2_a21oi_1 _2866_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1525_),
    .A2(net703),
    .Y(_0370_),
    .B1(net694));
 sg13g2_a221oi_1 _2867_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0370_),
    .C1(net599),
    .B1(_0369_),
    .A1(net31),
    .Y(_0371_),
    .A2(net694));
 sg13g2_a21oi_1 _2868_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1508_),
    .A2(net599),
    .Y(_0033_),
    .B1(_0371_));
 sg13g2_nand2b_1 _2869_ (.Y(_0372_),
    .B(net703),
    .A_N(\sap_3_inst.alu_inst.act[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2870_ (.Y(_0373_),
    .A(net789),
    .B(\sap_3_inst.alu_inst.tmp[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2871_ (.B(\sap_3_inst.alu_inst.tmp[1] ),
    .A(net789),
    .X(_0374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2872_ (.Y(_0375_),
    .B(_0374_),
    .A_N(_0341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2873_ (.B(_0374_),
    .A(_0341_),
    .X(_0376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2874_ (.A(net575),
    .B(_0376_),
    .Y(_0377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2875_ (.A(net793),
    .B_N(\sap_3_inst.alu_inst.tmp[0] ),
    .Y(_0378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2876_ (.Y(_0379_),
    .A(_0374_),
    .B(_0378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _2877_ (.X(_0380_),
    .A(net748),
    .B(_0343_),
    .C(_0379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2878_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net748),
    .A2(_0343_),
    .Y(_0381_),
    .B1(_0379_));
 sg13g2_o21ai_1 _2879_ (.B1(_0348_),
    .VDD(VPWR),
    .Y(_0382_),
    .VSS(VGND),
    .A1(_0380_),
    .A2(_0381_));
 sg13g2_nand3_1 _2880_ (.B(\sap_3_inst.alu_inst.tmp[1] ),
    .C(_0363_),
    .A(net790),
    .Y(_0383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2881_ (.Y(_0384_),
    .A(net792),
    .B(net692),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2882_ (.Y(_0385_),
    .A(net789),
    .B(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2883_ (.B(net709),
    .A(net789),
    .X(_0386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2884_ (.Y(_0387_),
    .A(net792),
    .B(_0386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2885_ (.B1(_2000_),
    .VDD(VPWR),
    .Y(_0388_),
    .VSS(VGND),
    .A1(net792),
    .A2(_0386_));
 sg13g2_inv_1 _2886_ (.VDD(VPWR),
    .Y(_0389_),
    .A(_0388_),
    .VSS(VGND));
 sg13g2_a221oi_1 _2887_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0389_),
    .C1(net703),
    .B1(_0387_),
    .A1(net786),
    .Y(_0390_),
    .A2(net691));
 sg13g2_or2_1 _2888_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0391_),
    .B(_0379_),
    .A(_0346_));
 sg13g2_o21ai_1 _2889_ (.B1(_0361_),
    .VDD(VPWR),
    .Y(_0392_),
    .VSS(VGND),
    .A1(net790),
    .A2(\sap_3_inst.alu_inst.tmp[1] ));
 sg13g2_nand3_1 _2890_ (.B(_0342_),
    .C(_0374_),
    .A(net748),
    .Y(_0393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2891_ (.B1(_0376_),
    .VDD(VPWR),
    .Y(_0394_),
    .VSS(VGND),
    .A1(_1487_),
    .A2(_0343_));
 sg13g2_nand3_1 _2892_ (.B(_0393_),
    .C(_0394_),
    .A(_0344_),
    .Y(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2893_ (.A(_0355_),
    .B_N(_0374_),
    .Y(_0396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2894_ (.B(_0390_),
    .C(_0395_),
    .A(_0384_),
    .Y(_0397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2895_ (.B1(_0382_),
    .VDD(VPWR),
    .Y(_0398_),
    .VSS(VGND),
    .A1(net789),
    .A2(_0335_));
 sg13g2_nor4_1 _2896_ (.A(_0377_),
    .B(_0396_),
    .C(_0397_),
    .D(_0398_),
    .Y(_0399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2897_ (.B(_0391_),
    .C(_0392_),
    .A(_0383_),
    .Y(_0400_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0399_));
 sg13g2_a21o_1 _2898_ (.A2(_0400_),
    .A1(_0372_),
    .B1(net694),
    .X(_0401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2899_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2051_),
    .A2(net694),
    .Y(_0402_),
    .B1(net599));
 sg13g2_a22oi_1 _2900_ (.Y(_0403_),
    .B1(_0401_),
    .B2(_0402_),
    .A2(net599),
    .A1(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2901_ (.VDD(VPWR),
    .Y(_0034_),
    .A(_0403_),
    .VSS(VGND));
 sg13g2_nand3_1 _2902_ (.B(\sap_3_inst.alu_inst.tmp[2] ),
    .C(_0363_),
    .A(net786),
    .Y(_0404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2903_ (.Y(_0405_),
    .A(net786),
    .B(\sap_3_inst.alu_inst.tmp[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2904_ (.B1(_0404_),
    .VDD(VPWR),
    .Y(_0406_),
    .VSS(VGND),
    .A1(_0355_),
    .A2(_0405_));
 sg13g2_o21ai_1 _2905_ (.B1(_0361_),
    .VDD(VPWR),
    .Y(_0407_),
    .VSS(VGND),
    .A1(net787),
    .A2(\sap_3_inst.alu_inst.tmp[2] ));
 sg13g2_o21ai_1 _2906_ (.B1(_0407_),
    .VDD(VPWR),
    .Y(_0408_),
    .VSS(VGND),
    .A1(net786),
    .A2(_0334_));
 sg13g2_nor2_1 _2907_ (.A(_0406_),
    .B(_0408_),
    .Y(_0409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2908_ (.Y(_0410_),
    .B(net790),
    .A_N(\sap_3_inst.alu_inst.tmp[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2909_ (.B1(_0410_),
    .VDD(VPWR),
    .Y(_0411_),
    .VSS(VGND),
    .A1(_0374_),
    .A2(_0378_));
 sg13g2_xor2_1 _2910_ (.B(_0411_),
    .A(_0405_),
    .X(_0412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2911_ (.A(_0380_),
    .B(_0405_),
    .X(_0413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2912_ (.Y(_0414_),
    .A(_0348_),
    .B(_0413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2913_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0373_),
    .A2(_0375_),
    .Y(_0415_),
    .B1(_0405_));
 sg13g2_nand3_1 _2914_ (.B(_0375_),
    .C(_0405_),
    .A(_0373_),
    .Y(_0416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2915_ (.A(_0415_),
    .B_N(_0416_),
    .Y(_0417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2916_ (.A(_0393_),
    .B_N(_0417_),
    .Y(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2917_ (.VDD(VPWR),
    .Y(_0419_),
    .A(_0418_),
    .VSS(VGND));
 sg13g2_xnor2_1 _2918_ (.Y(_0420_),
    .A(_0393_),
    .B(_0417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2919_ (.Y(_0421_),
    .B1(_0420_),
    .B2(_0344_),
    .A2(_0413_),
    .A1(_0348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2920_ (.Y(_0422_),
    .A(net786),
    .B(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2921_ (.Y(_0423_),
    .A(net786),
    .B(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2922_ (.B(_0387_),
    .C(_0423_),
    .A(_0385_),
    .Y(_0424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2923_ (.A2(_0387_),
    .A1(_0385_),
    .B1(_0423_),
    .X(_0425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2924_ (.X(_0426_),
    .A(net704),
    .B(_0424_),
    .C(_0425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2925_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net783),
    .C1(_0426_),
    .B1(net691),
    .A1(net789),
    .Y(_0427_),
    .A2(net692));
 sg13g2_o21ai_1 _2926_ (.B1(_0346_),
    .VDD(VPWR),
    .Y(_0428_),
    .VSS(VGND),
    .A1(_0349_),
    .A2(_0380_));
 sg13g2_nand4_1 _2927_ (.B(_0409_),
    .C(_0421_),
    .A(net575),
    .Y(_0429_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0427_));
 sg13g2_a21oi_1 _2928_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0412_),
    .A2(_0428_),
    .Y(_0430_),
    .B1(_0429_));
 sg13g2_nor2_1 _2929_ (.A(net575),
    .B(_0417_),
    .Y(_0431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2930_ (.A(net702),
    .B(_0430_),
    .C(_0431_),
    .Y(_0432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2931_ (.Y(_0433_),
    .A(\sap_3_inst.alu_inst.act[2] ),
    .B(net702),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2932_ (.A(net693),
    .B(_0432_),
    .Y(_0434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2933_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0434_),
    .C1(net598),
    .B1(_0433_),
    .A1(_0227_),
    .Y(_0435_),
    .A2(net693));
 sg13g2_a21o_1 _2934_ (.A2(net598),
    .A1(net787),
    .B1(_0435_),
    .X(_0035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2935_ (.A(net32),
    .B_N(net693),
    .Y(_0436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2936_ (.A(net784),
    .B(\sap_3_inst.alu_inst.tmp[3] ),
    .Y(_0437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2937_ (.Y(_0438_),
    .A(net784),
    .B(\sap_3_inst.alu_inst.tmp[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2938_ (.Y(_0439_),
    .B(_0438_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0437_));
 sg13g2_inv_1 _2939_ (.VDD(VPWR),
    .Y(_0440_),
    .A(_0439_),
    .VSS(VGND));
 sg13g2_nor2b_1 _2940_ (.A(\sap_3_inst.alu_inst.tmp[2] ),
    .B_N(net787),
    .Y(_0441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2941_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0405_),
    .A2(_0411_),
    .Y(_0442_),
    .B1(_0441_));
 sg13g2_nor2_1 _2942_ (.A(_0440_),
    .B(_0442_),
    .Y(_0443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2943_ (.Y(_0444_),
    .A(_0439_),
    .B(_0442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2944_ (.A(_0414_),
    .B(_0444_),
    .Y(_0445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2945_ (.B(\sap_3_inst.alu_inst.tmp[3] ),
    .C(_0363_),
    .A(net784),
    .Y(_0446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2946_ (.B1(_0446_),
    .VDD(VPWR),
    .Y(_0447_),
    .VSS(VGND),
    .A1(_0355_),
    .A2(_0439_));
 sg13g2_nand2b_1 _2947_ (.Y(_0448_),
    .B(_0361_),
    .A_N(_0437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2948_ (.Y(_0449_),
    .B1(net691),
    .B2(net781),
    .A2(net692),
    .A1(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2949_ (.Y(_0450_),
    .A(_0448_),
    .B(_0449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2950_ (.A(_0445_),
    .B(_0447_),
    .C(_0450_),
    .Y(_0451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2951_ (.B1(_0346_),
    .VDD(VPWR),
    .Y(_0452_),
    .VSS(VGND),
    .A1(_0349_),
    .A2(_0413_));
 sg13g2_nand2_1 _2952_ (.Y(_0453_),
    .A(_0422_),
    .B(_0425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2953_ (.Y(_0454_),
    .A(net783),
    .B(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2954_ (.Y(_0455_),
    .A(net783),
    .B(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2955_ (.Y(_0456_),
    .A(_0453_),
    .B(_0455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2956_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net787),
    .A2(\sap_3_inst.alu_inst.tmp[2] ),
    .Y(_0457_),
    .B1(_0415_));
 sg13g2_xnor2_1 _2957_ (.Y(_0458_),
    .A(_0439_),
    .B(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2958_ (.A(_0419_),
    .B(_0458_),
    .Y(_0459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2959_ (.Y(_0460_),
    .A(_0418_),
    .B(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2960_ (.Y(_0461_),
    .B1(_0460_),
    .B2(_0344_),
    .A2(_0456_),
    .A1(net704),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2961_ (.B1(_0461_),
    .VDD(VPWR),
    .Y(_0462_),
    .VSS(VGND),
    .A1(net783),
    .A2(_0334_));
 sg13g2_a21oi_1 _2962_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0444_),
    .A2(_0452_),
    .Y(_0463_),
    .B1(_0462_));
 sg13g2_nand3_1 _2963_ (.B(_0451_),
    .C(_0463_),
    .A(net575),
    .Y(_0464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2964_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0353_),
    .A2(_0458_),
    .Y(_0465_),
    .B1(net702));
 sg13g2_a221oi_1 _2965_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0465_),
    .C1(net693),
    .B1(_0464_),
    .A1(\sap_3_inst.alu_inst.act[3] ),
    .Y(_0466_),
    .A2(_0320_));
 sg13g2_nor3_1 _2966_ (.A(net598),
    .B(_0436_),
    .C(_0466_),
    .Y(_0467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2967_ (.A2(net598),
    .A1(net783),
    .B1(_0467_),
    .X(_0036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2968_ (.Y(_0468_),
    .A(net781),
    .B(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2969_ (.B1(_0453_),
    .VDD(VPWR),
    .Y(_0469_),
    .VSS(VGND),
    .A1(net783),
    .A2(net708));
 sg13g2_nand3_1 _2970_ (.B(_0468_),
    .C(_0469_),
    .A(_0454_),
    .Y(_0470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2971_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0454_),
    .A2(_0469_),
    .Y(_0471_),
    .B1(_0468_));
 sg13g2_nand2_1 _2972_ (.Y(_0472_),
    .A(net704),
    .B(_0470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2973_ (.A(net782),
    .B(\sap_3_inst.alu_inst.tmp[4] ),
    .X(_0473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2974_ (.Y(_0474_),
    .A(net781),
    .B(\sap_3_inst.alu_inst.tmp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2975_ (.VDD(VPWR),
    .Y(_0475_),
    .A(_0474_),
    .VSS(VGND));
 sg13g2_nor2b_1 _2976_ (.A(\sap_3_inst.alu_inst.tmp[3] ),
    .B_N(net784),
    .Y(_0476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2977_ (.B1(_0474_),
    .VDD(VPWR),
    .Y(_0477_),
    .VSS(VGND),
    .A1(_0443_),
    .A2(_0476_));
 sg13g2_or3_1 _2978_ (.A(_0443_),
    .B(_0474_),
    .C(_0476_),
    .X(_0478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2979_ (.A(_0477_),
    .B(_0478_),
    .X(_0479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2980_ (.VDD(VPWR),
    .Y(_0480_),
    .A(_0479_),
    .VSS(VGND));
 sg13g2_nand2_2 _2981_ (.Y(_0481_),
    .A(_0413_),
    .B(_0439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2982_ (.B(_0481_),
    .A(_0479_),
    .X(_0482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2983_ (.B1(_0361_),
    .VDD(VPWR),
    .Y(_0483_),
    .VSS(VGND),
    .A1(net782),
    .A2(\sap_3_inst.alu_inst.tmp[4] ));
 sg13g2_o21ai_1 _2984_ (.B1(_0483_),
    .VDD(VPWR),
    .Y(_0484_),
    .VSS(VGND),
    .A1(_0349_),
    .A2(_0482_));
 sg13g2_nand2_1 _2985_ (.Y(_0485_),
    .A(_0363_),
    .B(_0473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2986_ (.B1(_0485_),
    .VDD(VPWR),
    .Y(_0486_),
    .VSS(VGND),
    .A1(_0346_),
    .A2(_0480_));
 sg13g2_a22oi_1 _2987_ (.Y(_0487_),
    .B1(net691),
    .B2(net778),
    .A2(net692),
    .A1(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2988_ (.B1(_0487_),
    .VDD(VPWR),
    .Y(_0488_),
    .VSS(VGND),
    .A1(net781),
    .A2(_0334_));
 sg13g2_a21oi_1 _2989_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0438_),
    .A2(_0457_),
    .Y(_0489_),
    .B1(_0437_));
 sg13g2_xnor2_1 _2990_ (.Y(_0490_),
    .A(_0474_),
    .B(_0489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2991_ (.Y(_0491_),
    .A(_0459_),
    .B(_0490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2992_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0492_),
    .B(_0490_),
    .A(_0459_));
 sg13g2_nand3_1 _2993_ (.B(_0491_),
    .C(_0492_),
    .A(_0344_),
    .Y(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2994_ (.B1(_0493_),
    .VDD(VPWR),
    .Y(_0494_),
    .VSS(VGND),
    .A1(_0355_),
    .A2(_0474_));
 sg13g2_nor4_1 _2995_ (.A(_0484_),
    .B(_0486_),
    .C(_0488_),
    .D(_0494_),
    .Y(_0495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2996_ (.B1(_0495_),
    .VDD(VPWR),
    .Y(_0496_),
    .VSS(VGND),
    .A1(_0471_),
    .A2(_0472_));
 sg13g2_mux2_1 _2997_ (.A0(_0490_),
    .A1(_0496_),
    .S(net575),
    .X(_0497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2998_ (.Y(_0498_),
    .B(_0497_),
    .A_N(net702),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2999_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu_inst.act[4] ),
    .A2(net702),
    .Y(_0499_),
    .B1(net693));
 sg13g2_a221oi_1 _3000_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0499_),
    .C1(net599),
    .B1(_0498_),
    .A1(_1991_),
    .Y(_0500_),
    .A2(_0330_));
 sg13g2_a21o_1 _3001_ (.A2(_0340_),
    .A1(net781),
    .B1(_0500_),
    .X(_0037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3002_ (.A2(net708),
    .A1(net782),
    .B1(_0471_),
    .X(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3003_ (.Y(_0502_),
    .A(net778),
    .B(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3004_ (.B(net709),
    .A(net778),
    .X(_0503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3005_ (.B1(net704),
    .VDD(VPWR),
    .Y(_0504_),
    .VSS(VGND),
    .A1(_0501_),
    .A2(_0503_));
 sg13g2_a21oi_1 _3006_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0501_),
    .A2(_0503_),
    .Y(_0505_),
    .B1(_0504_));
 sg13g2_nor2_1 _3007_ (.A(net778),
    .B(\sap_3_inst.alu_inst.tmp[5] ),
    .Y(_0506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3008_ (.Y(_0507_),
    .A(net778),
    .B(\sap_3_inst.alu_inst.tmp[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3009_ (.A(_0506_),
    .B_N(_0507_),
    .Y(_0508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3010_ (.A(_0355_),
    .B_N(_0507_),
    .Y(_0509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3011_ (.A(_0361_),
    .B(_0509_),
    .Y(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3012_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0511_),
    .B(_0510_),
    .A(_0506_));
 sg13g2_nand2b_1 _3013_ (.Y(_0512_),
    .B(net781),
    .A_N(\sap_3_inst.alu_inst.tmp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3014_ (.A(_0477_),
    .B(_0512_),
    .X(_0513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3015_ (.A(_0508_),
    .B(_0513_),
    .Y(_0514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3016_ (.B(_0513_),
    .A(_0508_),
    .X(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3017_ (.A(net780),
    .B(_0336_),
    .Y(_0516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3018_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0347_),
    .A2(_0515_),
    .Y(_0517_),
    .B1(_0516_));
 sg13g2_a21oi_1 _3019_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0475_),
    .A2(_0489_),
    .Y(_0518_),
    .B1(_0473_));
 sg13g2_xor2_1 _3020_ (.B(_0518_),
    .A(_0508_),
    .X(_0519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3021_ (.A(_0491_),
    .B(_0519_),
    .Y(_0520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3022_ (.B(_0519_),
    .A(_0491_),
    .X(_0521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3023_ (.A(_0475_),
    .B(_0481_),
    .C(_0508_),
    .Y(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3024_ (.B1(_0515_),
    .VDD(VPWR),
    .Y(_0523_),
    .VSS(VGND),
    .A1(_0479_),
    .A2(_0481_));
 sg13g2_nand2b_1 _3025_ (.Y(_0524_),
    .B(_0523_),
    .A_N(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3026_ (.B(\sap_3_inst.alu_inst.tmp[5] ),
    .C(_0363_),
    .A(net778),
    .Y(_0525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3027_ (.Y(_0526_),
    .B1(_0359_),
    .B2(net775),
    .A2(net692),
    .A1(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3028_ (.Y(_0527_),
    .A(_0525_),
    .B(_0526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3029_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0348_),
    .C1(_0527_),
    .B1(_0524_),
    .A1(_0344_),
    .Y(_0528_),
    .A2(_0521_));
 sg13g2_nand4_1 _3030_ (.B(_0511_),
    .C(_0517_),
    .A(_0354_),
    .Y(_0529_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0528_));
 sg13g2_a21oi_1 _3031_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0353_),
    .A2(_0519_),
    .Y(_0530_),
    .B1(net702));
 sg13g2_o21ai_1 _3032_ (.B1(_0530_),
    .VDD(VPWR),
    .Y(_0531_),
    .VSS(VGND),
    .A1(_0505_),
    .A2(_0529_));
 sg13g2_a21oi_1 _3033_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu_inst.act[5] ),
    .A2(_0320_),
    .Y(_0532_),
    .B1(net693));
 sg13g2_a221oi_1 _3034_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0532_),
    .C1(net598),
    .B1(_0531_),
    .A1(net569),
    .Y(_0533_),
    .A2(_0330_));
 sg13g2_a21o_1 _3035_ (.A2(net598),
    .A1(net779),
    .B1(_0533_),
    .X(_0038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3036_ (.Y(_0534_),
    .A(net775),
    .B(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3037_ (.Y(_0535_),
    .A(net775),
    .B(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3038_ (.B1(_0501_),
    .VDD(VPWR),
    .Y(_0536_),
    .VSS(VGND),
    .A1(net778),
    .A2(net709));
 sg13g2_a21o_1 _3039_ (.A2(_0536_),
    .A1(_0502_),
    .B1(_0535_),
    .X(_0537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3040_ (.B(_0535_),
    .C(_0536_),
    .A(_0502_),
    .Y(_0538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3041_ (.B(_0537_),
    .C(_0538_),
    .A(net704),
    .Y(_0539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3042_ (.A(net775),
    .B(\sap_3_inst.alu_inst.tmp[6] ),
    .X(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3043_ (.Y(_0541_),
    .A(_0363_),
    .B(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3044_ (.B(\sap_3_inst.alu_inst.tmp[6] ),
    .A(net775),
    .X(_0542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3045_ (.B(_0333_),
    .C(_0542_),
    .A(_2012_),
    .Y(_0543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3046_ (.B1(_0361_),
    .VDD(VPWR),
    .Y(_0544_),
    .VSS(VGND),
    .A1(net776),
    .A2(\sap_3_inst.alu_inst.tmp[6] ));
 sg13g2_a21oi_1 _3047_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net778),
    .A2(_1527_),
    .Y(_0545_),
    .B1(_0514_));
 sg13g2_nor2_1 _3048_ (.A(_0542_),
    .B(_0545_),
    .Y(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3049_ (.B(_0545_),
    .A(_0542_),
    .X(_0547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3050_ (.Y(_0548_),
    .B1(net691),
    .B2(net772),
    .A2(_0357_),
    .A1(net780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3051_ (.B1(_0548_),
    .VDD(VPWR),
    .Y(_0549_),
    .VSS(VGND),
    .A1(net775),
    .A2(_0334_));
 sg13g2_a21oi_1 _3052_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0347_),
    .A2(_0547_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_nand4_1 _3053_ (.B(_0543_),
    .C(_0544_),
    .A(_0541_),
    .Y(_0551_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0550_));
 sg13g2_nor2b_1 _3054_ (.A(_0547_),
    .B_N(_0522_),
    .Y(_0552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3055_ (.Y(_0553_),
    .A(_0522_),
    .B(_0547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3056_ (.B1(_0507_),
    .VDD(VPWR),
    .Y(_0554_),
    .VSS(VGND),
    .A1(_0506_),
    .A2(_0518_));
 sg13g2_xor2_1 _3057_ (.B(_0554_),
    .A(_0542_),
    .X(_0555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3058_ (.Y(_0556_),
    .A(_0542_),
    .B(_0554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3059_ (.Y(_0557_),
    .A(_0520_),
    .B(_0555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3060_ (.B1(_0344_),
    .VDD(VPWR),
    .Y(_0558_),
    .VSS(VGND),
    .A1(_0520_),
    .A2(_0555_));
 sg13g2_nand2b_1 _3061_ (.Y(_0559_),
    .B(_0557_),
    .A_N(_0558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3062_ (.B1(_0559_),
    .VDD(VPWR),
    .Y(_0560_),
    .VSS(VGND),
    .A1(_0349_),
    .A2(_0553_));
 sg13g2_nor3_1 _3063_ (.A(_0353_),
    .B(_0551_),
    .C(_0560_),
    .Y(_0561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3064_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0539_),
    .C1(net702),
    .B1(_0561_),
    .A1(_0353_),
    .Y(_0562_),
    .A2(_0556_));
 sg13g2_a21oi_1 _3065_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu_inst.act[6] ),
    .A2(net702),
    .Y(_0563_),
    .B1(net693));
 sg13g2_nand2b_1 _3066_ (.Y(_0564_),
    .B(_0563_),
    .A_N(_0562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3067_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1941_),
    .A2(net693),
    .Y(_0565_),
    .B1(net598));
 sg13g2_a22oi_1 _3068_ (.Y(_0566_),
    .B1(_0564_),
    .B2(_0565_),
    .A2(net598),
    .A1(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3069_ (.VDD(VPWR),
    .Y(_0039_),
    .A(_0566_),
    .VSS(VGND));
 sg13g2_nand2_1 _3070_ (.Y(_0567_),
    .A(_0534_),
    .B(_0537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3071_ (.Y(_0568_),
    .A(net772),
    .B(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3072_ (.Y(_0569_),
    .A(_0567_),
    .B(_0568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3073_ (.A(net772),
    .B(\sap_3_inst.alu_inst.tmp[7] ),
    .Y(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3074_ (.Y(_0571_),
    .A(net772),
    .B(\sap_3_inst.alu_inst.tmp[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3075_ (.Y(_0572_),
    .B(_0571_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0570_));
 sg13g2_inv_1 _3076_ (.VDD(VPWR),
    .Y(_0573_),
    .A(_0572_),
    .VSS(VGND));
 sg13g2_a21oi_1 _3077_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0542_),
    .A2(_0554_),
    .Y(_0574_),
    .B1(_0540_));
 sg13g2_xnor2_1 _3078_ (.Y(_0575_),
    .A(_0573_),
    .B(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3079_ (.Y(_0576_),
    .A(_0557_),
    .B(_0575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3080_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net775),
    .A2(_1528_),
    .Y(_0577_),
    .B1(_0546_));
 sg13g2_xnor2_1 _3081_ (.Y(_0578_),
    .A(_0572_),
    .B(_0577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3082_ (.B(\sap_3_inst.alu_inst.tmp[7] ),
    .C(_0363_),
    .A(net772),
    .Y(_0579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3083_ (.Y(_0580_),
    .B1(_0358_),
    .B2(net691),
    .A2(net692),
    .A1(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3084_ (.Y(_0581_),
    .B(_0361_),
    .A_N(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3085_ (.A(_0355_),
    .B(_0572_),
    .Y(_0582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3086_ (.A(net772),
    .B(_0334_),
    .Y(_0583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3087_ (.A(_0582_),
    .B(_0583_),
    .Y(_0584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3088_ (.A(_0579_),
    .B(_0580_),
    .C(_0581_),
    .D(_0584_),
    .X(_0585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3089_ (.A(_0542_),
    .B(_0573_),
    .Y(_0586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3090_ (.B(_0522_),
    .C(_0586_),
    .A(_0348_),
    .Y(_0587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3091_ (.B1(_0346_),
    .VDD(VPWR),
    .Y(_0588_),
    .VSS(VGND),
    .A1(_0349_),
    .A2(_0552_));
 sg13g2_a22oi_1 _3092_ (.Y(_0589_),
    .B1(_0578_),
    .B2(_0588_),
    .A2(_0576_),
    .A1(_0344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3093_ (.B(_0585_),
    .C(_0587_),
    .A(net575),
    .Y(_0590_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0589_));
 sg13g2_a21oi_1 _3094_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2000_),
    .A2(_0569_),
    .Y(_0591_),
    .B1(_0590_));
 sg13g2_nor2_1 _3095_ (.A(net703),
    .B(_0591_),
    .Y(_0592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3096_ (.B1(_0592_),
    .VDD(VPWR),
    .Y(_0593_),
    .VSS(VGND),
    .A1(net575),
    .A2(_0575_));
 sg13g2_a21oi_1 _3097_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu_inst.act[7] ),
    .A2(net703),
    .Y(_0594_),
    .B1(net694));
 sg13g2_a221oi_1 _3098_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0594_),
    .C1(net599),
    .B1(_0593_),
    .A1(_1914_),
    .Y(_0595_),
    .A2(net694));
 sg13g2_a21o_1 _3099_ (.A2(net599),
    .A1(net773),
    .B1(_0595_),
    .X(_0040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3100_ (.Y(_0596_),
    .A(\sap_3_inst.out[0] ),
    .B(net705),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3101_ (.B1(_0596_),
    .VDD(VPWR),
    .Y(_0041_),
    .VSS(VGND),
    .A1(_1508_),
    .A2(net705));
 sg13g2_mux2_1 _3102_ (.A0(net789),
    .A1(\sap_3_inst.out[1] ),
    .S(net705),
    .X(_0042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3103_ (.A0(net786),
    .A1(\sap_3_inst.out[2] ),
    .S(net705),
    .X(_0043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3104_ (.A0(net783),
    .A1(\sap_3_inst.out[3] ),
    .S(net705),
    .X(_0044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3105_ (.Y(_0597_),
    .A(\sap_3_inst.out[4] ),
    .B(net706),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3106_ (.B1(_0597_),
    .VDD(VPWR),
    .Y(_0045_),
    .VSS(VGND),
    .A1(_1509_),
    .A2(net706));
 sg13g2_mux2_1 _3107_ (.A0(net779),
    .A1(\sap_3_inst.out[5] ),
    .S(net706),
    .X(_0046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3108_ (.A0(net775),
    .A1(\sap_3_inst.out[6] ),
    .S(net706),
    .X(_0047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3109_ (.A0(net774),
    .A1(\sap_3_inst.out[7] ),
    .S(net706),
    .X(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3110_ (.Y(_0598_),
    .A(net772),
    .B(_1529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3111_ (.B1(_0587_),
    .VDD(VPWR),
    .Y(_0599_),
    .VSS(VGND),
    .A1(net773),
    .A2(_1529_));
 sg13g2_a21o_1 _3112_ (.A2(_0598_),
    .A1(_0577_),
    .B1(_0599_),
    .X(_0600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3113_ (.A(_0475_),
    .B(_0508_),
    .X(_0601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3114_ (.B(_0542_),
    .C(_0573_),
    .A(_0459_),
    .Y(_0602_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0601_));
 sg13g2_nand3_1 _3115_ (.B(_2004_),
    .C(_2006_),
    .A(net761),
    .Y(_0603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3116_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.alu_flags[1] ),
    .A2(_2017_),
    .Y(_0604_),
    .B1(_0603_));
 sg13g2_a221oi_1 _3117_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net792),
    .C1(_0604_),
    .B1(net691),
    .A1(net772),
    .Y(_0605_),
    .A2(net692));
 sg13g2_o21ai_1 _3118_ (.B1(_0605_),
    .VDD(VPWR),
    .Y(_0606_),
    .VSS(VGND),
    .A1(_0345_),
    .A2(_0602_));
 sg13g2_a21oi_1 _3119_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0350_),
    .A2(_0600_),
    .Y(_0607_),
    .B1(_0606_));
 sg13g2_nor2_1 _3120_ (.A(_2002_),
    .B(_2023_),
    .Y(_0608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3121_ (.Y(_0609_),
    .A(_2022_),
    .B(_0351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3122_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0345_),
    .C1(_0570_),
    .B1(_0609_),
    .A1(_0571_),
    .Y(_0610_),
    .A2(_0574_));
 sg13g2_nor2b_1 _3123_ (.A(_0610_),
    .B_N(_0608_),
    .Y(_0611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3124_ (.A(\sap_3_inst.alu_inst.carry ),
    .B(_0608_),
    .Y(_0612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3125_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0607_),
    .A2(_0611_),
    .Y(_0049_),
    .B1(_0612_));
 sg13g2_a21oi_1 _3126_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net730),
    .A2(_1595_),
    .Y(_0613_),
    .B1(_1874_));
 sg13g2_nand2_1 _3127_ (.Y(_0614_),
    .A(net716),
    .B(_0613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3128_ (.B1(_1880_),
    .VDD(VPWR),
    .Y(_0615_),
    .VSS(VGND),
    .A1(_1800_),
    .A2(_0614_));
 sg13g2_mux2_1 _3129_ (.A0(net17),
    .A1(\sap_3_inst.alu_inst.tmp[0] ),
    .S(net701),
    .X(_0050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3130_ (.Y(_0616_),
    .A(\sap_3_inst.alu_inst.tmp[1] ),
    .B(net700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3131_ (.B1(_0616_),
    .VDD(VPWR),
    .Y(_0051_),
    .VSS(VGND),
    .A1(_2051_),
    .A2(net701));
 sg13g2_nand2_1 _3132_ (.Y(_0617_),
    .A(\sap_3_inst.alu_inst.tmp[2] ),
    .B(net700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3133_ (.B1(_0617_),
    .VDD(VPWR),
    .Y(_0052_),
    .VSS(VGND),
    .A1(_0227_),
    .A2(net700));
 sg13g2_mux2_1 _3134_ (.A0(net32),
    .A1(\sap_3_inst.alu_inst.tmp[3] ),
    .S(net700),
    .X(_0053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3135_ (.Y(_0618_),
    .A(\sap_3_inst.alu_inst.tmp[4] ),
    .B(net700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3136_ (.B1(_0618_),
    .VDD(VPWR),
    .Y(_0054_),
    .VSS(VGND),
    .A1(_1991_),
    .A2(net701));
 sg13g2_nand2_1 _3137_ (.Y(_0619_),
    .A(\sap_3_inst.alu_inst.tmp[5] ),
    .B(net700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3138_ (.B1(_0619_),
    .VDD(VPWR),
    .Y(_0055_),
    .VSS(VGND),
    .A1(_1967_),
    .A2(net701));
 sg13g2_nand2_1 _3139_ (.Y(_0620_),
    .A(\sap_3_inst.alu_inst.tmp[6] ),
    .B(net700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3140_ (.B1(_0620_),
    .VDD(VPWR),
    .Y(_0056_),
    .VSS(VGND),
    .A1(net570),
    .A2(net700));
 sg13g2_nor2_1 _3141_ (.A(net24),
    .B(net701),
    .Y(_0621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3142_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1529_),
    .A2(net701),
    .Y(_0057_),
    .B1(_0621_));
 sg13g2_mux2_1 _3143_ (.A0(\sap_3_inst.controller_inst.opcode[0] ),
    .A1(net31),
    .S(net717),
    .X(_0058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3144_ (.A(net769),
    .B(net718),
    .Y(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3145_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net717),
    .A2(_2051_),
    .Y(_0059_),
    .B1(_0622_));
 sg13g2_nand2_1 _3146_ (.Y(_0623_),
    .A(net718),
    .B(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3147_ (.B1(_0623_),
    .VDD(VPWR),
    .Y(_0060_),
    .VSS(VGND),
    .A1(_1494_),
    .A2(_1585_));
 sg13g2_nand2_1 _3148_ (.Y(_0624_),
    .A(net717),
    .B(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3149_ (.B1(_0624_),
    .VDD(VPWR),
    .Y(_0061_),
    .VSS(VGND),
    .A1(_1493_),
    .A2(net717));
 sg13g2_nor2_1 _3150_ (.A(net759),
    .B(net717),
    .Y(_0625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3151_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net717),
    .A2(_1991_),
    .Y(_0062_),
    .B1(_0625_));
 sg13g2_nor2_1 _3152_ (.A(net758),
    .B(net717),
    .Y(_0626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3153_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net717),
    .A2(net569),
    .Y(_0063_),
    .B1(_0626_));
 sg13g2_nor2_1 _3154_ (.A(net756),
    .B(net718),
    .Y(_0627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3155_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net718),
    .A2(_1941_),
    .Y(_0064_),
    .B1(_0627_));
 sg13g2_nor2_1 _3156_ (.A(net754),
    .B(net718),
    .Y(_0628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3157_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1585_),
    .A2(_1914_),
    .Y(_0065_),
    .B1(_0628_));
 sg13g2_nand3_1 _3158_ (.B(_1633_),
    .C(_1667_),
    .A(_1627_),
    .Y(_0629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3159_ (.Y(_0630_),
    .B(_1627_),
    .A_N(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3160_ (.Y(_0631_),
    .B(_1635_),
    .A_N(net724),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3161_ (.B(_0630_),
    .C(_0631_),
    .A(_0629_),
    .Y(_0632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3162_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1634_),
    .A2(_1709_),
    .Y(_0633_),
    .B1(_1653_));
 sg13g2_a22oi_1 _3163_ (.Y(_0634_),
    .B1(net720),
    .B2(_1634_),
    .A2(_1666_),
    .A1(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3164_ (.Y(_0635_),
    .A(_1762_),
    .B(_1875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3165_ (.B(_1645_),
    .C(_1692_),
    .A(net761),
    .Y(_0636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3166_ (.Y(_0637_),
    .B1(_0636_),
    .B2(_1634_),
    .A2(_1776_),
    .A1(_1646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3167_ (.B1(_1659_),
    .VDD(VPWR),
    .Y(_0638_),
    .VSS(VGND),
    .A1(_1633_),
    .A2(_1705_));
 sg13g2_a22oi_1 _3168_ (.Y(_0639_),
    .B1(_1822_),
    .B2(_1875_),
    .A2(_1699_),
    .A1(_1633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3169_ (.B(_1889_),
    .C(_0638_),
    .A(_1816_),
    .Y(_0640_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0639_));
 sg13g2_nor4_1 _3170_ (.A(_0633_),
    .B(_0634_),
    .C(_0637_),
    .D(_0640_),
    .Y(_0641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3171_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net715),
    .C1(net719),
    .B1(_0632_),
    .A1(net759),
    .Y(_0642_),
    .A2(_1886_));
 sg13g2_nor3_1 _3172_ (.A(net750),
    .B(net728),
    .C(_1761_),
    .Y(_0643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3173_ (.A(_1573_),
    .B(net729),
    .C(_1616_),
    .Y(_0644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3174_ (.B1(net759),
    .VDD(VPWR),
    .Y(_0645_),
    .VSS(VGND),
    .A1(_0643_),
    .A2(_0644_));
 sg13g2_a21o_1 _3175_ (.A2(_0645_),
    .A1(net719),
    .B1(net739),
    .X(_0646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3176_ (.A2(_0642_),
    .A1(_0641_),
    .B1(_0646_),
    .X(_0647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3177_ (.Y(_0648_),
    .A(net740),
    .B(_0647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3178_ (.Y(_0649_),
    .A(net741),
    .B(_1823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3179_ (.B(_1869_),
    .C(_0649_),
    .A(_1555_),
    .Y(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3180_ (.VDD(VPWR),
    .Y(_0651_),
    .A(_0650_),
    .VSS(VGND));
 sg13g2_a21oi_2 _3181_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0650_),
    .Y(_0652_),
    .A2(_0647_),
    .A1(net740));
 sg13g2_a21o_2 _3182_ (.A2(_0647_),
    .A1(_1567_),
    .B1(_0650_),
    .X(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3183_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net752),
    .A2(_1627_),
    .Y(_0654_),
    .B1(_1777_));
 sg13g2_a21oi_1 _3184_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1658_),
    .A2(_0654_),
    .Y(_0655_),
    .B1(net721));
 sg13g2_nand2_1 _3185_ (.Y(_0656_),
    .A(_1731_),
    .B(_1782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3186_ (.A(net750),
    .B(net727),
    .C(_1837_),
    .Y(_0657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3187_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net764),
    .C1(_0657_),
    .B1(_1886_),
    .A1(_1629_),
    .Y(_0658_),
    .A2(net734));
 sg13g2_nor4_1 _3188_ (.A(_1491_),
    .B(net746),
    .C(_1493_),
    .D(_1680_),
    .Y(_0659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3189_ (.B1(_1659_),
    .VDD(VPWR),
    .Y(_0660_),
    .VSS(VGND),
    .A1(net722),
    .A2(_0659_));
 sg13g2_nand3_1 _3190_ (.B(_0658_),
    .C(_0660_),
    .A(_0656_),
    .Y(_0661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3191_ (.B1(net740),
    .VDD(VPWR),
    .Y(_0662_),
    .VSS(VGND),
    .A1(_0655_),
    .A2(_0661_));
 sg13g2_or4_1 _3192_ (.A(net754),
    .B(_1563_),
    .C(net721),
    .D(_1837_),
    .X(_0663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3193_ (.A(_0662_),
    .B(_0663_),
    .X(_0664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3194_ (.Y(_0665_),
    .A(_0662_),
    .B(_0663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3195_ (.A(_0652_),
    .B(_0665_),
    .Y(_0666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3196_ (.Y(_0667_),
    .A(_0653_),
    .B(_0664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3197_ (.Y(_0668_),
    .A(net705),
    .B(_0630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3198_ (.A(net714),
    .B(net705),
    .C(_0630_),
    .D(_0631_),
    .X(_0669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3199_ (.Y(_0670_),
    .A(_1649_),
    .B(_1670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3200_ (.Y(_0671_),
    .A(_1587_),
    .B(_1679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3201_ (.Y(_0672_),
    .A(_1673_),
    .B(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3202_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0673_),
    .B(_0671_),
    .A(net735));
 sg13g2_nand4_1 _3203_ (.B(_1673_),
    .C(net720),
    .A(net726),
    .Y(_0674_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0671_));
 sg13g2_nand3_1 _3204_ (.B(_1670_),
    .C(_0674_),
    .A(_1649_),
    .Y(_0675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3205_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net727),
    .A2(net720),
    .Y(_0676_),
    .B1(_1691_));
 sg13g2_nand3_1 _3206_ (.B(_1652_),
    .C(_1666_),
    .A(_1644_),
    .Y(_0677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3207_ (.Y(_0678_),
    .B1(_0677_),
    .B2(_0672_),
    .A2(_0676_),
    .A1(_1670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3208_ (.X(_0679_),
    .A(_0673_),
    .B(_0675_),
    .C(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3209_ (.A(_1639_),
    .B(_1699_),
    .Y(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3210_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0279_),
    .A2(_0680_),
    .Y(_0681_),
    .B1(_1752_));
 sg13g2_nor2_1 _3211_ (.A(net715),
    .B(_0681_),
    .Y(_0682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3212_ (.A(_1495_),
    .B(_0636_),
    .Y(_0683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3213_ (.B1(_1645_),
    .VDD(VPWR),
    .Y(_0684_),
    .VSS(VGND),
    .A1(_1612_),
    .A2(_1672_));
 sg13g2_o21ai_1 _3214_ (.B1(_0684_),
    .VDD(VPWR),
    .Y(_0685_),
    .VSS(VGND),
    .A1(_1660_),
    .A2(_1752_));
 sg13g2_nor4_1 _3215_ (.A(net714),
    .B(_0681_),
    .C(_0683_),
    .D(_0685_),
    .Y(_0686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3216_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0679_),
    .A2(_0686_),
    .Y(_0687_),
    .B1(_0669_));
 sg13g2_o21ai_1 _3217_ (.B1(_0288_),
    .VDD(VPWR),
    .Y(_0688_),
    .VSS(VGND),
    .A1(_1621_),
    .A2(_0687_));
 sg13g2_a22oi_1 _3218_ (.Y(_0689_),
    .B1(_0644_),
    .B2(_1557_),
    .A2(net737),
    .A1(net743),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3219_ (.Y(_0690_),
    .A(_0688_),
    .B(_0689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3220_ (.A(_1699_),
    .B(_1782_),
    .Y(_0691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3221_ (.B(_1666_),
    .C(_1700_),
    .A(_1644_),
    .Y(_0692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3222_ (.B(_1650_),
    .C(_1652_),
    .A(_1640_),
    .Y(_0693_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1691_));
 sg13g2_o21ai_1 _3223_ (.B1(_1633_),
    .VDD(VPWR),
    .Y(_0694_),
    .VSS(VGND),
    .A1(_0692_),
    .A2(_0693_));
 sg13g2_a21oi_1 _3224_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net734),
    .A2(_1735_),
    .Y(_0695_),
    .B1(_1815_));
 sg13g2_nand2_1 _3225_ (.Y(_0696_),
    .A(net758),
    .B(_1886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3226_ (.B1(_1634_),
    .VDD(VPWR),
    .Y(_0697_),
    .VSS(VGND),
    .A1(_1656_),
    .A2(_1693_));
 sg13g2_a22oi_1 _3227_ (.Y(_0698_),
    .B1(_0697_),
    .B2(_1645_),
    .A2(_1875_),
    .A1(_1775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3228_ (.B(_0695_),
    .C(_0696_),
    .A(_0694_),
    .Y(_0699_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0698_));
 sg13g2_a21oi_1 _3229_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1627_),
    .A2(_1633_),
    .Y(_0700_),
    .B1(_1657_));
 sg13g2_a21oi_1 _3230_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1491_),
    .A2(_1493_),
    .Y(_0701_),
    .B1(_1683_));
 sg13g2_nor3_1 _3231_ (.A(_1633_),
    .B(_0659_),
    .C(_0701_),
    .Y(_0702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3232_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0703_),
    .B(_0702_),
    .A(_0700_));
 sg13g2_nand2_1 _3233_ (.Y(_0704_),
    .A(net730),
    .B(net719),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3234_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0703_),
    .A2(_0704_),
    .Y(_0705_),
    .B1(_1656_));
 sg13g2_a221oi_1 _3235_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1759_),
    .C1(_0705_),
    .B1(_0699_),
    .A1(net741),
    .Y(_0706_),
    .A2(_1775_));
 sg13g2_nor2_2 _3236_ (.A(_1870_),
    .B(_0706_),
    .Y(_0707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3237_ (.Y(_0708_),
    .B(_1869_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0706_));
 sg13g2_nand3_1 _3238_ (.B(_0689_),
    .C(_0708_),
    .A(_0688_),
    .Y(_0709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3239_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0663_),
    .C1(_0650_),
    .B1(_0662_),
    .A1(net740),
    .Y(_0710_),
    .A2(_0647_));
 sg13g2_and2_1 _3240_ (.A(_0707_),
    .B(_0710_),
    .X(_0711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3241_ (.A(_0667_),
    .B(net689),
    .Y(_0712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3242_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0713_),
    .B(net689),
    .A(_0667_));
 sg13g2_a21o_1 _3243_ (.A2(_0670_),
    .A1(net735),
    .B1(_1709_),
    .X(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3244_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0715_),
    .B(_1744_),
    .A(_1691_));
 sg13g2_nor2_1 _3245_ (.A(_1651_),
    .B(_0631_),
    .Y(_0716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3246_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net764),
    .A2(_0644_),
    .Y(_0717_),
    .B1(_0716_));
 sg13g2_or2_1 _3247_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0718_),
    .B(_1744_),
    .A(_1650_));
 sg13g2_and4_1 _3248_ (.A(_0714_),
    .B(_0715_),
    .C(_0717_),
    .D(_0718_),
    .X(_0719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3249_ (.B(_0715_),
    .C(_0717_),
    .A(_0714_),
    .Y(_0720_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0718_));
 sg13g2_a21oi_1 _3250_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net726),
    .A2(net720),
    .Y(_0721_),
    .B1(_0670_));
 sg13g2_nand2_1 _3251_ (.Y(_0722_),
    .A(_0279_),
    .B(_0684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3252_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net725),
    .A2(_1733_),
    .Y(_0723_),
    .B1(_1660_));
 sg13g2_o21ai_1 _3253_ (.B1(_1620_),
    .VDD(VPWR),
    .Y(_0724_),
    .VSS(VGND),
    .A1(_1613_),
    .A2(_1776_));
 sg13g2_nor4_1 _3254_ (.A(_0668_),
    .B(_0722_),
    .C(_0723_),
    .D(_0724_),
    .Y(_0725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3255_ (.B1(_1753_),
    .VDD(VPWR),
    .Y(_0726_),
    .VSS(VGND),
    .A1(_1651_),
    .A2(_0692_));
 sg13g2_nand3_1 _3256_ (.B(_0725_),
    .C(_0726_),
    .A(_0715_),
    .Y(_0727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3257_ (.B1(_0288_),
    .VDD(VPWR),
    .Y(_0728_),
    .VSS(VGND),
    .A1(_0721_),
    .A2(_0727_));
 sg13g2_a22oi_1 _3258_ (.Y(_0729_),
    .B1(_0644_),
    .B2(_1493_),
    .A2(_1586_),
    .A1(_1551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3259_ (.A(_0728_),
    .B(_0729_),
    .X(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3260_ (.Y(_0731_),
    .A(net659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3261_ (.Y(_0732_),
    .A(_0719_),
    .B(net659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3262_ (.Y(_0733_),
    .B1(_0654_),
    .B2(_0691_),
    .A2(_1783_),
    .A1(_1634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3263_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1681_),
    .A2(net721),
    .Y(_0734_),
    .B1(_1653_));
 sg13g2_nand2_1 _3264_ (.Y(_0735_),
    .A(_0635_),
    .B(_0695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3265_ (.A(_1873_),
    .B(_0733_),
    .C(_0734_),
    .D(_0735_),
    .Y(_0736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3266_ (.A(_0319_),
    .B(_0736_),
    .Y(_0737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3267_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0738_),
    .B(_0737_),
    .A(_0643_));
 sg13g2_a21oi_1 _3268_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1569_),
    .A2(_0738_),
    .Y(_0739_),
    .B1(net741));
 sg13g2_nor4_1 _3269_ (.A(_1556_),
    .B(_1870_),
    .C(_0328_),
    .D(_0739_),
    .Y(_0740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3270_ (.B1(net664),
    .VDD(VPWR),
    .Y(_0741_),
    .VSS(VGND),
    .A1(_0732_),
    .A2(_0740_));
 sg13g2_inv_2 _3271_ (.Y(_0742_),
    .A(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3272_ (.Y(_0743_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][0] ),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3273_ (.A(_0719_),
    .B(_0731_),
    .Y(_0744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3274_ (.Y(_0745_),
    .A(_0720_),
    .B(net659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3275_ (.Y(_0746_),
    .A(_0653_),
    .B(_0665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3276_ (.A(_0652_),
    .B(_0664_),
    .C(_0708_),
    .Y(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3277_ (.A(_0653_),
    .B(_0665_),
    .Y(_0748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3278_ (.Y(_0749_),
    .A(_0652_),
    .B(_0664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3279_ (.A(_0653_),
    .B(_0665_),
    .C(_0708_),
    .Y(_0750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3280_ (.Y(_0751_),
    .A(_0707_),
    .B(_0748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3281_ (.Y(_0752_),
    .B1(net681),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .A2(net684),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3282_ (.A(_0652_),
    .B(_0665_),
    .C(_0708_),
    .Y(_0753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3283_ (.Y(_0754_),
    .A(_0666_),
    .B(_0707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3284_ (.Y(_0755_),
    .B1(net677),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .A2(net688),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3285_ (.X(_0756_),
    .A(net662),
    .B(_0752_),
    .C(_0755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3286_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0689_),
    .C1(_0665_),
    .B1(_0688_),
    .A1(_0648_),
    .Y(_0757_),
    .A2(_0651_));
 sg13g2_nand2_2 _3287_ (.Y(_0758_),
    .A(_0666_),
    .B(_0690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3288_ (.A(_0690_),
    .B(_0748_),
    .X(_0759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3289_ (.Y(_0760_),
    .A(_0690_),
    .B(_0748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3290_ (.Y(_0761_),
    .B1(net649),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ),
    .A2(net673),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3291_ (.A(net689),
    .B(_0746_),
    .Y(_0762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3292_ (.A(_0688_),
    .B(_0689_),
    .C(_0708_),
    .D(_0710_),
    .X(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3293_ (.Y(_0764_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .B(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3294_ (.A(net689),
    .B(_0749_),
    .Y(_0765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3295_ (.Y(_0766_),
    .B(_0748_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net689));
 sg13g2_a22oi_1 _3296_ (.Y(_0767_),
    .B1(net639),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .A2(net642),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3297_ (.B(_0761_),
    .C(_0764_),
    .A(_0756_),
    .Y(_0768_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0767_));
 sg13g2_nand2b_1 _3298_ (.Y(_0769_),
    .B(net664),
    .A_N(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3299_ (.A(_0768_),
    .B(_0769_),
    .X(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3300_ (.Y(_0771_),
    .A(_0768_),
    .B(_0769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3301_ (.Y(_0772_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .B(net648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3302_ (.Y(_0773_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .B(net641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3303_ (.Y(_0774_),
    .B1(net680),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .A2(net683),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3304_ (.Y(_0775_),
    .B1(net669),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .A2(net686),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3305_ (.Y(_0776_),
    .B1(net675),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .A2(net665),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3306_ (.Y(_0777_),
    .B1(net638),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .A2(net671),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3307_ (.A(_0774_),
    .B(_0775_),
    .C(_0776_),
    .D(_0777_),
    .X(_0778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3308_ (.X(_0779_),
    .A(_0772_),
    .B(_0773_),
    .C(_0778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3309_ (.B(_0773_),
    .C(_0778_),
    .A(_0772_),
    .Y(_0780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3310_ (.Y(_0781_),
    .B1(net683),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .A2(net686),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3311_ (.Y(_0782_),
    .B1(net638),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3312_ (.Y(_0783_),
    .B1(net669),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .A2(net680),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3313_ (.Y(_0784_),
    .B1(net675),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .A2(net664),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3314_ (.B(_0782_),
    .C(_0783_),
    .A(_0781_),
    .Y(_0785_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0784_));
 sg13g2_a221oi_1 _3315_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .C1(_0785_),
    .B1(net651),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .Y(_0786_),
    .A2(net671));
 sg13g2_a22oi_1 _3316_ (.Y(_0787_),
    .B1(net681),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .A2(net686),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3317_ (.Y(_0788_),
    .B1(net678),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .A2(net684),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3318_ (.Y(_0789_),
    .B1(net642),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .A2(net665),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3319_ (.Y(_0790_),
    .B1(net669),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .A2(net672),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3320_ (.X(_0791_),
    .A(_0787_),
    .B(_0788_),
    .C(_0790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3321_ (.Y(_0792_),
    .B1(net639),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .A2(net649),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3322_ (.X(_0793_),
    .A(_0789_),
    .B(_0791_),
    .C(_0792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3323_ (.B(_0791_),
    .C(_0792_),
    .A(_0789_),
    .Y(_0794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3324_ (.Y(_0795_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .B(net672),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3325_ (.B(_0690_),
    .C(_0748_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .Y(_0796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3326_ (.Y(_0797_),
    .B1(net680),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .A2(net684),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3327_ (.Y(_0798_),
    .B1(net678),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .A2(net686),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3328_ (.A(_0795_),
    .B(_0796_),
    .C(_0797_),
    .D(_0798_),
    .X(_0799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3329_ (.Y(_0800_),
    .B1(net640),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3330_ (.Y(_0801_),
    .B1(net669),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .A2(net665),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3331_ (.X(_0802_),
    .A(_0799_),
    .B(_0800_),
    .C(_0801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3332_ (.B(_0800_),
    .C(_0801_),
    .A(_0799_),
    .Y(_0803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3333_ (.Y(_0804_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .B(net672),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3334_ (.B(_0690_),
    .C(_0748_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .Y(_0805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3335_ (.Y(_0806_),
    .B1(net684),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .A2(net687),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3336_ (.Y(_0807_),
    .B1(net677),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .A2(net682),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3337_ (.B(_0805_),
    .C(_0806_),
    .A(_0804_),
    .Y(_0808_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0807_));
 sg13g2_and2_1 _3338_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .B(net639),
    .X(_0809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3339_ (.A(_1499_),
    .B(net662),
    .Y(_0810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3340_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .B(_0763_),
    .X(_0811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3341_ (.A2(net642),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .B1(_0811_),
    .X(_0812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3342_ (.A(_0808_),
    .B(_0809_),
    .C(_0810_),
    .Y(_0813_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0812_));
 sg13g2_or4_1 _3343_ (.A(_0808_),
    .B(_0809_),
    .C(_0810_),
    .D(_0812_),
    .X(_0814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3344_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .B(net649),
    .X(_0815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3345_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ),
    .B(net673),
    .X(_0816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3346_ (.Y(_0817_),
    .B1(net681),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .A2(net687),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3347_ (.Y(_0818_),
    .B1(net677),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .A2(net684),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3348_ (.Y(_0819_),
    .A(_0817_),
    .B(_0818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3349_ (.A(_1522_),
    .B(net690),
    .C(_0749_),
    .Y(_0820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3350_ (.A(_1523_),
    .B(net690),
    .C(_0746_),
    .Y(_0821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3351_ (.A(_1524_),
    .B(_0667_),
    .C(net690),
    .Y(_0822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3352_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .B(net670),
    .X(_0823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _3353_ (.A(_0820_),
    .B(_0821_),
    .C(_0822_),
    .D(_0823_),
    .X(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3354_ (.A(_0815_),
    .B(_0816_),
    .C(_0819_),
    .Y(_0825_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0824_));
 sg13g2_nand3_1 _3355_ (.B(_0690_),
    .C(_0748_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .Y(_0826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3356_ (.Y(_0827_),
    .B1(net681),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .A2(net688),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3357_ (.Y(_0828_),
    .B1(net677),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .A2(net684),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3358_ (.Y(_0829_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .B(net673),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3359_ (.A(_0826_),
    .B(_0827_),
    .C(_0828_),
    .D(_0829_),
    .X(_0830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3360_ (.A(_1507_),
    .B(_0667_),
    .C(net690),
    .Y(_0831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3361_ (.A(_1506_),
    .B(net690),
    .C(_0746_),
    .Y(_0832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3362_ (.A(_1505_),
    .B(net690),
    .C(_0749_),
    .Y(_0833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3363_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .B(net670),
    .X(_0834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3364_ (.A(_0831_),
    .B(_0832_),
    .C(_0833_),
    .D(_0834_),
    .Y(_0835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3365_ (.A(_0830_),
    .B(_0835_),
    .X(_0836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3366_ (.B(_0690_),
    .C(_0748_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .Y(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3367_ (.Y(_0838_),
    .B1(net680),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .A2(net688),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3368_ (.Y(_0839_),
    .B1(net677),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .A2(net683),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3369_ (.Y(_0840_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .B(net671),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3370_ (.A(_0837_),
    .B(_0838_),
    .C(_0839_),
    .D(_0840_),
    .X(_0841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3371_ (.A(_1519_),
    .B(_0667_),
    .C(net689),
    .Y(_0842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3372_ (.A(_1517_),
    .B(net689),
    .C(_0749_),
    .Y(_0843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3373_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .B(net670),
    .X(_0844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3374_ (.A(_1518_),
    .B(net689),
    .C(_0746_),
    .Y(_0845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3375_ (.A(_0842_),
    .B(_0843_),
    .C(_0844_),
    .D(_0845_),
    .Y(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3376_ (.A(_0841_),
    .B(_0846_),
    .X(_0847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3377_ (.Y(_0848_),
    .A(net589),
    .B(_0847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3378_ (.B(_0836_),
    .C(_0847_),
    .A(net591),
    .Y(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3379_ (.A(_0813_),
    .B(net591),
    .C(_0836_),
    .D(_0847_),
    .X(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3380_ (.B(_0802_),
    .C(_0850_),
    .A(_0793_),
    .Y(_0851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3381_ (.B(_0793_),
    .C(_0802_),
    .A(_0786_),
    .Y(_0852_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0850_));
 sg13g2_nor3_1 _3382_ (.A(_0770_),
    .B(_0780_),
    .C(_0852_),
    .Y(_0853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3383_ (.B1(_0770_),
    .VDD(VPWR),
    .Y(_0854_),
    .VSS(VGND),
    .A1(_0780_),
    .A2(_0852_));
 sg13g2_nand2b_2 _3384_ (.Y(_0855_),
    .B(_0854_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0853_));
 sg13g2_nor2_1 _3385_ (.A(net612),
    .B(_0855_),
    .Y(_0856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3386_ (.A(_0720_),
    .B(net659),
    .Y(_0857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3387_ (.Y(_0858_),
    .A(_0719_),
    .B(_0731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3388_ (.Y(_0859_),
    .B1(_0841_),
    .B2(_0846_),
    .A2(_0835_),
    .A1(_0830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3389_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0860_),
    .B(_0847_),
    .A(_0836_));
 sg13g2_nand2_2 _3390_ (.Y(_0861_),
    .A(_0814_),
    .B(_0859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3391_ (.B(_0814_),
    .C(_0859_),
    .A(_0803_),
    .Y(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3392_ (.B(_0803_),
    .C(_0814_),
    .A(_0794_),
    .Y(_0863_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0859_));
 sg13g2_or2_1 _3393_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0864_),
    .B(_0863_),
    .A(_0786_));
 sg13g2_nor4_2 _3394_ (.A(_0771_),
    .B(_0779_),
    .C(_0786_),
    .Y(_0865_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0863_));
 sg13g2_or2_1 _3395_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0866_),
    .B(_0862_),
    .A(net591));
 sg13g2_nor2_1 _3396_ (.A(net589),
    .B(_0863_),
    .Y(_0867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3397_ (.A(_0779_),
    .B(net589),
    .C(_0864_),
    .Y(_0868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3398_ (.Y(_0869_),
    .A(_0770_),
    .B(_0868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3399_ (.Y(_0870_),
    .A(net608),
    .B(_0869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3400_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1645_),
    .C1(_0723_),
    .B1(_0672_),
    .A1(net734),
    .Y(_0871_),
    .A2(_1705_));
 sg13g2_and3_1 _3401_ (.X(_0872_),
    .A(_0679_),
    .B(_0682_),
    .C(_0871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3402_ (.B1(_1620_),
    .VDD(VPWR),
    .Y(_0873_),
    .VSS(VGND),
    .A1(_0669_),
    .A2(_0872_));
 sg13g2_a221oi_1 _3403_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0873_),
    .C1(_0644_),
    .B1(_0288_),
    .A1(_1551_),
    .Y(_0874_),
    .A2(net737));
 sg13g2_nor2_2 _3404_ (.A(net660),
    .B(net668),
    .Y(_0875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3405_ (.Y(_0876_),
    .B(net664),
    .A_N(net668),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3406_ (.Y(_0877_),
    .A(net31),
    .B(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3407_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net9),
    .A2(_0875_),
    .Y(_0878_),
    .B1(_0732_));
 sg13g2_a21oi_1 _3408_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0877_),
    .A2(_0878_),
    .Y(_0879_),
    .B1(net596));
 sg13g2_nand2_1 _3409_ (.Y(_0880_),
    .A(_0870_),
    .B(_0879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3410_ (.Y(_0881_),
    .A(_0720_),
    .B(_0731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3411_ (.B1(_0743_),
    .VDD(VPWR),
    .Y(_0066_),
    .VSS(VGND),
    .A1(_0856_),
    .A2(_0880_));
 sg13g2_or2_1 _3412_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0882_),
    .B(_0847_),
    .A(net589));
 sg13g2_nand2_2 _3413_ (.Y(_0883_),
    .A(_0848_),
    .B(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3414_ (.Y(_0884_),
    .A(net660),
    .B(_0883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3415_ (.Y(_0885_),
    .B1(net683),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .A2(net688),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3416_ (.Y(_0886_),
    .B1(net675),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .A2(net680),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3417_ (.B(_0885_),
    .C(_0886_),
    .A(net660),
    .Y(_0887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3418_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ),
    .C1(_0887_),
    .B1(net648),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ),
    .Y(_0888_),
    .A2(net671));
 sg13g2_nor2_1 _3419_ (.A(_1518_),
    .B(net637),
    .Y(_0889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3420_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .C1(_0889_),
    .B1(net670),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .Y(_0890_),
    .A2(net641));
 sg13g2_a22oi_1 _3421_ (.Y(_0891_),
    .B1(_0888_),
    .B2(_0890_),
    .A2(net665),
    .A1(_1510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3422_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0892_),
    .B(_0891_),
    .A(_0770_));
 sg13g2_or3_1 _3423_ (.A(_0780_),
    .B(_0852_),
    .C(_0892_),
    .X(_0893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3424_ (.Y(_0894_),
    .A(_0853_),
    .B(_0891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3425_ (.B1(_0884_),
    .VDD(VPWR),
    .Y(_0895_),
    .VSS(VGND),
    .A1(net660),
    .A2(_0894_));
 sg13g2_nand2_1 _3426_ (.Y(_0896_),
    .A(net594),
    .B(_0895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3427_ (.Y(_0897_),
    .A(_0865_),
    .B(_0891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3428_ (.A(net589),
    .B(_0897_),
    .Y(_0898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3429_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0770_),
    .A2(_0868_),
    .Y(_0899_),
    .B1(_0891_));
 sg13g2_or2_1 _3430_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0900_),
    .B(_0899_),
    .A(_0898_));
 sg13g2_inv_1 _3431_ (.VDD(VPWR),
    .Y(_0901_),
    .A(_0900_),
    .VSS(VGND));
 sg13g2_a21oi_1 _3432_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net664),
    .A2(_0900_),
    .Y(_0902_),
    .B1(net587));
 sg13g2_nor2_1 _3433_ (.A(net10),
    .B(net605),
    .Y(_0903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3434_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2051_),
    .A2(net605),
    .Y(_0904_),
    .B1(_0903_));
 sg13g2_nor3_1 _3435_ (.A(net596),
    .B(_0902_),
    .C(_0904_),
    .Y(_0905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3436_ (.Y(_0067_),
    .B1(_0896_),
    .B2(_0905_),
    .A2(net596),
    .A1(_1510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3437_ (.Y(_0906_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][2] ),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3438_ (.Y(_0907_),
    .B1(net677),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .A2(net688),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3439_ (.Y(_0908_),
    .B1(net681),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .A2(net684),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3440_ (.X(_0909_),
    .A(net662),
    .B(_0907_),
    .C(_0908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3441_ (.Y(_0910_),
    .B1(net649),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ),
    .A2(net673),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3442_ (.Y(_0911_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .B(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3443_ (.Y(_0912_),
    .B1(net639),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .A2(net642),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3444_ (.B(_0910_),
    .C(_0911_),
    .A(_0909_),
    .Y(_0913_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0912_));
 sg13g2_o21ai_1 _3445_ (.B1(_0913_),
    .VDD(VPWR),
    .Y(_0914_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][2] ),
    .A2(net662));
 sg13g2_inv_1 _3446_ (.VDD(VPWR),
    .Y(_0915_),
    .A(_0914_),
    .VSS(VGND));
 sg13g2_nand2b_1 _3447_ (.Y(_0916_),
    .B(_0914_),
    .A_N(_0893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3448_ (.Y(_0917_),
    .A(_0893_),
    .B(_0915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3449_ (.A(net660),
    .B(_0917_),
    .Y(_0918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3450_ (.Y(_0919_),
    .A(_0836_),
    .B(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3451_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net661),
    .A2(_0919_),
    .Y(_0920_),
    .B1(_0918_));
 sg13g2_nand2_1 _3452_ (.Y(_0921_),
    .A(_0227_),
    .B(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3453_ (.Y(_0922_),
    .B(_0875_),
    .A_N(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3454_ (.Y(_0923_),
    .A(_0836_),
    .B(_0847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3455_ (.A(_0719_),
    .B(net648),
    .Y(_0924_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3456_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net659),
    .Y(_0925_),
    .A2(_0924_),
    .A1(_0923_));
 sg13g2_a221oi_1 _3457_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0922_),
    .C1(_0925_),
    .B1(_0921_),
    .A1(net594),
    .Y(_0926_),
    .A2(_0920_));
 sg13g2_nand3_1 _3458_ (.B(_0891_),
    .C(_0915_),
    .A(_0865_),
    .Y(_0927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3459_ (.Y(_0928_),
    .A(_0898_),
    .B(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3460_ (.A(net587),
    .B(_0928_),
    .Y(_0929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3461_ (.A(net591),
    .B(_0860_),
    .Y(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3462_ (.Y(_0931_),
    .A(_0836_),
    .B(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3463_ (.B1(_0742_),
    .VDD(VPWR),
    .Y(_0932_),
    .VSS(VGND),
    .A1(net587),
    .A2(_0928_));
 sg13g2_o21ai_1 _3464_ (.B1(_0906_),
    .VDD(VPWR),
    .Y(_0068_),
    .VSS(VGND),
    .A1(_0926_),
    .A2(_0932_));
 sg13g2_a22oi_1 _3465_ (.Y(_0933_),
    .B1(net685),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .A2(net687),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3466_ (.Y(_0934_),
    .B1(net678),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .A2(net682),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3467_ (.X(_0935_),
    .A(net662),
    .B(_0933_),
    .C(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3468_ (.Y(_0936_),
    .B1(net650),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ),
    .A2(net673),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3469_ (.Y(_0937_),
    .B1(net639),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .A2(net642),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3470_ (.Y(_0938_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .B(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3471_ (.B(_0936_),
    .C(_0937_),
    .A(_0935_),
    .Y(_0939_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0938_));
 sg13g2_o21ai_1 _3472_ (.B1(_0939_),
    .VDD(VPWR),
    .Y(_0940_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][3] ),
    .A2(net662));
 sg13g2_inv_1 _3473_ (.VDD(VPWR),
    .Y(_0941_),
    .A(_0940_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3474_ (.B1(_0940_),
    .VDD(VPWR),
    .Y(_0942_),
    .VSS(VGND),
    .A1(_0825_),
    .A2(_0927_));
 sg13g2_nand4_1 _3475_ (.B(_0891_),
    .C(_0915_),
    .A(_0865_),
    .Y(_0943_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0941_));
 sg13g2_nor2_1 _3476_ (.A(net590),
    .B(net571),
    .Y(_0944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3477_ (.B1(_0942_),
    .VDD(VPWR),
    .Y(_0945_),
    .VSS(VGND),
    .A1(_0825_),
    .A2(net572));
 sg13g2_xnor2_1 _3478_ (.Y(_0946_),
    .A(_0813_),
    .B(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3479_ (.B1(net611),
    .VDD(VPWR),
    .Y(_0947_),
    .VSS(VGND),
    .A1(net665),
    .A2(_0946_));
 sg13g2_a21oi_1 _3480_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net665),
    .A2(_0945_),
    .Y(_0948_),
    .B1(_0947_));
 sg13g2_nand2_1 _3481_ (.Y(_0949_),
    .A(_0914_),
    .B(_0940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3482_ (.A(_0780_),
    .B(_0852_),
    .C(_0892_),
    .Y(_0950_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0949_));
 sg13g2_xnor2_1 _3483_ (.Y(_0951_),
    .A(_0916_),
    .B(_0940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3484_ (.Y(_0952_),
    .A(_0813_),
    .B(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3485_ (.A2(_0952_),
    .A1(_0713_),
    .B1(net613),
    .X(_0953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3486_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net665),
    .A2(_0951_),
    .Y(_0954_),
    .B1(_0953_));
 sg13g2_nor2_1 _3487_ (.A(net32),
    .B(_0875_),
    .Y(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3488_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0303_),
    .A2(_0875_),
    .Y(_0956_),
    .B1(_0955_));
 sg13g2_a21oi_1 _3489_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0813_),
    .A2(_0860_),
    .Y(_0957_),
    .B1(_0881_));
 sg13g2_nor4_1 _3490_ (.A(net597),
    .B(_0948_),
    .C(_0954_),
    .D(_0956_),
    .Y(_0958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3491_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1497_),
    .A2(net597),
    .Y(_0069_),
    .B1(_0958_));
 sg13g2_nand2_1 _3492_ (.Y(_0959_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][4] ),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3493_ (.Y(_0960_),
    .B1(net678),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .A2(net686),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3494_ (.Y(_0961_),
    .B1(net682),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .A2(net685),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3495_ (.B(_0960_),
    .C(_0961_),
    .A(net661),
    .Y(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3496_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .C1(_0962_),
    .B1(net647),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .Y(_0963_),
    .A2(net674));
 sg13g2_nand2_1 _3497_ (.Y(_0964_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .B(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3498_ (.Y(_0965_),
    .B1(net669),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3499_ (.B(_0964_),
    .C(_0965_),
    .A(_0963_),
    .Y(_0966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3500_ (.B1(_0966_),
    .VDD(VPWR),
    .Y(_0967_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][4] ),
    .A2(net661));
 sg13g2_xor2_1 _3501_ (.B(net573),
    .A(_0950_),
    .X(_0968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3502_ (.Y(_0969_),
    .A(_0802_),
    .B(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3503_ (.B1(net592),
    .VDD(VPWR),
    .Y(_0970_),
    .VSS(VGND),
    .A1(net663),
    .A2(_0969_));
 sg13g2_a21oi_1 _3504_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net663),
    .A2(_0968_),
    .Y(_0971_),
    .B1(_0970_));
 sg13g2_mux2_1 _3505_ (.A0(net21),
    .A1(net13),
    .S(_0875_),
    .X(_0972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3506_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0802_),
    .A2(_0861_),
    .Y(_0973_),
    .B1(net585));
 sg13g2_nand2_1 _3507_ (.Y(_0974_),
    .A(_0862_),
    .B(_0973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3508_ (.Y(_0975_),
    .A(net588),
    .B(_0974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3509_ (.A(_0971_),
    .B(_0972_),
    .C(_0975_),
    .Y(_0976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3510_ (.A(net571),
    .B(net574),
    .Y(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3511_ (.A(net590),
    .B(net571),
    .C(net573),
    .Y(_0978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3512_ (.Y(_0979_),
    .A(_0944_),
    .B(net573),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3513_ (.B1(_0742_),
    .VDD(VPWR),
    .Y(_0980_),
    .VSS(VGND),
    .A1(net586),
    .A2(_0979_));
 sg13g2_o21ai_1 _3514_ (.B1(_0802_),
    .VDD(VPWR),
    .Y(_0981_),
    .VSS(VGND),
    .A1(net591),
    .A2(_0861_));
 sg13g2_o21ai_1 _3515_ (.B1(_0959_),
    .VDD(VPWR),
    .Y(_0070_),
    .VSS(VGND),
    .A1(_0976_),
    .A2(_0980_));
 sg13g2_nand2_1 _3516_ (.Y(_0982_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][5] ),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3517_ (.Y(_0983_),
    .B1(net681),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .A2(net684),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3518_ (.Y(_0984_),
    .B1(net678),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .A2(net687),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3519_ (.B(_0983_),
    .C(_0984_),
    .A(net662),
    .Y(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3520_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .C1(_0985_),
    .B1(net649),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .Y(_0986_),
    .A2(net672));
 sg13g2_nand2_1 _3521_ (.Y(_0987_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .B(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3522_ (.Y(_0988_),
    .B1(net640),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .A2(net642),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3523_ (.B(_0987_),
    .C(_0988_),
    .A(_0986_),
    .Y(_0989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3524_ (.B1(_0989_),
    .VDD(VPWR),
    .Y(_0990_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][5] ),
    .A2(net661));
 sg13g2_and2_1 _3525_ (.A(net573),
    .B(_0990_),
    .X(_0991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3526_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0950_),
    .A2(net574),
    .Y(_0992_),
    .B1(_0990_));
 sg13g2_a21oi_2 _3527_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0992_),
    .Y(_0993_),
    .A2(_0991_),
    .A1(_0950_));
 sg13g2_a21o_1 _3528_ (.A2(_0850_),
    .A1(_0802_),
    .B1(_0793_),
    .X(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3529_ (.Y(_0995_),
    .A(_0851_),
    .B(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3530_ (.B1(net593),
    .VDD(VPWR),
    .Y(_0996_),
    .VSS(VGND),
    .A1(net663),
    .A2(_0995_));
 sg13g2_a21oi_1 _3531_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net663),
    .A2(_0993_),
    .Y(_0997_),
    .B1(_0996_));
 sg13g2_nor2_1 _3532_ (.A(net14),
    .B(net605),
    .Y(_0998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3533_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net569),
    .A2(net606),
    .Y(_0999_),
    .B1(_0998_));
 sg13g2_a21oi_1 _3534_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0793_),
    .A2(_0862_),
    .Y(_1000_),
    .B1(net585));
 sg13g2_nand2_1 _3535_ (.Y(_1001_),
    .A(_0863_),
    .B(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3536_ (.Y(_1002_),
    .A(net588),
    .B(_1001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3537_ (.A(_0997_),
    .B(_0999_),
    .C(_1002_),
    .Y(_1003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3538_ (.A(net571),
    .B(net574),
    .C(_0990_),
    .Y(_1004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _3539_ (.A(net590),
    .B(net571),
    .C(net573),
    .D(_0990_),
    .X(_1005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3540_ (.Y(_1006_),
    .A(_0978_),
    .B(_0990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3541_ (.A(net586),
    .B(_1006_),
    .Y(_1007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3542_ (.B1(_0742_),
    .VDD(VPWR),
    .Y(_1008_),
    .VSS(VGND),
    .A1(net586),
    .A2(_1006_));
 sg13g2_xnor2_1 _3543_ (.Y(_1009_),
    .A(_0793_),
    .B(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3544_ (.B1(_0982_),
    .VDD(VPWR),
    .Y(_0071_),
    .VSS(VGND),
    .A1(_1003_),
    .A2(_1008_));
 sg13g2_a22oi_1 _3545_ (.Y(_1010_),
    .B1(net680),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .A2(net683),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3546_ (.Y(_1011_),
    .B1(net675),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .A2(net686),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3547_ (.B(_1010_),
    .C(_1011_),
    .A(net661),
    .Y(_1012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3548_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ),
    .C1(_1012_),
    .B1(net647),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .Y(_1013_),
    .A2(net671));
 sg13g2_a22oi_1 _3549_ (.Y(_1014_),
    .B1(net640),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3550_ (.Y(_1015_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .B(net669),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3551_ (.B(_1014_),
    .C(_1015_),
    .A(_1013_),
    .Y(_1016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3552_ (.B1(_1016_),
    .VDD(VPWR),
    .Y(_1017_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][6] ),
    .A2(net661));
 sg13g2_nor4_1 _3553_ (.A(net571),
    .B(net573),
    .C(_0990_),
    .D(_1017_),
    .Y(_1018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3554_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1019_),
    .B(_1017_),
    .A(_0990_));
 sg13g2_nor4_1 _3555_ (.A(net590),
    .B(net571),
    .C(net573),
    .D(_1019_),
    .Y(_1020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3556_ (.A2(_1017_),
    .A1(_1005_),
    .B1(_1020_),
    .X(_1021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3557_ (.Y(_1022_),
    .A(_0786_),
    .B(_0867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3558_ (.B1(net609),
    .VDD(VPWR),
    .Y(_1023_),
    .VSS(VGND),
    .A1(net663),
    .A2(_1022_));
 sg13g2_a21oi_1 _3559_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net663),
    .A2(_1021_),
    .Y(_1024_),
    .B1(_1023_));
 sg13g2_nand3_1 _3560_ (.B(_0991_),
    .C(_1017_),
    .A(_0950_),
    .Y(_1025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3561_ (.A2(_0991_),
    .A1(_0950_),
    .B1(_1017_),
    .X(_1026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3562_ (.A(_1025_),
    .B(_1026_),
    .X(_1027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3563_ (.B(_0851_),
    .A(_0786_),
    .X(_1028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3564_ (.B1(net592),
    .VDD(VPWR),
    .Y(_1029_),
    .VSS(VGND),
    .A1(net663),
    .A2(_1028_));
 sg13g2_a21oi_1 _3565_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net663),
    .A2(_1027_),
    .Y(_1030_),
    .B1(_1029_));
 sg13g2_nor2_1 _3566_ (.A(net15),
    .B(net605),
    .Y(_1031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3567_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net570),
    .A2(net605),
    .Y(_1032_),
    .B1(_1031_));
 sg13g2_nor4_1 _3568_ (.A(net597),
    .B(_1024_),
    .C(_1030_),
    .D(_1032_),
    .Y(_1033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3569_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1539_),
    .A2(net597),
    .Y(_0072_),
    .B1(_1033_));
 sg13g2_a22oi_1 _3570_ (.Y(_1034_),
    .B1(net675),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .A2(net683),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3571_ (.Y(_1035_),
    .B1(net680),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .A2(net686),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3572_ (.B(_1034_),
    .C(_1035_),
    .A(net660),
    .Y(_1036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3573_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .C1(_1036_),
    .B1(net648),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .Y(_1037_),
    .A2(net671));
 sg13g2_and2_1 _3574_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .B(net669),
    .X(_1038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3575_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .C1(_1038_),
    .B1(net638),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .Y(_1039_),
    .A2(net641));
 sg13g2_a22oi_1 _3576_ (.Y(_1040_),
    .B1(_1037_),
    .B2(_1039_),
    .A2(net664),
    .A1(_1545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3577_ (.B(_1040_),
    .A(_1025_),
    .X(_1041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3578_ (.Y(_1042_),
    .A(net664),
    .B(_1041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3579_ (.Y(_1043_),
    .A(_0779_),
    .B(_0852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3580_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net660),
    .A2(_1043_),
    .Y(_1044_),
    .B1(net612));
 sg13g2_xor2_1 _3581_ (.B(_1040_),
    .A(_1020_),
    .X(_1045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3582_ (.B1(_0779_),
    .VDD(VPWR),
    .Y(_1046_),
    .VSS(VGND),
    .A1(net589),
    .A2(_0864_));
 sg13g2_nor2b_2 _3583_ (.A(_0868_),
    .B_N(_1046_),
    .Y(_1047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3584_ (.A0(_1045_),
    .A1(_1047_),
    .S(net660),
    .X(_1048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3585_ (.A(_0306_),
    .B(net605),
    .Y(_1049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3586_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net24),
    .A2(net606),
    .Y(_1050_),
    .B1(_1049_));
 sg13g2_nand2_1 _3587_ (.Y(_1051_),
    .A(_0742_),
    .B(_1050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3588_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net607),
    .C1(_1051_),
    .B1(_1048_),
    .A1(_1042_),
    .Y(_1052_),
    .A2(_1044_));
 sg13g2_a21oi_1 _3589_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1545_),
    .A2(net597),
    .Y(_0073_),
    .B1(_1052_));
 sg13g2_nor2_1 _3590_ (.A(net641),
    .B(_0875_),
    .Y(_1053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3591_ (.Y(_1054_),
    .B(net606),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net642));
 sg13g2_and2_1 _3592_ (.A(net595),
    .B(net589),
    .X(_1055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3593_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0720_),
    .A2(net589),
    .Y(_1056_),
    .B1(net659));
 sg13g2_nor3_2 _3594_ (.A(net31),
    .B(_1055_),
    .C(_1056_),
    .Y(_1057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3595_ (.A(net591),
    .B(net588),
    .Y(_1058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3596_ (.A(net583),
    .B(_1057_),
    .C(_1058_),
    .X(_1059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3597_ (.B1(_1059_),
    .VDD(VPWR),
    .Y(_0074_),
    .VSS(VGND),
    .A1(_1524_),
    .A2(_1054_));
 sg13g2_nor2_2 _3598_ (.A(net588),
    .B(_0883_),
    .Y(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3599_ (.A(net583),
    .B(_1060_),
    .Y(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3600_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0848_),
    .A2(_0882_),
    .Y(_1062_),
    .B1(net612));
 sg13g2_nor2b_2 _3601_ (.A(_1062_),
    .B_N(_2051_),
    .Y(_1063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3602_ (.Y(_0075_),
    .B1(_1061_),
    .B2(_1063_),
    .A2(net583),
    .A1(_1519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3603_ (.A(net613),
    .B(_0919_),
    .Y(_1064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3604_ (.A(net19),
    .B(_1064_),
    .Y(_1065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3605_ (.A(net588),
    .B(_0931_),
    .Y(_1066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3606_ (.A(net583),
    .B(_1066_),
    .Y(_1067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3607_ (.Y(_0076_),
    .B1(_1065_),
    .B2(_1067_),
    .A2(net583),
    .A1(_1507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3608_ (.A(net613),
    .B(_0952_),
    .Y(_1068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3609_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1069_),
    .B(_1068_),
    .A(net32));
 sg13g2_a21oi_2 _3610_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1069_),
    .Y(_1070_),
    .A2(_0957_),
    .A1(_0861_));
 sg13g2_and2_1 _3611_ (.A(net611),
    .B(_0946_),
    .X(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3612_ (.A(net583),
    .B(_1071_),
    .Y(_1072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3613_ (.Y(_0077_),
    .B1(_1070_),
    .B2(_1072_),
    .A2(net583),
    .A1(_1499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3614_ (.A(net592),
    .B(_0969_),
    .X(_1073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3615_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1074_),
    .B(_1073_),
    .A(net21));
 sg13g2_nand3_1 _3616_ (.B(_0866_),
    .C(_0981_),
    .A(net611),
    .Y(_1075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3617_ (.A(net583),
    .B(_1074_),
    .Y(_1076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3618_ (.Y(_0078_),
    .B1(_1075_),
    .B2(_1076_),
    .A2(net584),
    .A1(_1535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3619_ (.Y(_1077_),
    .A(net595),
    .B(_0995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3620_ (.A(net569),
    .B(_1077_),
    .X(_1078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3621_ (.Y(_1079_),
    .B(_1078_),
    .A_N(_1002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3622_ (.Y(_1080_),
    .A(net611),
    .B(_1009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3623_ (.Y(_1081_),
    .A(_1079_),
    .B(_1080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3624_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ),
    .B(_1054_),
    .Y(_1082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3625_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1054_),
    .A2(_1081_),
    .Y(_0079_),
    .B1(_1082_));
 sg13g2_nand2_1 _3626_ (.Y(_1083_),
    .A(net593),
    .B(_1028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3627_ (.Y(_1084_),
    .A(net570),
    .B(_1083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3628_ (.Y(_1085_),
    .A(net609),
    .B(_1022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3629_ (.A(net584),
    .B(_1084_),
    .Y(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3630_ (.Y(_0080_),
    .B1(_1085_),
    .B2(_1086_),
    .A2(net584),
    .A1(_1544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3631_ (.A(net612),
    .B(_1043_),
    .Y(_1087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3632_ (.Y(_1088_),
    .A(_0779_),
    .B(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3633_ (.B1(net587),
    .VDD(VPWR),
    .Y(_1089_),
    .VSS(VGND),
    .A1(net585),
    .A2(_1088_));
 sg13g2_nor3_2 _3634_ (.A(net24),
    .B(_1087_),
    .C(_1089_),
    .Y(_1090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3635_ (.Y(_1091_),
    .B(net610),
    .A_N(_1047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3636_ (.Y(_1092_),
    .A(_1091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3637_ (.A(net584),
    .B(_1090_),
    .C(_1092_),
    .Y(_1093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3638_ (.A2(net584),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .B1(_1093_),
    .X(_0081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3639_ (.Y(_1094_),
    .A(net595),
    .B(_0855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3640_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net595),
    .A2(_0855_),
    .Y(_1095_),
    .B1(_1056_));
 sg13g2_nor2_1 _3641_ (.A(net636),
    .B(net668),
    .Y(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3642_ (.Y(_1097_),
    .A(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3643_ (.Y(_1098_),
    .A(_0301_),
    .B(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3644_ (.B1(_1098_),
    .VDD(VPWR),
    .Y(_1099_),
    .VSS(VGND),
    .A1(net31),
    .A2(net604));
 sg13g2_nand2_1 _3645_ (.Y(_1100_),
    .A(net637),
    .B(_1055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3646_ (.B(_1099_),
    .C(_1100_),
    .A(_1095_),
    .Y(_1101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3647_ (.B(_0870_),
    .C(_1101_),
    .A(net639),
    .Y(_1102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3648_ (.B1(_1102_),
    .VDD(VPWR),
    .Y(_0082_),
    .VSS(VGND),
    .A1(_1523_),
    .A2(net639));
 sg13g2_nand2_1 _3649_ (.Y(_1103_),
    .A(net594),
    .B(_0894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3650_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1104_),
    .B(net668),
    .A(_0302_));
 sg13g2_a21oi_1 _3651_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net18),
    .A2(_1097_),
    .Y(_1105_),
    .B1(_0732_));
 sg13g2_a221oi_1 _3652_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1105_),
    .C1(net636),
    .B1(_1104_),
    .A1(net607),
    .Y(_1106_),
    .A2(_0900_));
 sg13g2_a22oi_1 _3653_ (.Y(_1107_),
    .B1(_1103_),
    .B2(_1106_),
    .A2(net636),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3654_ (.VDD(VPWR),
    .Y(_0083_),
    .A(_1107_),
    .VSS(VGND));
 sg13g2_nand2_1 _3655_ (.Y(_1108_),
    .A(net637),
    .B(_0919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3656_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0917_),
    .A2(_1108_),
    .Y(_1109_),
    .B1(net613));
 sg13g2_nand2_1 _3657_ (.Y(_1110_),
    .A(_0227_),
    .B(net668),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3658_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net11),
    .C1(_0732_),
    .B1(net604),
    .A1(net19),
    .Y(_1111_),
    .A2(_0874_));
 sg13g2_or4_1 _3659_ (.A(net637),
    .B(_0929_),
    .C(_1109_),
    .D(_1111_),
    .X(_1112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3660_ (.B1(_1112_),
    .VDD(VPWR),
    .Y(_0084_),
    .VSS(VGND),
    .A1(_1506_),
    .A2(net639));
 sg13g2_a21oi_1 _3661_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net32),
    .A2(_1097_),
    .Y(_1113_),
    .B1(_0732_));
 sg13g2_o21ai_1 _3662_ (.B1(_1113_),
    .VDD(VPWR),
    .Y(_1114_),
    .VSS(VGND),
    .A1(_0303_),
    .A2(net668));
 sg13g2_a221oi_1 _3663_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net595),
    .C1(_0766_),
    .B1(_0951_),
    .A1(_0857_),
    .Y(_1115_),
    .A2(_0945_));
 sg13g2_a22oi_1 _3664_ (.Y(_1116_),
    .B1(_1114_),
    .B2(_1115_),
    .A2(net637),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3665_ (.VDD(VPWR),
    .Y(_0085_),
    .A(_1116_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3666_ (.B1(net592),
    .VDD(VPWR),
    .Y(_1117_),
    .VSS(VGND),
    .A1(net638),
    .A2(_0969_));
 sg13g2_nor2_1 _3667_ (.A(_0968_),
    .B(_1117_),
    .Y(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3668_ (.A(net609),
    .B(_0979_),
    .X(_1119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3669_ (.Y(_1120_),
    .A(net609),
    .B(_0979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3670_ (.A(net13),
    .B(_1097_),
    .Y(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3671_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1991_),
    .A2(_1097_),
    .Y(_1122_),
    .B1(_1121_));
 sg13g2_nor3_1 _3672_ (.A(net636),
    .B(_1118_),
    .C(_1122_),
    .Y(_1123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3673_ (.Y(_0086_),
    .B1(_1120_),
    .B2(_1123_),
    .A2(net636),
    .A1(_1534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3674_ (.A(net610),
    .B(_1006_),
    .X(_1124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3675_ (.Y(_1125_),
    .A(net609),
    .B(_1006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3676_ (.A(net638),
    .B(_0995_),
    .Y(_1126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3677_ (.Y(_1127_),
    .A(net14),
    .B(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3678_ (.B1(_1127_),
    .VDD(VPWR),
    .Y(_1128_),
    .VSS(VGND),
    .A1(net569),
    .A2(net604));
 sg13g2_nor3_1 _3679_ (.A(net612),
    .B(_0993_),
    .C(_1126_),
    .Y(_1129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3680_ (.A(net636),
    .B(_1128_),
    .C(_1129_),
    .Y(_1130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3681_ (.Y(_0087_),
    .B1(_1125_),
    .B2(_1130_),
    .A2(net637),
    .A1(_1538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3682_ (.Y(_1131_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .B(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3683_ (.Y(_1132_),
    .A(net609),
    .B(_1021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3684_ (.Y(_1133_),
    .A(net638),
    .B(_1132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3685_ (.B1(net592),
    .VDD(VPWR),
    .Y(_1134_),
    .VSS(VGND),
    .A1(net638),
    .A2(_1028_));
 sg13g2_nor2_1 _3686_ (.A(_1027_),
    .B(_1134_),
    .Y(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3687_ (.A(net15),
    .B(_1097_),
    .Y(_1136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3688_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net570),
    .A2(_1097_),
    .Y(_1137_),
    .B1(_1136_));
 sg13g2_nand2_1 _3689_ (.Y(_1138_),
    .A(_0786_),
    .B(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3690_ (.A(_0720_),
    .B(_0731_),
    .C(_0864_),
    .D(_1138_),
    .X(_1139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3691_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1140_),
    .B(_1139_),
    .A(net609));
 sg13g2_nor3_1 _3692_ (.A(_1135_),
    .B(_1137_),
    .C(_1140_),
    .Y(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3693_ (.B1(_1131_),
    .VDD(VPWR),
    .Y(_0088_),
    .VSS(VGND),
    .A1(_1133_),
    .A2(_1141_));
 sg13g2_nor2_1 _3694_ (.A(net612),
    .B(_1041_),
    .Y(_1142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3695_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0306_),
    .C1(_0732_),
    .B1(net604),
    .A1(_1914_),
    .Y(_1143_),
    .A2(net668));
 sg13g2_nor3_1 _3696_ (.A(net636),
    .B(_1142_),
    .C(_1143_),
    .Y(_1144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3697_ (.Y(_1145_),
    .A(net608),
    .B(_1045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3698_ (.Y(_0089_),
    .B1(_1144_),
    .B2(_1145_),
    .A2(net636),
    .A1(_1548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3699_ (.A(net670),
    .B(net604),
    .Y(_1146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3700_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1147_),
    .B(net604),
    .A(net669));
 sg13g2_or3_1 _3701_ (.A(_1057_),
    .B(_1058_),
    .C(net582),
    .X(_1148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3702_ (.B1(_1148_),
    .VDD(VPWR),
    .Y(_0090_),
    .VSS(VGND),
    .A1(_1522_),
    .A2(_1147_));
 sg13g2_o21ai_1 _3703_ (.B1(_0731_),
    .VDD(VPWR),
    .Y(_1149_),
    .VSS(VGND),
    .A1(_0719_),
    .A2(_0847_));
 sg13g2_and2_1 _3704_ (.A(_1063_),
    .B(_1149_),
    .X(_1150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3705_ (.Y(_1151_),
    .A(net607),
    .B(_0883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3706_ (.A(net582),
    .B(_1150_),
    .Y(_1152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3707_ (.Y(_1153_),
    .B1(_1151_),
    .B2(_1152_),
    .A2(net582),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3708_ (.VDD(VPWR),
    .Y(_0091_),
    .A(_1153_),
    .VSS(VGND));
 sg13g2_nand2b_2 _3709_ (.Y(_1154_),
    .B(_1065_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0925_));
 sg13g2_and2_1 _3710_ (.A(net611),
    .B(_0931_),
    .X(_1155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3711_ (.A(net582),
    .B(_1155_),
    .Y(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3712_ (.Y(_1157_),
    .B1(_1154_),
    .B2(_1156_),
    .A2(net582),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3713_ (.VDD(VPWR),
    .Y(_0092_),
    .A(_1157_),
    .VSS(VGND));
 sg13g2_nor2_1 _3714_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .B(_1147_),
    .Y(_1158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3715_ (.A(_1069_),
    .B(_1071_),
    .Y(_1159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3716_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1147_),
    .A2(_1159_),
    .Y(_0093_),
    .B1(_1158_));
 sg13g2_nand3b_1 _3717_ (.B(_1075_),
    .C(_0974_),
    .Y(_1160_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1074_));
 sg13g2_mux2_1 _3718_ (.A0(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .A1(_1160_),
    .S(_1147_),
    .X(_0094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3719_ (.Y(_1161_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .B(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3720_ (.B1(_1161_),
    .VDD(VPWR),
    .Y(_0095_),
    .VSS(VGND),
    .A1(_1081_),
    .A2(net582));
 sg13g2_nand3_1 _3721_ (.B(_1083_),
    .C(_1085_),
    .A(net570),
    .Y(_1162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3722_ (.A0(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .A1(_1162_),
    .S(_1147_),
    .X(_0096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3723_ (.A(_1090_),
    .B(_1092_),
    .C(net582),
    .Y(_1163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3724_ (.A2(_1146_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .B1(_1163_),
    .X(_0097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3725_ (.A(net655),
    .B(net668),
    .Y(_1164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3726_ (.Y(_1165_),
    .A(_0301_),
    .B(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3727_ (.B1(_1165_),
    .VDD(VPWR),
    .Y(_1166_),
    .VSS(VGND),
    .A1(net31),
    .A2(net603));
 sg13g2_a21oi_1 _3728_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net655),
    .A2(_1055_),
    .Y(_1167_),
    .B1(_1056_));
 sg13g2_nand3_1 _3729_ (.B(_1166_),
    .C(_1167_),
    .A(_1094_),
    .Y(_1168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3730_ (.B(_0870_),
    .C(_1168_),
    .A(net677),
    .Y(_1169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3731_ (.B1(_1169_),
    .VDD(VPWR),
    .Y(_0098_),
    .VSS(VGND),
    .A1(_1521_),
    .A2(net677));
 sg13g2_nand2b_1 _3732_ (.Y(_1170_),
    .B(net594),
    .A_N(_0894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3733_ (.Y(_1171_),
    .A(_0302_),
    .B(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3734_ (.B1(_1171_),
    .VDD(VPWR),
    .Y(_1172_),
    .VSS(VGND),
    .A1(net18),
    .A2(net602));
 sg13g2_nand2_1 _3735_ (.Y(_1173_),
    .A(net655),
    .B(_1062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3736_ (.B(_1170_),
    .C(_1172_),
    .A(_1149_),
    .Y(_1174_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1173_));
 sg13g2_a21oi_1 _3737_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net607),
    .A2(_0900_),
    .Y(_1175_),
    .B1(net655));
 sg13g2_a22oi_1 _3738_ (.Y(_1176_),
    .B1(_1174_),
    .B2(_1175_),
    .A2(net655),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3739_ (.VDD(VPWR),
    .Y(_0099_),
    .A(_1176_),
    .VSS(VGND));
 sg13g2_nand2_1 _3740_ (.Y(_1177_),
    .A(net594),
    .B(_0917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3741_ (.A(_0732_),
    .B(net603),
    .Y(_1178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3742_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1179_),
    .B(_1178_),
    .A(net11));
 sg13g2_a221oi_1 _3743_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1179_),
    .C1(net655),
    .B1(_1110_),
    .A1(net608),
    .Y(_1180_),
    .A2(_0928_));
 sg13g2_a22oi_1 _3744_ (.Y(_0100_),
    .B1(_1177_),
    .B2(_1180_),
    .A2(net655),
    .A1(_1504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3745_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .B(net678),
    .Y(_1181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3746_ (.Y(_1182_),
    .B(net595),
    .A_N(_0951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3747_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1183_),
    .B(_0945_),
    .A(net588));
 sg13g2_nand2_1 _3748_ (.Y(_1184_),
    .A(_0303_),
    .B(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3749_ (.B1(_1184_),
    .VDD(VPWR),
    .Y(_1185_),
    .VSS(VGND),
    .A1(net20),
    .A2(net603));
 sg13g2_nand4_1 _3750_ (.B(_1182_),
    .C(_1183_),
    .A(net678),
    .Y(_1186_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1185_));
 sg13g2_nor2b_1 _3751_ (.A(_1181_),
    .B_N(_1186_),
    .Y(_0101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3752_ (.A(net676),
    .B(_0969_),
    .Y(_1187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3753_ (.B1(net592),
    .VDD(VPWR),
    .Y(_1188_),
    .VSS(VGND),
    .A1(_0968_),
    .A2(_1187_));
 sg13g2_a21oi_1 _3754_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net13),
    .A2(net602),
    .Y(_1189_),
    .B1(net593));
 sg13g2_o21ai_1 _3755_ (.B1(_1189_),
    .VDD(VPWR),
    .Y(_1190_),
    .VSS(VGND),
    .A1(_1991_),
    .A2(net602));
 sg13g2_a21oi_1 _3756_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1188_),
    .A2(_1190_),
    .Y(_1191_),
    .B1(net656));
 sg13g2_a22oi_1 _3757_ (.Y(_0102_),
    .B1(_1120_),
    .B2(_1191_),
    .A2(net656),
    .A1(_1533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3758_ (.Y(_1192_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .B(net656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3759_ (.B1(net594),
    .VDD(VPWR),
    .Y(_1193_),
    .VSS(VGND),
    .A1(net676),
    .A2(_0995_));
 sg13g2_nor2_1 _3760_ (.A(_0993_),
    .B(_1193_),
    .Y(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3761_ (.A0(net569),
    .A1(_0304_),
    .S(net603),
    .X(_1195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3762_ (.Y(_1196_),
    .B(_1195_),
    .A_N(_1002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3763_ (.B1(net675),
    .VDD(VPWR),
    .Y(_1197_),
    .VSS(VGND),
    .A1(_1194_),
    .A2(_1196_));
 sg13g2_o21ai_1 _3764_ (.B1(_1192_),
    .VDD(VPWR),
    .Y(_0103_),
    .VSS(VGND),
    .A1(_1007_),
    .A2(_1197_));
 sg13g2_nand2_1 _3765_ (.Y(_1198_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .B(net656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3766_ (.B1(net592),
    .VDD(VPWR),
    .Y(_1199_),
    .VSS(VGND),
    .A1(net676),
    .A2(_1028_));
 sg13g2_nor2_1 _3767_ (.A(_1027_),
    .B(_1199_),
    .Y(_1200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3768_ (.A0(net23),
    .A1(net15),
    .S(net602),
    .X(_1201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3769_ (.A(_1140_),
    .B(_1200_),
    .C(_1201_),
    .Y(_1202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3770_ (.Y(_1203_),
    .A(net676),
    .B(_1132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3771_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1204_),
    .B(_1021_),
    .A(net586));
 sg13g2_o21ai_1 _3772_ (.B1(_1198_),
    .VDD(VPWR),
    .Y(_0104_),
    .VSS(VGND),
    .A1(_1202_),
    .A2(_1203_));
 sg13g2_nor2_1 _3773_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .B(net675),
    .Y(_1205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3774_ (.Y(_1206_),
    .A(_0306_),
    .B(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3775_ (.B1(_1206_),
    .VDD(VPWR),
    .Y(_1207_),
    .VSS(VGND),
    .A1(net24),
    .A2(net602));
 sg13g2_a21oi_1 _3776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net655),
    .A2(_1043_),
    .Y(_1208_),
    .B1(net612));
 sg13g2_nand2b_1 _3777_ (.Y(_1209_),
    .B(_1208_),
    .A_N(_1041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3778_ (.B(_1145_),
    .C(_1207_),
    .A(net675),
    .Y(_1210_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1209_));
 sg13g2_nor2b_1 _3779_ (.A(_1205_),
    .B_N(_1210_),
    .Y(_0105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3780_ (.A(net683),
    .B(net602),
    .Y(_1211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3781_ (.A(_1057_),
    .B(_1058_),
    .C(net580),
    .Y(_1212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3782_ (.A2(net580),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .B1(_1212_),
    .X(_0106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3783_ (.A(_1060_),
    .B(net580),
    .Y(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3784_ (.Y(_0107_),
    .B1(_1213_),
    .B2(_1063_),
    .A2(net580),
    .A1(_1516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3785_ (.A(_1155_),
    .B(net580),
    .Y(_1214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3786_ (.Y(_1215_),
    .B1(_1214_),
    .B2(_1154_),
    .A2(net580),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3787_ (.VDD(VPWR),
    .Y(_0108_),
    .A(_1215_),
    .VSS(VGND));
 sg13g2_nand2b_1 _3788_ (.Y(_1216_),
    .B(_1070_),
    .A_N(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3789_ (.A0(_1216_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .S(net580),
    .X(_0109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3790_ (.A0(_1160_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .S(net581),
    .X(_0110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3791_ (.Y(_1217_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .B(net581),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3792_ (.B1(_1217_),
    .VDD(VPWR),
    .Y(_0111_),
    .VSS(VGND),
    .A1(_1081_),
    .A2(net580));
 sg13g2_mux2_1 _3793_ (.A0(_1162_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .S(net581),
    .X(_0112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3794_ (.B1(net607),
    .VDD(VPWR),
    .Y(_1218_),
    .VSS(VGND),
    .A1(net683),
    .A2(_1047_));
 sg13g2_nor3_1 _3795_ (.A(net24),
    .B(_1087_),
    .C(net581),
    .Y(_1219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3796_ (.Y(_0113_),
    .B1(_1218_),
    .B2(_1219_),
    .A2(net581),
    .A1(_1547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3797_ (.A(net658),
    .B(_1057_),
    .Y(_1220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3798_ (.Y(_1221_),
    .B1(_0870_),
    .B2(_1220_),
    .A2(net657),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3799_ (.VDD(VPWR),
    .Y(_0114_),
    .A(_1221_),
    .VSS(VGND));
 sg13g2_nor2_1 _3800_ (.A(net587),
    .B(_0900_),
    .Y(_1222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3801_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net607),
    .A2(_0901_),
    .Y(_1223_),
    .B1(net657));
 sg13g2_a22oi_1 _3802_ (.Y(_0115_),
    .B1(_1063_),
    .B2(_1223_),
    .A2(net657),
    .A1(_1515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3803_ (.Y(_1224_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .B(net658),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3804_ (.Y(_1225_),
    .A(net681),
    .B(_1154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3805_ (.B1(_1224_),
    .VDD(VPWR),
    .Y(_0116_),
    .VSS(VGND),
    .A1(_0929_),
    .A2(_1225_));
 sg13g2_a21oi_1 _3806_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1070_),
    .A2(_1183_),
    .Y(_1226_),
    .B1(net658));
 sg13g2_a21o_1 _3807_ (.A2(net658),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .B1(_1226_),
    .X(_0117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3808_ (.A(net657),
    .B(_1074_),
    .Y(_1227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3809_ (.Y(_0118_),
    .B1(_1120_),
    .B2(_1227_),
    .A2(net657),
    .A1(_1532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3810_ (.Y(_1228_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .B(net658),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3811_ (.Y(_1229_),
    .A(net681),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3812_ (.B1(_1228_),
    .VDD(VPWR),
    .Y(_0119_),
    .VSS(VGND),
    .A1(_1007_),
    .A2(_1229_));
 sg13g2_nor2_1 _3813_ (.A(net657),
    .B(_1084_),
    .Y(_1230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3814_ (.Y(_0120_),
    .B1(_1204_),
    .B2(_1230_),
    .A2(net657),
    .A1(_1543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3815_ (.Y(_1231_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .B(net657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3816_ (.B1(net680),
    .VDD(VPWR),
    .Y(_1232_),
    .VSS(VGND),
    .A1(net586),
    .A2(_1045_));
 sg13g2_o21ai_1 _3817_ (.B1(_1231_),
    .VDD(VPWR),
    .Y(_0121_),
    .VSS(VGND),
    .A1(_1090_),
    .A2(_1232_));
 sg13g2_a21oi_2 _3818_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net688),
    .Y(_1233_),
    .A2(_1705_),
    .A1(_1659_));
 sg13g2_nor3_1 _3819_ (.A(_1057_),
    .B(_1058_),
    .C(net634),
    .Y(_1234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3820_ (.A2(net635),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .B1(_1234_),
    .X(_0122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3821_ (.A(_1060_),
    .B(net635),
    .Y(_1235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3822_ (.Y(_0123_),
    .B1(_1235_),
    .B2(_1063_),
    .A2(net635),
    .A1(_1514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3823_ (.A(_1066_),
    .B(net634),
    .Y(_1236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3824_ (.Y(_0124_),
    .B1(_1236_),
    .B2(_1065_),
    .A2(net635),
    .A1(_1503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3825_ (.A0(_1216_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .S(net635),
    .X(_0125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3826_ (.A0(_1160_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .S(net634),
    .X(_0126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3827_ (.B1(_1078_),
    .VDD(VPWR),
    .Y(_1237_),
    .VSS(VGND),
    .A1(net588),
    .A2(_1009_));
 sg13g2_mux2_1 _3828_ (.A0(_1237_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .S(net634),
    .X(_0127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3829_ (.Y(_1238_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .B(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3830_ (.Y(_1239_),
    .B(_1022_),
    .A_N(net686),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3831_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net610),
    .A2(_1239_),
    .Y(_1240_),
    .B1(net634));
 sg13g2_o21ai_1 _3832_ (.B1(_1240_),
    .VDD(VPWR),
    .Y(_1241_),
    .VSS(VGND),
    .A1(_1084_),
    .A2(_1140_));
 sg13g2_nand2_1 _3833_ (.Y(_0128_),
    .A(_1238_),
    .B(_1241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3834_ (.A(_1090_),
    .B(_1092_),
    .C(net634),
    .Y(_1242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3835_ (.A2(net634),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .B1(_1242_),
    .X(_0129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3836_ (.Y(_1243_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .B(net654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3837_ (.Y(_1244_),
    .A(net673),
    .B(_0870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3838_ (.B1(_0771_),
    .VDD(VPWR),
    .Y(_1245_),
    .VSS(VGND),
    .A1(_0779_),
    .A2(_0864_));
 sg13g2_nor2_1 _3839_ (.A(_0865_),
    .B(net585),
    .Y(_1246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3840_ (.Y(_1247_),
    .A(_0301_),
    .B(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3841_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0719_),
    .C1(_1055_),
    .B1(_1247_),
    .A1(_1245_),
    .Y(_1248_),
    .A2(_1246_));
 sg13g2_o21ai_1 _3842_ (.B1(_1243_),
    .VDD(VPWR),
    .Y(_0130_),
    .VSS(VGND),
    .A1(_1244_),
    .A2(_1248_));
 sg13g2_xnor2_1 _3843_ (.Y(_1249_),
    .A(_0865_),
    .B(_0891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3844_ (.A(net585),
    .B(_1249_),
    .Y(_1250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3845_ (.A(net652),
    .B(_1222_),
    .C(_1250_),
    .Y(_1251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3846_ (.Y(_0131_),
    .B1(_1251_),
    .B2(_0302_),
    .A2(net652),
    .A1(_1513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3847_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0897_),
    .A2(_0914_),
    .Y(_1252_),
    .B1(_0881_));
 sg13g2_or3_1 _3848_ (.A(net11),
    .B(_0857_),
    .C(_1064_),
    .X(_1253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3849_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0927_),
    .A2(_1252_),
    .Y(_1254_),
    .B1(_1253_));
 sg13g2_nor3_1 _3850_ (.A(_0758_),
    .B(_0929_),
    .C(_1254_),
    .Y(_1255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3851_ (.A2(net654),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .B1(_1255_),
    .X(_0132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3852_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0927_),
    .A2(_0940_),
    .Y(_1256_),
    .B1(_0881_));
 sg13g2_nand2_1 _3853_ (.Y(_1257_),
    .A(_0303_),
    .B(net673),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3854_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net572),
    .A2(_1256_),
    .Y(_1258_),
    .B1(_1257_));
 sg13g2_a22oi_1 _3855_ (.Y(_0133_),
    .B1(_1183_),
    .B2(_1258_),
    .A2(net654),
    .A1(_1498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3856_ (.A(net652),
    .B(_1119_),
    .Y(_1259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3857_ (.A(net572),
    .B(net574),
    .X(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3858_ (.A(net585),
    .B(_0977_),
    .C(_1260_),
    .Y(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3859_ (.A(net13),
    .B(_1073_),
    .C(_1261_),
    .Y(_1262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3860_ (.Y(_0134_),
    .B1(_1259_),
    .B2(_1262_),
    .A2(net652),
    .A1(_1531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3861_ (.B1(_0990_),
    .VDD(VPWR),
    .Y(_1263_),
    .VSS(VGND),
    .A1(net571),
    .A2(net573));
 sg13g2_nor2_1 _3862_ (.A(net585),
    .B(_1004_),
    .Y(_1264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3863_ (.Y(_1265_),
    .A(_0304_),
    .B(net674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3864_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1263_),
    .A2(_1264_),
    .Y(_1266_),
    .B1(_1265_));
 sg13g2_a22oi_1 _3865_ (.Y(_0135_),
    .B1(_1125_),
    .B2(_1266_),
    .A2(net653),
    .A1(_1537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3866_ (.A(_1004_),
    .B_N(_1017_),
    .Y(_1267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3867_ (.A(net585),
    .B(_1018_),
    .C(_1267_),
    .Y(_1268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3868_ (.B(net586),
    .C(_1083_),
    .A(_0305_),
    .Y(_1269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3869_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net609),
    .A2(_1021_),
    .Y(_1270_),
    .B1(net653));
 sg13g2_o21ai_1 _3870_ (.B1(_1270_),
    .VDD(VPWR),
    .Y(_1271_),
    .VSS(VGND),
    .A1(_1268_),
    .A2(_1269_));
 sg13g2_o21ai_1 _3871_ (.B1(_1271_),
    .VDD(VPWR),
    .Y(_0136_),
    .VSS(VGND),
    .A1(_1542_),
    .A2(net674));
 sg13g2_nand2_1 _3872_ (.Y(_1272_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .B(net652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3873_ (.Y(_1273_),
    .A(_1018_),
    .B(_1040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3874_ (.A(net659),
    .B(_1273_),
    .Y(_1274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3875_ (.A(net16),
    .B(net607),
    .C(_1087_),
    .D(_1274_),
    .Y(_1275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3876_ (.B1(net671),
    .VDD(VPWR),
    .Y(_1276_),
    .VSS(VGND),
    .A1(net587),
    .A2(_1045_));
 sg13g2_o21ai_1 _3877_ (.B1(_1272_),
    .VDD(VPWR),
    .Y(_0137_),
    .VSS(VGND),
    .A1(_1275_),
    .A2(_1276_));
 sg13g2_nor3_1 _3878_ (.A(net654),
    .B(_1057_),
    .C(_1058_),
    .Y(_1277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3879_ (.A2(net654),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ),
    .B1(_1277_),
    .X(_0138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3880_ (.Y(_1278_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .B(net652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3881_ (.Y(_1279_),
    .A(net671),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3882_ (.B1(_1278_),
    .VDD(VPWR),
    .Y(_0139_),
    .VSS(VGND),
    .A1(_1150_),
    .A2(_1279_));
 sg13g2_nor2_1 _3883_ (.A(net654),
    .B(_1155_),
    .Y(_1280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3884_ (.Y(_1281_),
    .B1(_1154_),
    .B2(_1280_),
    .A2(_0758_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3885_ (.VDD(VPWR),
    .Y(_0140_),
    .A(_1281_),
    .VSS(VGND));
 sg13g2_mux2_1 _3886_ (.A0(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .A1(_1216_),
    .S(net672),
    .X(_0141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3887_ (.A0(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .A1(_1160_),
    .S(net672),
    .X(_0142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3888_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .B(net672),
    .Y(_1282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3889_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net672),
    .A2(_1081_),
    .Y(_0143_),
    .B1(_1282_));
 sg13g2_nor3_1 _3890_ (.A(net653),
    .B(_1139_),
    .C(_1162_),
    .Y(_1283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3891_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1541_),
    .A2(net653),
    .Y(_0144_),
    .B1(_1283_));
 sg13g2_nor3_1 _3892_ (.A(net652),
    .B(_1090_),
    .C(_1092_),
    .Y(_1284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3893_ (.A2(net652),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .B1(_1284_),
    .X(_0145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3894_ (.Y(_1285_),
    .A(_0719_),
    .B(net648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3895_ (.VDD(VPWR),
    .Y(_1286_),
    .A(_1285_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3896_ (.B1(_1095_),
    .VDD(VPWR),
    .Y(_1287_),
    .VSS(VGND),
    .A1(_0301_),
    .A2(_1285_));
 sg13g2_nand3_1 _3897_ (.B(_0870_),
    .C(_1287_),
    .A(net649),
    .Y(_1288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3898_ (.B1(_1288_),
    .VDD(VPWR),
    .Y(_0146_),
    .VSS(VGND),
    .A1(_1520_),
    .A2(net649));
 sg13g2_nand2_1 _3899_ (.Y(_1289_),
    .A(net659),
    .B(net648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3900_ (.B1(net612),
    .VDD(VPWR),
    .Y(_1290_),
    .VSS(VGND),
    .A1(_0302_),
    .A2(_1289_));
 sg13g2_a221oi_1 _3901_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1290_),
    .C1(net643),
    .B1(_1103_),
    .A1(net607),
    .Y(_1291_),
    .A2(_0901_));
 sg13g2_a21oi_1 _3902_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1512_),
    .A2(net643),
    .Y(_0147_),
    .B1(_1291_));
 sg13g2_nand2b_1 _3903_ (.Y(_1292_),
    .B(net648),
    .A_N(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3904_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net643),
    .A2(_0931_),
    .Y(_1293_),
    .B1(net587));
 sg13g2_a221oi_1 _3905_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1293_),
    .C1(_1292_),
    .B1(_0928_),
    .A1(net595),
    .Y(_1294_),
    .A2(_0917_));
 sg13g2_a21oi_1 _3906_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1502_),
    .A2(net645),
    .Y(_0148_),
    .B1(_1294_));
 sg13g2_nor2_1 _3907_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ),
    .B(net650),
    .Y(_1295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3908_ (.B(net649),
    .C(_1182_),
    .A(_0303_),
    .Y(_1296_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1183_));
 sg13g2_nor2b_1 _3909_ (.A(_1295_),
    .B_N(_1296_),
    .Y(_0149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3910_ (.B1(net647),
    .VDD(VPWR),
    .Y(_1297_),
    .VSS(VGND),
    .A1(net586),
    .A2(_0979_));
 sg13g2_o21ai_1 _3911_ (.B1(net593),
    .VDD(VPWR),
    .Y(_1298_),
    .VSS(VGND),
    .A1(net647),
    .A2(_0969_));
 sg13g2_a21oi_1 _3912_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net13),
    .A2(_1286_),
    .Y(_1299_),
    .B1(_0975_));
 sg13g2_o21ai_1 _3913_ (.B1(_1299_),
    .VDD(VPWR),
    .Y(_1300_),
    .VSS(VGND),
    .A1(_0968_),
    .A2(_1298_));
 sg13g2_nor2b_1 _3914_ (.A(_1297_),
    .B_N(_1300_),
    .Y(_1301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3915_ (.A2(net643),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .B1(_1301_),
    .X(_0150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3916_ (.B1(net594),
    .VDD(VPWR),
    .Y(_1302_),
    .VSS(VGND),
    .A1(net647),
    .A2(_0995_));
 sg13g2_nor2_1 _3917_ (.A(_0993_),
    .B(_1302_),
    .Y(_1303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3918_ (.B1(_1001_),
    .VDD(VPWR),
    .Y(_1304_),
    .VSS(VGND),
    .A1(_0304_),
    .A2(_1285_));
 sg13g2_nor4_1 _3919_ (.A(net643),
    .B(_1124_),
    .C(_1303_),
    .D(_1304_),
    .Y(_1305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3920_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1536_),
    .A2(net643),
    .Y(_0151_),
    .B1(_1305_));
 sg13g2_o21ai_1 _3921_ (.B1(net592),
    .VDD(VPWR),
    .Y(_1306_),
    .VSS(VGND),
    .A1(net647),
    .A2(_1028_));
 sg13g2_nor2_1 _3922_ (.A(_1027_),
    .B(_1306_),
    .Y(_1307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3923_ (.A(net15),
    .B(net644),
    .Y(_1308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3924_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net570),
    .A2(net644),
    .Y(_1309_),
    .B1(_1308_));
 sg13g2_o21ai_1 _3925_ (.B1(net647),
    .VDD(VPWR),
    .Y(_1310_),
    .VSS(VGND),
    .A1(net586),
    .A2(_1021_));
 sg13g2_nor4_1 _3926_ (.A(_1139_),
    .B(_1307_),
    .C(_1309_),
    .D(_1310_),
    .Y(_1311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3927_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1540_),
    .A2(net644),
    .Y(_0152_),
    .B1(_1311_));
 sg13g2_nor3_1 _3928_ (.A(net16),
    .B(net643),
    .C(_1142_),
    .Y(_1312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3929_ (.Y(_0153_),
    .B1(_1145_),
    .B2(_1312_),
    .A2(net643),
    .A1(_1546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3930_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1313_),
    .B(\sap_3_inst.reg_file_inst.array_serializer_inst.state[1] ),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.state[0] ));
 sg13g2_inv_4 _3931_ (.A(net798),
    .Y(_0154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3932_ (.Y(_1314_),
    .B(net78),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\sap_3_inst.reg_file_inst.array_serializer_inst.state[1] ));
 sg13g2_nor2b_2 _3933_ (.A(net78),
    .B_N(\sap_3_inst.reg_file_inst.array_serializer_inst.state[1] ),
    .Y(_1315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3934_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ),
    .B(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .X(_1316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3935_ (.Y(_1317_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ),
    .B(_1316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3936_ (.Y(_1318_),
    .A(_1315_),
    .B(_1317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3937_ (.Y(_0155_),
    .A(_1314_),
    .B(_1318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3938_ (.A(net803),
    .B(_1315_),
    .Y(_1319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3939_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net803),
    .A2(_0155_),
    .Y(_0156_),
    .B1(_1319_));
 sg13g2_a21oi_1 _3940_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net803),
    .A2(_0155_),
    .Y(_1320_),
    .B1(net54));
 sg13g2_nand2_1 _3941_ (.Y(_1321_),
    .A(net61),
    .B(_1314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3942_ (.Y(_1322_),
    .A(_1315_),
    .B(_1316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3943_ (.B1(_1314_),
    .VDD(VPWR),
    .Y(_1323_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ),
    .A2(_1322_));
 sg13g2_nor2_1 _3944_ (.A(_1320_),
    .B(_1323_),
    .Y(_0157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3945_ (.Y(_0158_),
    .A(net62),
    .B(_1322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3946_ (.A2(regFile_serial_start),
    .A1(net73),
    .B1(_0154_),
    .X(_0159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3947_ (.A(net70),
    .B(_0155_),
    .Y(_1324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3948_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net803),
    .A2(_1549_),
    .Y(_1325_),
    .B1(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ));
 sg13g2_o21ai_1 _3949_ (.B1(_1325_),
    .VDD(VPWR),
    .Y(_1326_),
    .VSS(VGND),
    .A1(net803),
    .A2(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[1] ));
 sg13g2_nor2b_1 _3950_ (.A(net803),
    .B_N(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ),
    .Y(_1327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3951_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[3] ),
    .C1(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ),
    .B1(_1327_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[4] ),
    .Y(_1328_),
    .A2(_1316_));
 sg13g2_nand2_1 _3952_ (.Y(_1329_),
    .A(net803),
    .B(_1550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3953_ (.B1(_1329_),
    .VDD(VPWR),
    .Y(_1330_),
    .VSS(VGND),
    .A1(net803),
    .A2(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[5] ));
 sg13g2_o21ai_1 _3954_ (.B1(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ),
    .VDD(VPWR),
    .Y(_1331_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ),
    .A2(_1330_));
 sg13g2_a21oi_1 _3955_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[7] ),
    .A2(_1327_),
    .Y(_1332_),
    .B1(_1331_));
 sg13g2_a21oi_1 _3956_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1326_),
    .A2(_1328_),
    .Y(_1333_),
    .B1(_1332_));
 sg13g2_a22oi_1 _3957_ (.Y(_1334_),
    .B1(_1333_),
    .B2(_1315_),
    .A2(_1318_),
    .A1(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3958_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0155_),
    .A2(_1334_),
    .Y(_0160_),
    .B1(_1324_));
 sg13g2_nand2b_2 _3959_ (.Y(_1335_),
    .B(net802),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net801));
 sg13g2_nand2_2 _3960_ (.Y(_1336_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .B(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3961_ (.A(_1335_),
    .B(_1336_),
    .Y(_1337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3962_ (.A(net801),
    .B(net802),
    .C(_1336_),
    .Y(_1338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3963_ (.Y(_1339_),
    .B(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ));
 sg13g2_nor2_2 _3964_ (.A(_1335_),
    .B(_1339_),
    .Y(_1340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3965_ (.Y(_1341_),
    .B(net801),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net802));
 sg13g2_nor4_1 _3966_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .B(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .C(net801),
    .D(net802),
    .Y(_1342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3967_ (.A2(net802),
    .A1(net801),
    .B1(_1342_),
    .X(_1343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3968_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1342_),
    .Y(_1344_),
    .A2(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ));
 sg13g2_nand2b_2 _3969_ (.Y(_1345_),
    .B(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ));
 sg13g2_nor2_2 _3970_ (.A(_1341_),
    .B(_1345_),
    .Y(_1346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3971_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .B(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .C(_1335_),
    .Y(_1347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3972_ (.A(net801),
    .B(net802),
    .C(_1345_),
    .Y(_1348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3973_ (.A(net801),
    .B(net802),
    .C(_1339_),
    .Y(_1349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3974_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .B(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .C(_1341_),
    .Y(_1350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3975_ (.A(_1339_),
    .B(_1341_),
    .Y(_1351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3976_ (.A(_1335_),
    .B(_1345_),
    .Y(_1352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3977_ (.A(_1336_),
    .B(_1341_),
    .Y(_1353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3978_ (.Y(_1354_),
    .B1(_1352_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .A2(net797),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3979_ (.Y(_1355_),
    .B1(_1349_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .A2(_1347_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3980_ (.Y(_1356_),
    .B1(_1346_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ),
    .A2(_1340_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3981_ (.Y(_1357_),
    .B1(_1350_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .A2(_1348_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3982_ (.Y(_1358_),
    .B1(_1351_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ),
    .A2(net796),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3983_ (.B(_1356_),
    .C(_1357_),
    .A(_1354_),
    .Y(_1359_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1358_));
 sg13g2_a21oi_1 _3984_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .A2(_1353_),
    .Y(_1360_),
    .B1(net794));
 sg13g2_nand2_1 _3985_ (.Y(_1361_),
    .A(_1355_),
    .B(_1360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3986_ (.A(_1359_),
    .B(_1361_),
    .Y(_1362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3987_ (.B1(_0154_),
    .VDD(VPWR),
    .Y(_1363_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][0] ),
    .A2(_1344_));
 sg13g2_nand2_1 _3988_ (.Y(_1364_),
    .A(net48),
    .B(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3989_ (.B1(_1364_),
    .VDD(VPWR),
    .Y(_0161_),
    .VSS(VGND),
    .A1(_1362_),
    .A2(_1363_));
 sg13g2_a22oi_1 _3990_ (.Y(_1365_),
    .B1(_1346_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .A2(_1340_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3991_ (.Y(_1366_),
    .B1(_1351_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ),
    .A2(net796),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3992_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .A2(_1352_),
    .Y(_1367_),
    .B1(net794));
 sg13g2_a22oi_1 _3993_ (.Y(_1368_),
    .B1(_1349_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .A2(net797),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3994_ (.B(_1366_),
    .C(_1367_),
    .A(_1365_),
    .Y(_1369_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1368_));
 sg13g2_a22oi_1 _3995_ (.Y(_1370_),
    .B1(_1353_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .A2(_1347_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3996_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ),
    .C1(_1369_),
    .B1(_1350_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .Y(_1371_),
    .A2(_1348_));
 sg13g2_a221oi_1 _3997_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1371_),
    .C1(net798),
    .B1(_1370_),
    .A1(_1510_),
    .Y(_1372_),
    .A2(net794));
 sg13g2_a21o_1 _3998_ (.A2(net798),
    .A1(net66),
    .B1(_1372_),
    .X(_0162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3999_ (.Y(_1373_),
    .B1(_1348_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .A2(net797),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4000_ (.Y(_1374_),
    .B1(_1349_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .A2(net796),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4001_ (.Y(_1375_),
    .B1(_1353_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .A2(_1347_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4002_ (.Y(_1376_),
    .B1(_1352_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .A2(_1340_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4003_ (.Y(_1377_),
    .A(_1375_),
    .B(_1376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4004_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ),
    .A2(_1351_),
    .Y(_1378_),
    .B1(net795));
 sg13g2_a22oi_1 _4005_ (.Y(_1379_),
    .B1(_1350_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .A2(_1346_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4006_ (.B(_1374_),
    .C(_1378_),
    .A(_1373_),
    .Y(_1380_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1379_));
 sg13g2_a21oi_1 _4007_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1501_),
    .A2(net795),
    .Y(_1381_),
    .B1(_1313_));
 sg13g2_o21ai_1 _4008_ (.B1(_1381_),
    .VDD(VPWR),
    .Y(_1382_),
    .VSS(VGND),
    .A1(_1377_),
    .A2(_1380_));
 sg13g2_o21ai_1 _4009_ (.B1(_1382_),
    .VDD(VPWR),
    .Y(_0163_),
    .VSS(VGND),
    .A1(_1549_),
    .A2(_0154_));
 sg13g2_a22oi_1 _4010_ (.Y(_1383_),
    .B1(_1338_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .A2(_1337_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4011_ (.Y(_1384_),
    .B1(_1353_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .A2(_1347_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4012_ (.Y(_1385_),
    .B1(_1352_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .A2(_1340_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4013_ (.Y(_1386_),
    .A(_1384_),
    .B(_1385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4014_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ),
    .A2(_1351_),
    .Y(_1387_),
    .B1(net795));
 sg13g2_a22oi_1 _4015_ (.Y(_1388_),
    .B1(_1350_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .A2(_1349_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4016_ (.Y(_1389_),
    .B1(_1348_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .A2(_1346_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4017_ (.B(_1387_),
    .C(_1388_),
    .A(_1383_),
    .Y(_1390_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1389_));
 sg13g2_nor2_1 _4018_ (.A(_1386_),
    .B(_1390_),
    .Y(_1391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4019_ (.B1(_0154_),
    .VDD(VPWR),
    .Y(_1392_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][3] ),
    .A2(_1344_));
 sg13g2_nand2_1 _4020_ (.Y(_1393_),
    .A(net49),
    .B(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4021_ (.B1(_1393_),
    .VDD(VPWR),
    .Y(_0164_),
    .VSS(VGND),
    .A1(_1391_),
    .A2(_1392_));
 sg13g2_a21oi_1 _4022_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .A2(_1347_),
    .Y(_1394_),
    .B1(net794));
 sg13g2_a22oi_1 _4023_ (.Y(_1395_),
    .B1(_1340_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .A2(net796),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4024_ (.Y(_1396_),
    .B1(_1349_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .A2(_1346_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4025_ (.Y(_1397_),
    .B1(_1353_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .A2(net797),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4026_ (.Y(_1398_),
    .B1(_1351_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .A2(_1350_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4027_ (.B(_1395_),
    .C(_1397_),
    .A(_1394_),
    .Y(_1399_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1398_));
 sg13g2_a221oi_1 _4028_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .C1(_1399_),
    .B1(_1352_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .Y(_1400_),
    .A2(_1348_));
 sg13g2_o21ai_1 _4029_ (.B1(_0154_),
    .VDD(VPWR),
    .Y(_1401_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][4] ),
    .A2(_1344_));
 sg13g2_a21oi_1 _4030_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1396_),
    .A2(_1400_),
    .Y(_1402_),
    .B1(_1401_));
 sg13g2_a21o_1 _4031_ (.A2(net798),
    .A1(net63),
    .B1(_1402_),
    .X(_0165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4032_ (.Y(_1403_),
    .B1(_1351_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .A2(_1350_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4033_ (.Y(_1404_),
    .B1(_1340_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .A2(net796),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4034_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ),
    .A2(_1348_),
    .Y(_1405_),
    .B1(net795));
 sg13g2_a22oi_1 _4035_ (.Y(_1406_),
    .B1(_1353_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .A2(_1346_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4036_ (.Y(_1407_),
    .B1(_1349_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .A2(net797),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4037_ (.B(_1405_),
    .C(_1406_),
    .A(_1403_),
    .Y(_1408_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1407_));
 sg13g2_a221oi_1 _4038_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .C1(_1408_),
    .B1(_1352_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .Y(_1409_),
    .A2(_1347_));
 sg13g2_o21ai_1 _4039_ (.B1(_0154_),
    .VDD(VPWR),
    .Y(_1410_),
    .VSS(VGND),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][5] ),
    .A2(_1344_));
 sg13g2_a21oi_1 _4040_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1404_),
    .A2(_1409_),
    .Y(_1411_),
    .B1(_1410_));
 sg13g2_a21o_1 _4041_ (.A2(_1313_),
    .A1(net51),
    .B1(_1411_),
    .X(_0166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4042_ (.Y(_1412_),
    .B1(_1350_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .A2(net797),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4043_ (.Y(_1413_),
    .B1(_1353_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .A2(_1352_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4044_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ),
    .A2(_1348_),
    .Y(_1414_),
    .B1(net794));
 sg13g2_a22oi_1 _4045_ (.Y(_1415_),
    .B1(_1347_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .A2(_1340_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4046_ (.Y(_1416_),
    .B1(_1351_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ),
    .A2(_1346_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4047_ (.Y(_1417_),
    .A(_1412_),
    .B(_1416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4048_ (.Y(_1418_),
    .B1(_1349_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .A2(net796),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4049_ (.B(_1414_),
    .C(_1415_),
    .A(_1413_),
    .Y(_1419_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1418_));
 sg13g2_a21oi_1 _4050_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1539_),
    .A2(net794),
    .Y(_1420_),
    .B1(net798));
 sg13g2_o21ai_1 _4051_ (.B1(_1420_),
    .VDD(VPWR),
    .Y(_1421_),
    .VSS(VGND),
    .A1(_1417_),
    .A2(_1419_));
 sg13g2_o21ai_1 _4052_ (.B1(_1421_),
    .VDD(VPWR),
    .Y(_0167_),
    .VSS(VGND),
    .A1(_1550_),
    .A2(_0154_));
 sg13g2_a22oi_1 _4053_ (.Y(_1422_),
    .B1(_1353_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .A2(_1348_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4054_ (.Y(_1423_),
    .B1(_1340_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .A2(net797),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4055_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .A2(_1351_),
    .Y(_1424_),
    .B1(net794));
 sg13g2_a22oi_1 _4056_ (.Y(_1425_),
    .B1(_1349_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .A2(_1347_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4057_ (.Y(_1426_),
    .B1(_1352_),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .A2(_1346_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4058_ (.B(_1424_),
    .C(_1425_),
    .A(_1423_),
    .Y(_1427_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1426_));
 sg13g2_a221oi_1 _4059_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .C1(_1427_),
    .B1(_1350_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .Y(_1428_),
    .A2(net796));
 sg13g2_a221oi_1 _4060_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1428_),
    .C1(net798),
    .B1(_1422_),
    .A1(_1545_),
    .Y(_1429_),
    .A2(net794));
 sg13g2_a21o_1 _4061_ (.A2(_1313_),
    .A1(net53),
    .B1(_1429_),
    .X(_0168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4062_ (.A(net645),
    .B(_1057_),
    .C(_1058_),
    .Y(_1430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4063_ (.A2(net645),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .B1(_1430_),
    .X(_0169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4064_ (.A(net645),
    .B(_1060_),
    .Y(_1431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4065_ (.Y(_0170_),
    .B1(_1063_),
    .B2(_1431_),
    .A2(net645),
    .A1(_1511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4066_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0730_),
    .C1(net645),
    .B1(_1065_),
    .A1(net611),
    .Y(_1432_),
    .A2(_0931_));
 sg13g2_a21o_1 _4067_ (.A2(net645),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .B1(_1432_),
    .X(_0171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4068_ (.Y(_1433_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .B(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4069_ (.B1(_1433_),
    .VDD(VPWR),
    .Y(_0172_),
    .VSS(VGND),
    .A1(net646),
    .A2(_1159_));
 sg13g2_nor2_1 _4070_ (.A(net644),
    .B(_1074_),
    .Y(_1434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4071_ (.Y(_0173_),
    .B1(_1075_),
    .B2(_1434_),
    .A2(net646),
    .A1(_1530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4072_ (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .B(net650),
    .Y(_1435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4073_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net650),
    .A2(_1081_),
    .Y(_0174_),
    .B1(_1435_));
 sg13g2_mux2_1 _4074_ (.A0(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .A1(_1162_),
    .S(net647),
    .X(_0175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4075_ (.Y(_1436_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .B(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4076_ (.Y(_1437_),
    .A(net651),
    .B(_1091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4077_ (.B1(_1436_),
    .VDD(VPWR),
    .Y(_0176_),
    .VSS(VGND),
    .A1(_1090_),
    .A2(_1437_));
 sg13g2_a22oi_1 _4078_ (.Y(_1438_),
    .B1(_0321_),
    .B2(_0322_),
    .A2(net723),
    .A1(_1592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _4079_ (.Y(_1439_),
    .A(net698),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4080_ (.A(_2013_),
    .B(_2054_),
    .Y(_1440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4081_ (.A0(_1440_),
    .A1(net694),
    .S(_2002_),
    .X(_1441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4082_ (.B1(_1441_),
    .VDD(VPWR),
    .Y(_1442_),
    .VSS(VGND),
    .A1(_0331_),
    .A2(_1439_));
 sg13g2_nor2_1 _4083_ (.A(net793),
    .B(net698),
    .Y(_1443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4084_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0343_),
    .A2(net698),
    .Y(_1444_),
    .B1(_1443_));
 sg13g2_nor2_1 _4085_ (.A(net579),
    .B(_1444_),
    .Y(_1445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4086_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1525_),
    .A2(net579),
    .Y(_0177_),
    .B1(_1445_));
 sg13g2_nand2_1 _4087_ (.Y(_1446_),
    .A(_0379_),
    .B(net698),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4088_ (.B1(_1446_),
    .VDD(VPWR),
    .Y(_1447_),
    .VSS(VGND),
    .A1(net790),
    .A2(net698));
 sg13g2_nand2_1 _4089_ (.Y(_1448_),
    .A(\sap_3_inst.alu_inst.act[1] ),
    .B(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4090_ (.B1(_1448_),
    .VDD(VPWR),
    .Y(_0178_),
    .VSS(VGND),
    .A1(net579),
    .A2(_1447_));
 sg13g2_nand2b_1 _4091_ (.Y(_1449_),
    .B(net698),
    .A_N(_0412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4092_ (.B1(_1449_),
    .VDD(VPWR),
    .Y(_1450_),
    .VSS(VGND),
    .A1(net787),
    .A2(net699));
 sg13g2_nand2_1 _4093_ (.Y(_1451_),
    .A(\sap_3_inst.alu_inst.act[2] ),
    .B(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4094_ (.B1(_1451_),
    .VDD(VPWR),
    .Y(_0179_),
    .VSS(VGND),
    .A1(net578),
    .A2(_1450_));
 sg13g2_nand2b_1 _4095_ (.Y(_1452_),
    .B(net699),
    .A_N(_0444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4096_ (.B1(_1452_),
    .VDD(VPWR),
    .Y(_1453_),
    .VSS(VGND),
    .A1(net784),
    .A2(net699));
 sg13g2_nand2_1 _4097_ (.Y(_1454_),
    .A(\sap_3_inst.alu_inst.act[3] ),
    .B(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4098_ (.B1(_1454_),
    .VDD(VPWR),
    .Y(_0180_),
    .VSS(VGND),
    .A1(net578),
    .A2(_1453_));
 sg13g2_mux2_1 _4099_ (.A0(_1509_),
    .A1(_0480_),
    .S(net698),
    .X(_1455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4100_ (.Y(_1456_),
    .A(\sap_3_inst.alu_inst.act[4] ),
    .B(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4101_ (.B1(_1456_),
    .VDD(VPWR),
    .Y(_0181_),
    .VSS(VGND),
    .A1(net578),
    .A2(_1455_));
 sg13g2_nand2b_1 _4102_ (.Y(_1457_),
    .B(net699),
    .A_N(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4103_ (.B1(_1457_),
    .VDD(VPWR),
    .Y(_1458_),
    .VSS(VGND),
    .A1(net779),
    .A2(net699));
 sg13g2_nand2_1 _4104_ (.Y(_1459_),
    .A(\sap_3_inst.alu_inst.act[5] ),
    .B(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4105_ (.B1(_1459_),
    .VDD(VPWR),
    .Y(_0182_),
    .VSS(VGND),
    .A1(_1442_),
    .A2(_1458_));
 sg13g2_or2_1 _4106_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1460_),
    .B(net699),
    .A(net776));
 sg13g2_o21ai_1 _4107_ (.B1(_1460_),
    .VDD(VPWR),
    .Y(_1461_),
    .VSS(VGND),
    .A1(_0547_),
    .A2(_1439_));
 sg13g2_nand2_1 _4108_ (.Y(_1462_),
    .A(\sap_3_inst.alu_inst.act[6] ),
    .B(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4109_ (.B1(_1462_),
    .VDD(VPWR),
    .Y(_0183_),
    .VSS(VGND),
    .A1(net578),
    .A2(_1461_));
 sg13g2_nand2_1 _4110_ (.Y(_1463_),
    .A(_0578_),
    .B(net698),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4111_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net773),
    .A2(_1439_),
    .Y(_1464_),
    .B1(net579));
 sg13g2_a22oi_1 _4112_ (.Y(_0184_),
    .B1(_1463_),
    .B2(_1464_),
    .A2(net579),
    .A1(_1526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4113_ (.A(\u_ser.state[0] ),
    .B(_1489_),
    .Y(_1465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4114_ (.Y(_1466_),
    .A(\u_ser.bit_pos[1] ),
    .B(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4115_ (.Y(_1467_),
    .A(_1465_),
    .B(_1466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4116_ (.B1(_1465_),
    .VDD(VPWR),
    .Y(_1468_),
    .VSS(VGND),
    .A1(_1490_),
    .A2(_1466_));
 sg13g2_o21ai_1 _4117_ (.B1(_1468_),
    .VDD(VPWR),
    .Y(_0186_),
    .VSS(VGND),
    .A1(_1488_),
    .A2(\u_ser.state[1] ));
 sg13g2_nand3b_1 _4118_ (.B(\u_ser.shadow_reg[7] ),
    .C(\u_ser.bit_pos[1] ),
    .Y(_1469_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net800));
 sg13g2_nand2b_1 _4119_ (.Y(_1470_),
    .B(net800),
    .A_N(\u_ser.shadow_reg[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4120_ (.B1(_1470_),
    .VDD(VPWR),
    .Y(_1471_),
    .VSS(VGND),
    .A1(net800),
    .A2(\u_ser.shadow_reg[5] ));
 sg13g2_o21ai_1 _4121_ (.B1(_1469_),
    .VDD(VPWR),
    .Y(_1472_),
    .VSS(VGND),
    .A1(\u_ser.bit_pos[1] ),
    .A2(_1471_));
 sg13g2_nand3_1 _4122_ (.B(_1465_),
    .C(_1472_),
    .A(\u_ser.bit_pos[2] ),
    .Y(_1473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _4123_ (.S0(\u_ser.bit_pos[0] ),
    .A0(\u_ser.shadow_reg[1] ),
    .A1(\u_ser.shadow_reg[2] ),
    .A2(\u_ser.shadow_reg[3] ),
    .A3(\u_ser.shadow_reg[4] ),
    .S1(\u_ser.bit_pos[1] ),
    .X(_1474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4124_ (.B(_1465_),
    .C(_1474_),
    .A(_1490_),
    .Y(_1475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4125_ (.B1(\u_ser.shadow_reg[0] ),
    .VDD(VPWR),
    .Y(_1476_),
    .VSS(VGND),
    .A1(\u_ser.state[0] ),
    .A2(_1489_));
 sg13g2_nand4_1 _4126_ (.B(_1473_),
    .C(_1475_),
    .A(_0186_),
    .Y(_1477_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1476_));
 sg13g2_o21ai_1 _4127_ (.B1(_1477_),
    .VDD(VPWR),
    .Y(_1478_),
    .VSS(VGND),
    .A1(net75),
    .A2(_0186_));
 sg13g2_inv_1 _4128_ (.VDD(VPWR),
    .Y(_0187_),
    .A(_1478_),
    .VSS(VGND));
 sg13g2_a21o_1 _4129_ (.A2(net64),
    .A1(\u_ser.state[1] ),
    .B1(net799),
    .X(_0188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4130_ (.X(_1479_),
    .A(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ),
    .B(_1315_),
    .C(_1316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4131_ (.B(_1479_),
    .A(net77),
    .X(_0189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4132_ (.Y(_1480_),
    .B(_1479_),
    .A_N(_1336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4133_ (.A2(_1479_),
    .A1(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .B1(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .X(_1481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4134_ (.A(_1480_),
    .B(_1481_),
    .X(_0190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4135_ (.Y(_1482_),
    .B1(_1480_),
    .B2(net802),
    .A2(_1479_),
    .A1(net796),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4136_ (.VDD(VPWR),
    .Y(_0191_),
    .A(_1482_),
    .VSS(VGND));
 sg13g2_a22oi_1 _4137_ (.Y(_1483_),
    .B1(_1480_),
    .B2(net801),
    .A2(_1479_),
    .A1(net797),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4138_ (.VDD(VPWR),
    .Y(_0192_),
    .A(_1483_),
    .VSS(VGND));
 sg13g2_nor2_1 _4139_ (.A(net800),
    .B(_1465_),
    .Y(_1484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4140_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_0186_),
    .Y(_0193_),
    .B1(_1484_));
 sg13g2_a21oi_1 _4141_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_0186_),
    .Y(_1485_),
    .B1(net71));
 sg13g2_a21oi_1 _4142_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1467_),
    .A2(_0186_),
    .Y(_0194_),
    .B1(_1485_));
 sg13g2_nand3_1 _4143_ (.B(net800),
    .C(_1465_),
    .A(\u_ser.bit_pos[1] ),
    .Y(_1486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4144_ (.Y(_0195_),
    .B1(_1490_),
    .B2(_1486_),
    .A2(_1489_),
    .A1(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4146__4 (.VDD(VPWR),
    .Y(net38),
    .A(\clknet_leaf_1_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4147__5 (.VDD(VPWR),
    .Y(net39),
    .A(\clknet_leaf_2_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4148__6 (.VDD(VPWR),
    .Y(net40),
    .A(\clknet_leaf_0_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4149__7 (.VDD(VPWR),
    .Y(net41),
    .A(\clknet_leaf_2_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4150__8 (.VDD(VPWR),
    .Y(net42),
    .A(\clknet_leaf_2_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4151__9 (.VDD(VPWR),
    .Y(net43),
    .A(\clknet_leaf_2_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4152__10 (.VDD(VPWR),
    .Y(net44),
    .A(\clknet_leaf_0_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4153__11 (.VDD(VPWR),
    .Y(net45),
    .A(\clknet_leaf_0_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4154__12 (.VDD(VPWR),
    .Y(net46),
    .A(\clknet_leaf_0_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_inv_1 _4155__13 (.VDD(VPWR),
    .Y(net47),
    .A(\clknet_leaf_1_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_regs_0_clk_div_two (.A(\sap_3_inst.alu_inst.clk ),
    .X(\sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _4156_ (.RESET_B(net817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0017_),
    .Q(\u_ser.shadow_reg[0] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _4157_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0018_),
    .Q(\u_ser.shadow_reg[1] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4158_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0019_),
    .Q(\u_ser.shadow_reg[2] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4159_ (.RESET_B(net822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0020_),
    .Q(\u_ser.shadow_reg[3] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4160_ (.RESET_B(net822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0021_),
    .Q(\u_ser.shadow_reg[4] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4161_ (.RESET_B(net822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0022_),
    .Q(\u_ser.shadow_reg[5] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4162_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0023_),
    .Q(\u_ser.shadow_reg[6] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4163_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0024_),
    .Q(\u_ser.shadow_reg[7] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4164_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0025_),
    .Q(\sap_3_inst.alu_flags[0] ),
    .CLK(net36));
 sg13g2_dfrbpq_1 _4165_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0026_),
    .Q(\sap_3_inst.alu_flags[2] ),
    .CLK(net37));
 sg13g2_dfrbpq_1 _4166_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0027_),
    .Q(\sap_3_inst.alu_flags[3] ),
    .CLK(net38));
 sg13g2_dfrbpq_1 _4167_ (.RESET_B(net817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0028_),
    .Q(\sap_3_inst.alu_flags[1] ),
    .CLK(net39));
 sg13g2_dfrbpq_2 _4168_ (.RESET_B(net804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0001_),
    .Q(\sap_3_inst.controller_inst.stage[0] ),
    .CLK(net40));
 sg13g2_dfrbpq_2 _4169_ (.RESET_B(net807),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0002_),
    .Q(\sap_3_inst.controller_inst.stage[1] ),
    .CLK(net41));
 sg13g2_dfrbpq_2 _4170_ (.RESET_B(net807),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0003_),
    .Q(\sap_3_inst.controller_inst.stage[2] ),
    .CLK(net42));
 sg13g2_dfrbpq_1 _4171_ (.RESET_B(net807),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0004_),
    .Q(\sap_3_inst.controller_inst.stage[3] ),
    .CLK(net43));
 sg13g2_dfrbpq_1 _4172_ (.RESET_B(net805),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0029_),
    .Q(\sap_3_inst.alu_flags[4] ),
    .CLK(net44));
 sg13g2_dfrbpq_1 _4173_ (.RESET_B(net804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0030_),
    .Q(\sap_3_inst.alu_flags[5] ),
    .CLK(net45));
 sg13g2_dfrbpq_1 _4174_ (.RESET_B(net805),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0031_),
    .Q(\sap_3_inst.alu_flags[6] ),
    .CLK(net46));
 sg13g2_dfrbpq_1 _4175_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0032_),
    .Q(\sap_3_inst.alu_flags[7] ),
    .CLK(net47));
 sg13g2_dfrbpq_1 _4176_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0033_),
    .Q(\sap_3_inst.alu_inst.acc[0] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4177_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0034_),
    .Q(\sap_3_inst.alu_inst.acc[1] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4178_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0035_),
    .Q(\sap_3_inst.alu_inst.acc[2] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4179_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0036_),
    .Q(\sap_3_inst.alu_inst.acc[3] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4180_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0037_),
    .Q(\sap_3_inst.alu_inst.acc[4] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4181_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0038_),
    .Q(\sap_3_inst.alu_inst.acc[5] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4182_ (.RESET_B(net825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0039_),
    .Q(\sap_3_inst.alu_inst.acc[6] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4183_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0040_),
    .Q(\sap_3_inst.alu_inst.acc[7] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4184_ (.RESET_B(net817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0041_),
    .Q(\sap_3_inst.out[0] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4185_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0042_),
    .Q(\sap_3_inst.out[1] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4186_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0043_),
    .Q(\sap_3_inst.out[2] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4187_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0044_),
    .Q(\sap_3_inst.out[3] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4188_ (.RESET_B(net822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0045_),
    .Q(\sap_3_inst.out[4] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4189_ (.RESET_B(net822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0046_),
    .Q(\sap_3_inst.out[5] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4190_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0047_),
    .Q(\sap_3_inst.out[6] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4191_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0048_),
    .Q(\sap_3_inst.out[7] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4192_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0049_),
    .Q(\sap_3_inst.alu_inst.carry ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4193_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0050_),
    .Q(\sap_3_inst.alu_inst.tmp[0] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4194_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0051_),
    .Q(\sap_3_inst.alu_inst.tmp[1] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4195_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0052_),
    .Q(\sap_3_inst.alu_inst.tmp[2] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4196_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0053_),
    .Q(\sap_3_inst.alu_inst.tmp[3] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4197_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0054_),
    .Q(\sap_3_inst.alu_inst.tmp[4] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4198_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0055_),
    .Q(\sap_3_inst.alu_inst.tmp[5] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4199_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0056_),
    .Q(\sap_3_inst.alu_inst.tmp[6] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4200_ (.RESET_B(net817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0057_),
    .Q(\sap_3_inst.alu_inst.tmp[7] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4201_ (.RESET_B(net804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0058_),
    .Q(\sap_3_inst.controller_inst.opcode[0] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4202_ (.RESET_B(net804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0059_),
    .Q(\sap_3_inst.controller_inst.opcode[1] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4203_ (.RESET_B(net808),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0060_),
    .Q(\sap_3_inst.controller_inst.opcode[2] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4204_ (.RESET_B(net804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0061_),
    .Q(\sap_3_inst.controller_inst.opcode[3] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4205_ (.RESET_B(net804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0062_),
    .Q(\sap_3_inst.controller_inst.opcode[4] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4206_ (.RESET_B(net804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0063_),
    .Q(\sap_3_inst.controller_inst.opcode[5] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4207_ (.RESET_B(net808),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0064_),
    .Q(\sap_3_inst.controller_inst.opcode[6] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4208_ (.RESET_B(net808),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0065_),
    .Q(\sap_3_inst.controller_inst.opcode[7] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4209_ (.RESET_B(net813),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0066_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][0] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4210_ (.RESET_B(net805),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0067_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4211_ (.RESET_B(net813),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0068_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][2] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4212_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0069_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][3] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4213_ (.RESET_B(net810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0070_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][4] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4214_ (.RESET_B(net809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0071_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][5] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4215_ (.RESET_B(net810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0072_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][6] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4216_ (.RESET_B(net809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0073_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[0][7] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4217_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0074_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][0] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4218_ (.RESET_B(net808),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0075_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][1] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4219_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0076_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][2] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4220_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0077_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][3] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4221_ (.RESET_B(net815),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0078_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][4] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4222_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0079_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][5] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4223_ (.RESET_B(net811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0080_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][6] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4224_ (.RESET_B(net814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0081_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[1][7] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4225_ (.RESET_B(net816),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][0] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4226_ (.RESET_B(net805),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0083_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4227_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0084_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][2] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4228_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0085_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][3] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4229_ (.RESET_B(net810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0086_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][4] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4230_ (.RESET_B(net810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0087_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][5] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4231_ (.RESET_B(net812),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0088_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][6] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4232_ (.RESET_B(net809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0089_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[2][7] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4233_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0090_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][0] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4234_ (.RESET_B(net808),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0091_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][1] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4235_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0092_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][2] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4236_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0093_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][3] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4237_ (.RESET_B(net814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0094_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][4] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4238_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0095_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][5] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4239_ (.RESET_B(net814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0096_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][6] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4240_ (.RESET_B(net814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0097_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[3][7] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4241_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0098_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][0] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4242_ (.RESET_B(net805),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0099_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4243_ (.RESET_B(net806),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0100_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][2] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4244_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0101_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][3] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4245_ (.RESET_B(net810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0102_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][4] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4246_ (.RESET_B(net814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0103_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][5] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4247_ (.RESET_B(net812),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0104_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][6] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4248_ (.RESET_B(net809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0105_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[4][7] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4249_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0106_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][0] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4250_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0107_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][1] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4251_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0108_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][2] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4252_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0109_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][3] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4253_ (.RESET_B(net814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0110_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][4] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4254_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0111_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][5] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4255_ (.RESET_B(net811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0112_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][6] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4256_ (.RESET_B(net809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0113_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[5][7] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4257_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0114_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][0] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4258_ (.RESET_B(net804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0115_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][1] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4259_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0116_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][2] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4260_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0117_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][3] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4261_ (.RESET_B(net810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0118_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][4] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4262_ (.RESET_B(net815),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0119_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][5] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4263_ (.RESET_B(net811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0120_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][6] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4264_ (.RESET_B(net813),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0121_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[6][7] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4265_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0122_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][0] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4266_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0123_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][1] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4267_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0124_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][2] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4268_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0125_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][3] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4269_ (.RESET_B(net815),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0126_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][4] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4270_ (.RESET_B(net815),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0127_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][5] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4271_ (.RESET_B(net811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0128_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][6] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4272_ (.RESET_B(net811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0129_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[7][7] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4273_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0130_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][0] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4274_ (.RESET_B(net805),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4275_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0132_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][2] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4276_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0133_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][3] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4277_ (.RESET_B(net811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0134_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][4] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4278_ (.RESET_B(net810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0135_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][5] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4279_ (.RESET_B(net811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0136_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][6] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4280_ (.RESET_B(net809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0137_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[8][7] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4281_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0138_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][0] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4282_ (.RESET_B(net806),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0139_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][1] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4283_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0140_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][2] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4284_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0141_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][3] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4285_ (.RESET_B(net815),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0142_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][4] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4286_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0143_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][5] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4287_ (.RESET_B(net811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0144_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][6] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4288_ (.RESET_B(net814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0145_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[9][7] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4289_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0146_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][0] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4290_ (.RESET_B(net809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0147_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4291_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0148_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][2] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4292_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0149_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][3] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4293_ (.RESET_B(net810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0150_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][4] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4294_ (.RESET_B(net814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0151_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][5] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4295_ (.RESET_B(net812),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0152_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][6] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4296_ (.RESET_B(net809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0153_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[10][7] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4297_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0154_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.state[0] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _4298_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0155_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.state[1] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4299_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0156_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _4300_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net55),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _4301_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0158_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _4302_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net74),
    .Q(regFile_serial_start),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4303_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0160_),
    .Q(regFile_serial),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _4304_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0161_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[0] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4305_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0162_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[1] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4306_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0163_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[2] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4307_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0164_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[3] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _4308_ (.RESET_B(net835),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0165_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[4] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _4309_ (.RESET_B(net835),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0166_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[5] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _4310_ (.RESET_B(net835),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0167_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[6] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _4311_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0168_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[7] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _4312_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0169_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][0] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4313_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0170_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][1] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4314_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0171_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][2] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4315_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0172_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][3] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4316_ (.RESET_B(net815),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0173_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][4] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4317_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0174_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][5] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4318_ (.RESET_B(net812),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0175_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][6] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4319_ (.RESET_B(net816),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0176_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.data[11][7] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4320_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0177_),
    .Q(\sap_3_inst.alu_inst.act[0] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4321_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0178_),
    .Q(\sap_3_inst.alu_inst.act[1] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4322_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0179_),
    .Q(\sap_3_inst.alu_inst.act[2] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4323_ (.RESET_B(net825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0180_),
    .Q(\sap_3_inst.alu_inst.act[3] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4324_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0181_),
    .Q(\sap_3_inst.alu_inst.act[4] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4325_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0182_),
    .Q(\sap_3_inst.alu_inst.act[5] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4326_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0183_),
    .Q(\sap_3_inst.alu_inst.act[6] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_1 _4327_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0184_),
    .Q(\sap_3_inst.alu_inst.act[7] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs ));
 sg13g2_dfrbpq_2 _4328_ (.RESET_B(net817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net799),
    .Q(\u_ser.state[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _4329_ (.RESET_B(net817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0186_),
    .Q(\u_ser.state[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _4330_ (.RESET_B(net817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0187_),
    .Q(sap_3_outputReg_serial),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _4331_ (.RESET_B(net817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net65),
    .Q(sap_3_outputReg_start_sync),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _4332_ (.RESET_B(net835),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0189_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _4333_ (.RESET_B(net835),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0190_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[1] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _4334_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0191_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _4335_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _4336_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0193_),
    .Q(\u_ser.bit_pos[0] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _4337_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0194_),
    .Q(\u_ser.bit_pos[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _4338_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net69),
    .Q(\u_ser.bit_pos[2] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_tielo heichips25_sap3_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net34));
 sg13g2_inv_1 \clk_div_param_inst/_1__1  (.VDD(VPWR),
    .Y(net35),
    .A(clknet_1_1__leaf_clk_div_out),
    .VSS(VGND));
 sg13g2_buf_1 _4341_ (.A(mem_ram_we),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _4342_ (.A(mem_mar_we),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _4343_ (.A(sap_3_outputReg_serial),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _4344_ (.A(sap_3_outputReg_start_sync),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 _4345_ (.A(regFile_serial),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 _4346_ (.A(regFile_serial_start),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2133__2 (.VDD(VPWR),
    .Y(net36),
    .A(\clknet_leaf_1_sap_3_inst.alu_inst.clk ),
    .VSS(VGND));
 sg13g2_dfrbpq_1 \clk_div_param_inst/_2_  (.RESET_B(net808),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net35),
    .Q(clk_div_out),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_lgcp_1 \sap_3_inst.clock.clock_gate_inst  (.GATE(_0000_),
    .CLK(clknet_1_0__leaf_clk_div_out),
    .GCLK(\sap_3_inst.alu_inst.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout569 (.A(_1967_),
    .X(net569),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout570 (.A(_1941_),
    .X(net570),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout571 (.A(net572),
    .X(net571),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout572 (.A(_0943_),
    .X(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout573 (.A(_0967_),
    .X(net573),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout574 (.A(_0967_),
    .X(net574),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout575 (.A(_0354_),
    .X(net575),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout576 (.A(_1721_),
    .X(net576),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout577 (.A(_1721_),
    .X(net577),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout578 (.A(net579),
    .X(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout579 (.A(_1442_),
    .X(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout580 (.A(net581),
    .X(net580),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout581 (.A(_1211_),
    .X(net581),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout582 (.A(_1146_),
    .X(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout583 (.A(_1053_),
    .X(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout584 (.A(_1053_),
    .X(net584),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout585 (.A(_0881_),
    .X(net585),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout586 (.A(net587),
    .X(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout587 (.A(net588),
    .X(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout588 (.A(_0858_),
    .X(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout589 (.A(net591),
    .X(net589),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout590 (.A(net591),
    .X(net590),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout591 (.A(_0825_),
    .X(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout592 (.A(net593),
    .X(net592),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout594 (.A(net595),
    .X(net594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout595 (.A(_0744_),
    .X(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout596 (.A(net597),
    .X(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout597 (.A(_0741_),
    .X(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout599 (.A(_0340_),
    .X(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout600 (.A(_1862_),
    .X(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout601 (.A(_1850_),
    .X(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout602 (.A(net603),
    .X(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout603 (.A(_1164_),
    .X(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout604 (.A(_1096_),
    .X(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout605 (.A(net606),
    .X(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout606 (.A(_0876_),
    .X(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout607 (.A(net608),
    .X(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout608 (.A(net611),
    .X(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout609 (.A(net610),
    .X(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout610 (.A(net611),
    .X(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout611 (.A(_0857_),
    .X(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout612 (.A(_0745_),
    .X(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout613 (.A(_0745_),
    .X(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout614 (.A(net615),
    .X(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout615 (.A(_1864_),
    .X(net615),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout616 (.A(net617),
    .X(net616),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout617 (.A(_1860_),
    .X(net617),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout618 (.A(net619),
    .X(net618),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout619 (.A(_1859_),
    .X(net619),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout620 (.A(_1856_),
    .X(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout621 (.A(_1856_),
    .X(net621),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout622 (.A(net623),
    .X(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout623 (.A(_1853_),
    .X(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout624 (.A(_1852_),
    .X(net624),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout625 (.A(_1852_),
    .X(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout626 (.A(net627),
    .X(net626),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout627 (.A(_1849_),
    .X(net627),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout628 (.A(net629),
    .X(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout629 (.A(_1847_),
    .X(net629),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout630 (.A(net633),
    .X(net630),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout631 (.A(net632),
    .X(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout632 (.A(net633),
    .X(net632),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout633 (.A(_1845_),
    .X(net633),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout634 (.A(_1233_),
    .X(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout635 (.A(_1233_),
    .X(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout636 (.A(net637),
    .X(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout637 (.A(_0766_),
    .X(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout638 (.A(net640),
    .X(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout639 (.A(net640),
    .X(net639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout640 (.A(_0765_),
    .X(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout641 (.A(_0762_),
    .X(net641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout642 (.A(_0762_),
    .X(net642),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout643 (.A(net646),
    .X(net643),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout644 (.A(net646),
    .X(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout645 (.A(net646),
    .X(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout646 (.A(_0760_),
    .X(net646),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout647 (.A(net648),
    .X(net647),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout648 (.A(net651),
    .X(net648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout649 (.A(net651),
    .X(net649),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout650 (.A(net651),
    .X(net650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout651 (.A(_0759_),
    .X(net651),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout652 (.A(net654),
    .X(net652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout653 (.A(net654),
    .X(net653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout654 (.A(_0758_),
    .X(net654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout655 (.A(_0754_),
    .X(net655),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout656 (.A(_0754_),
    .X(net656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout657 (.A(_0751_),
    .X(net657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout658 (.A(_0751_),
    .X(net658),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout659 (.A(_0730_),
    .X(net659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout660 (.A(net661),
    .X(net660),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout661 (.A(net662),
    .X(net661),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout662 (.A(_0713_),
    .X(net662),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout663 (.A(net664),
    .X(net663),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout664 (.A(net665),
    .X(net664),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout665 (.A(_0712_),
    .X(net665),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout666 (.A(_1828_),
    .X(net666),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout667 (.A(_1809_),
    .X(net667),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout668 (.A(_0874_),
    .X(net668),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout669 (.A(net670),
    .X(net669),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout670 (.A(_0763_),
    .X(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout671 (.A(net674),
    .X(net671),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout672 (.A(net673),
    .X(net672),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout673 (.A(net674),
    .X(net673),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout674 (.A(_0757_),
    .X(net674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout675 (.A(net679),
    .X(net675),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout676 (.A(net679),
    .X(net676),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout677 (.A(net679),
    .X(net677),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout678 (.A(net679),
    .X(net678),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout679 (.A(_0753_),
    .X(net679),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout680 (.A(net682),
    .X(net680),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout681 (.A(net682),
    .X(net681),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout682 (.A(_0750_),
    .X(net682),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout683 (.A(net685),
    .X(net683),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout684 (.A(net685),
    .X(net684),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout685 (.A(_0747_),
    .X(net685),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout686 (.A(net688),
    .X(net686),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout687 (.A(net688),
    .X(net687),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout688 (.A(_0711_),
    .X(net688),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout689 (.A(_0709_),
    .X(net689),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout690 (.A(_0709_),
    .X(net690),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout691 (.A(_0359_),
    .X(net691),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout692 (.A(_0357_),
    .X(net692),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout693 (.A(_0330_),
    .X(net693),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout694 (.A(_0330_),
    .X(net694),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout695 (.A(_1899_),
    .X(net695),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout696 (.A(_1792_),
    .X(net696),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout697 (.A(_1792_),
    .X(net697),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout698 (.A(_1438_),
    .X(net698),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout699 (.A(_1438_),
    .X(net699),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout700 (.A(net701),
    .X(net700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout701 (.A(_0615_),
    .X(net701),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout702 (.A(net703),
    .X(net702),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout703 (.A(_0320_),
    .X(net703),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout704 (.A(_2000_),
    .X(net704),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout705 (.A(_0274_),
    .X(net705),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout706 (.A(_0274_),
    .X(net706),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout707 (.A(_1830_),
    .X(net707),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout708 (.A(net709),
    .X(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout709 (.A(_2014_),
    .X(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout710 (.A(_1915_),
    .X(net710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout711 (.A(net713),
    .X(net711),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout712 (.A(net713),
    .X(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout713 (.A(_1796_),
    .X(net713),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout714 (.A(net715),
    .X(net714),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout715 (.A(_1664_),
    .X(net715),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout716 (.A(_1601_),
    .X(net716),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout717 (.A(net718),
    .X(net717),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout718 (.A(_1585_),
    .X(net718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout719 (.A(_1760_),
    .X(net719),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout720 (.A(_1752_),
    .X(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout721 (.A(_1723_),
    .X(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout722 (.A(_1722_),
    .X(net722),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout723 (.A(_1722_),
    .X(net723),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout724 (.A(_1631_),
    .X(net724),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout725 (.A(_1613_),
    .X(net725),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout726 (.A(net727),
    .X(net726),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout727 (.A(_1583_),
    .X(net727),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout728 (.A(net729),
    .X(net728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout729 (.A(_1583_),
    .X(net729),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout730 (.A(_1582_),
    .X(net730),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout731 (.A(_1582_),
    .X(net731),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout732 (.A(_1671_),
    .X(net732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout733 (.A(_1662_),
    .X(net733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout734 (.A(_1661_),
    .X(net734),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout735 (.A(_1652_),
    .X(net735),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout736 (.A(_1610_),
    .X(net736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout737 (.A(_1586_),
    .X(net737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout738 (.A(_1584_),
    .X(net738),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout739 (.A(_1568_),
    .X(net739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout740 (.A(_1567_),
    .X(net740),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout741 (.A(_1566_),
    .X(net741),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout742 (.A(_1566_),
    .X(net742),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout743 (.A(_1551_),
    .X(net743),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout744 (.A(\sap_3_inst.controller_inst.stage[3] ),
    .X(net744),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout745 (.A(\sap_3_inst.controller_inst.stage[2] ),
    .X(net745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout746 (.A(\sap_3_inst.controller_inst.stage[1] ),
    .X(net746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout747 (.A(\sap_3_inst.controller_inst.stage[0] ),
    .X(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout748 (.A(\sap_3_inst.alu_flags[1] ),
    .X(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout749 (.A(_1625_),
    .X(net749),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout750 (.A(_1565_),
    .X(net750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout751 (.A(_1563_),
    .X(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout752 (.A(_1558_),
    .X(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout753 (.A(net754),
    .X(net753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout754 (.A(\sap_3_inst.controller_inst.opcode[7] ),
    .X(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout755 (.A(net756),
    .X(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout756 (.A(\sap_3_inst.controller_inst.opcode[6] ),
    .X(net756),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout757 (.A(net758),
    .X(net757),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout758 (.A(\sap_3_inst.controller_inst.opcode[5] ),
    .X(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout759 (.A(net761),
    .X(net759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout760 (.A(net761),
    .X(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout761 (.A(\sap_3_inst.controller_inst.opcode[4] ),
    .X(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout762 (.A(net763),
    .X(net762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout763 (.A(\sap_3_inst.controller_inst.opcode[3] ),
    .X(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout764 (.A(\sap_3_inst.controller_inst.opcode[3] ),
    .X(net764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout765 (.A(\sap_3_inst.controller_inst.opcode[2] ),
    .X(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout766 (.A(\sap_3_inst.controller_inst.opcode[2] ),
    .X(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout767 (.A(net768),
    .X(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout768 (.A(net769),
    .X(net768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout769 (.A(\sap_3_inst.controller_inst.opcode[1] ),
    .X(net769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout770 (.A(net771),
    .X(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout771 (.A(\sap_3_inst.controller_inst.opcode[0] ),
    .X(net771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout772 (.A(net773),
    .X(net772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout773 (.A(net774),
    .X(net773),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout774 (.A(\sap_3_inst.alu_inst.acc[7] ),
    .X(net774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout775 (.A(net776),
    .X(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout776 (.A(net777),
    .X(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout777 (.A(\sap_3_inst.alu_inst.acc[6] ),
    .X(net777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout778 (.A(net779),
    .X(net778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout779 (.A(net780),
    .X(net779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout780 (.A(\sap_3_inst.alu_inst.acc[5] ),
    .X(net780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout781 (.A(net782),
    .X(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout782 (.A(\sap_3_inst.alu_inst.acc[4] ),
    .X(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout783 (.A(net785),
    .X(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout784 (.A(net785),
    .X(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout785 (.A(\sap_3_inst.alu_inst.acc[3] ),
    .X(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout786 (.A(net788),
    .X(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout787 (.A(net788),
    .X(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout788 (.A(\sap_3_inst.alu_inst.acc[2] ),
    .X(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout789 (.A(net791),
    .X(net789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout790 (.A(net791),
    .X(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout791 (.A(\sap_3_inst.alu_inst.acc[1] ),
    .X(net791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout792 (.A(net793),
    .X(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout793 (.A(\sap_3_inst.alu_inst.acc[0] ),
    .X(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout794 (.A(_1343_),
    .X(net794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout795 (.A(_1343_),
    .X(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout796 (.A(_1338_),
    .X(net796),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout797 (.A(_1337_),
    .X(net797),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout798 (.A(_1313_),
    .X(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout799 (.A(_0185_),
    .X(net799),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout800 (.A(\u_ser.bit_pos[0] ),
    .X(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout801 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[3] ),
    .X(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout802 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[2] ),
    .X(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout803 (.A(net79),
    .X(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout804 (.A(net806),
    .X(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout805 (.A(net806),
    .X(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout806 (.A(net807),
    .X(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout807 (.A(net808),
    .X(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout808 (.A(net836),
    .X(net808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout809 (.A(net813),
    .X(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout810 (.A(net812),
    .X(net810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout811 (.A(net812),
    .X(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout812 (.A(net813),
    .X(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout813 (.A(net836),
    .X(net813),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout814 (.A(net816),
    .X(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout815 (.A(net816),
    .X(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout816 (.A(net836),
    .X(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout817 (.A(net818),
    .X(net817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout818 (.A(net826),
    .X(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout819 (.A(net826),
    .X(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout820 (.A(net826),
    .X(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout821 (.A(net825),
    .X(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout822 (.A(net825),
    .X(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout823 (.A(net825),
    .X(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout824 (.A(net825),
    .X(net824),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout825 (.A(net826),
    .X(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout826 (.A(net836),
    .X(net826),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout827 (.A(net829),
    .X(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout828 (.A(net832),
    .X(net828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout829 (.A(net832),
    .X(net829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout830 (.A(net832),
    .X(net830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout831 (.A(net832),
    .X(net831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout832 (.A(net836),
    .X(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout833 (.A(net834),
    .X(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout834 (.A(net835),
    .X(net834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout835 (.A(net836),
    .X(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout836 (.A(rst_n),
    .X(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net31),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net32),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout31 (.A(net17),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout32 (.A(net20),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_sap3_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net33));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload0 (.VDD(VPWR),
    .A(clknet_3_1__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_1 clkload1 (.A(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload2 (.VDD(VPWR),
    .A(clknet_3_3__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload4 (.VDD(VPWR),
    .A(clknet_3_5__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload5 (.VDD(VPWR),
    .A(clknet_3_6__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload6 (.VDD(VPWR),
    .A(clknet_3_7__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk_div_out (.A(clk_div_out),
    .X(clknet_0_clk_div_out),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_clk_div_out (.A(clknet_0_clk_div_out),
    .X(clknet_1_0__leaf_clk_div_out),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_1__f_clk_div_out (.A(clknet_0_clk_div_out),
    .X(clknet_1_1__leaf_clk_div_out),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload7 (.A(clknet_1_1__leaf_clk_div_out),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_leaf_0_sap_3_inst.alu_inst.clk  (.A(\clknet_1_0__leaf_sap_3_inst.alu_inst.clk ),
    .X(\clknet_leaf_0_sap_3_inst.alu_inst.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_leaf_1_sap_3_inst.alu_inst.clk  (.A(\clknet_1_1__leaf_sap_3_inst.alu_inst.clk ),
    .X(\clknet_leaf_1_sap_3_inst.alu_inst.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_leaf_2_sap_3_inst.alu_inst.clk  (.A(\clknet_1_0__leaf_sap_3_inst.alu_inst.clk ),
    .X(\clknet_leaf_2_sap_3_inst.alu_inst.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_0_sap_3_inst.alu_inst.clk  (.A(\sap_3_inst.alu_inst.clk ),
    .X(\clknet_0_sap_3_inst.alu_inst.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_1_0__f_sap_3_inst.alu_inst.clk  (.A(\clknet_0_sap_3_inst.alu_inst.clk ),
    .X(\clknet_1_0__leaf_sap_3_inst.alu_inst.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_1_1__f_sap_3_inst.alu_inst.clk  (.A(\clknet_0_sap_3_inst.alu_inst.clk ),
    .X(\clknet_1_1__leaf_sap_3_inst.alu_inst.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload8 (.A(\clknet_1_1__leaf_sap_3_inst.alu_inst.clk ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_0_sap_3_inst.alu_inst.clk_regs  (.A(\sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_0_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_0_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_1_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_1_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_2_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_2_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_3_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_3_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_4_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_4_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_5_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_5_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_6_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_6_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_7_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_7_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_8_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_8_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_9_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_9_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_10_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_10_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_11_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_11_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_12_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_12_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_13_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_13_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_14_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_14_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_4_15_0_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_4_15_0_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_0__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_0_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_0__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_1__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_0_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_2__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_1_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_2__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_3__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_1_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_4__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_2_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_4__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_5__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_2_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_6__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_3_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_7__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_3_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_7__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_8__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_4_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_8__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_9__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_4_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_10__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_5_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_10__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_11__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_5_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_12__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_6_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_12__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_13__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_6_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_14__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_7_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_14__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_15__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_7_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_15__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_16__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_8_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_16__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_17__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_8_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_18__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_9_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_18__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_19__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_9_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_19__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_20__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_10_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_20__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_21__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_10_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_22__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_11_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_22__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_23__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_11_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_24__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_12_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_24__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_25__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_12_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_26__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_13_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_26__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_27__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_13_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_27__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_28__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_14_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_28__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_29__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_14_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_30__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_15_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_30__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 \clkbuf_5_31__f_sap_3_inst.alu_inst.clk_regs  (.A(\clknet_4_15_0_sap_3_inst.alu_inst.clk_regs ),
    .X(\clknet_5_31__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload9 (.VDD(VPWR),
    .A(\clknet_5_1__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload10 (.VDD(VPWR),
    .A(\clknet_5_3__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload11 (.VDD(VPWR),
    .A(\clknet_5_5__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VSS(VGND));
 sg13g2_buf_1 clkload12 (.A(\clknet_5_6__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload13 (.VDD(VPWR),
    .A(\clknet_5_9__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VSS(VGND));
 sg13g2_buf_1 clkload14 (.A(\clknet_5_11__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload15 (.VDD(VPWR),
    .A(\clknet_5_13__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload16 (.VDD(VPWR),
    .A(\clknet_5_17__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload17 (.VDD(VPWR),
    .A(\clknet_5_21__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VSS(VGND));
 sg13g2_buf_1 clkload18 (.A(\clknet_5_23__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload19 (.VDD(VPWR),
    .A(\clknet_5_25__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VSS(VGND));
 sg13g2_inv_1 clkload20 (.VDD(VPWR),
    .A(\clknet_5_29__leaf_sap_3_inst.alu_inst.clk_regs ),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold2 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold3 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold4 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold5 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold6 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold7 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0157_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_ser.shadow_reg[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_ser.shadow_reg[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_ser.shadow_reg[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_ser.shadow_reg[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_ser.shadow_reg[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold14 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold15 (.A(_1321_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold16 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold17 (.A(sap_3_outputReg_start_sync),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0188_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold19 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.shadow_reg[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold20 (.A(\u_ser.shadow_reg[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_ser.state[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0195_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold23 (.A(regFile_serial),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u_ser.bit_pos[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_ser.shadow_reg[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold26 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.state[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0159_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold28 (.A(sap_3_outputReg_serial),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_ser.shadow_reg[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold30 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.word_index[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold31 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.state[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold32 (.A(\sap_3_inst.reg_file_inst.array_serializer_inst.bit_pos[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net79));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uo_out[6] = net33;
 assign uo_out[7] = net34;
endmodule
