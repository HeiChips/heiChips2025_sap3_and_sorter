* NGSPICE file created from heichips25_top_sorter.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

.subckt heichips25_top_sorter VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_277 VPWR VGND sg13g2_fill_2
XFILLER_36_951 VPWR VGND sg13g2_decap_8
XFILLER_35_1009 VPWR VGND sg13g2_decap_8
X_6776_ net189 VGND VPWR _0286_ s0.genblk1\[9\].modules.bubble clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
XFILLER_23_678 VPWR VGND sg13g2_decap_8
X_3988_ _1547_ VPWR _1548_ VGND net1490 net618 sg13g2_o21ai_1
X_5727_ _0317_ VPWR _0318_ VGND net1012 _0316_ sg13g2_o21ai_1
XFILLER_10_328 VPWR VGND sg13g2_decap_8
X_5658_ _3052_ net1308 net527 VPWR VGND sg13g2_nand2_1
X_5589_ net1325 VPWR _2992_ VGND _2909_ _2991_ sg13g2_o21ai_1
X_4609_ VGND VPWR net997 _2047_ _2105_ net1370 sg13g2_a21oi_1
Xhold351 _0196_ VPWR VGND net671 sg13g2_dlygate4sd3_1
Xhold340 s0.data_out\[18\]\[0\] VPWR VGND net660 sg13g2_dlygate4sd3_1
Xhold362 s0.data_out\[6\]\[2\] VPWR VGND net682 sg13g2_dlygate4sd3_1
Xhold373 s0.data_out\[15\]\[6\] VPWR VGND net693 sg13g2_dlygate4sd3_1
Xhold384 s0.data_new_delayed\[4\] VPWR VGND net704 sg13g2_dlygate4sd3_1
XFILLER_19_918 VPWR VGND sg13g2_decap_8
XFILLER_26_461 VPWR VGND sg13g2_fill_2
XFILLER_42_943 VPWR VGND sg13g2_decap_8
XFILLER_9_104 VPWR VGND sg13g2_decap_8
XFILLER_14_689 VPWR VGND sg13g2_fill_2
XFILLER_49_520 VPWR VGND sg13g2_decap_8
XFILLER_1_582 VPWR VGND sg13g2_decap_8
XFILLER_49_597 VPWR VGND sg13g2_decap_8
XFILLER_36_269 VPWR VGND sg13g2_fill_2
XFILLER_18_973 VPWR VGND sg13g2_decap_8
XFILLER_33_921 VPWR VGND sg13g2_fill_2
X_4960_ net1037 net1157 _2423_ VPWR VGND sg13g2_nor2b_1
XFILLER_44_280 VPWR VGND sg13g2_fill_1
X_4891_ _2356_ VPWR _2357_ VGND net1051 _2242_ sg13g2_o21ai_1
X_3911_ _1477_ net1177 net477 VPWR VGND sg13g2_nand2_1
XFILLER_33_965 VPWR VGND sg13g2_decap_8
X_3842_ _1419_ VPWR _1420_ VGND net1484 net621 sg13g2_o21ai_1
X_6630_ net208 VGND VPWR _0140_ s0.data_out\[12\]\[4\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_6561_ net283 VGND VPWR _0071_ s0.data_out\[18\]\[6\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_5512_ _2916_ net1315 _2917_ _2918_ VPWR VGND sg13g2_a21o_1
X_3773_ _1352_ net1190 net422 VPWR VGND sg13g2_nand2_1
X_6492_ net61 VGND VPWR _0002_ s0.valid_out\[23\][0] clknet_leaf_0_clk sg13g2_dfrbpq_2
X_5443_ VPWR _2861_ net578 VGND sg13g2_inv_1
X_5374_ VPWR _2792_ net352 VGND sg13g2_inv_1
X_4325_ VGND VPWR _1848_ _1839_ net1412 sg13g2_or2_1
XFILLER_47_18 VPWR VGND sg13g2_decap_8
X_4256_ VPWR _0185_ _1784_ VGND sg13g2_inv_1
X_4187_ _1720_ net1116 _1721_ _1722_ VPWR VGND sg13g2_a21o_1
X_6680__154 VPWR VGND net154 sg13g2_tiehi
XFILLER_27_203 VPWR VGND sg13g2_decap_8
XFILLER_43_718 VPWR VGND sg13g2_fill_1
XFILLER_43_707 VPWR VGND sg13g2_decap_4
XFILLER_43_729 VPWR VGND sg13g2_fill_2
XFILLER_42_217 VPWR VGND sg13g2_fill_2
XFILLER_24_932 VPWR VGND sg13g2_decap_4
XFILLER_11_604 VPWR VGND sg13g2_decap_8
XFILLER_23_453 VPWR VGND sg13g2_decap_4
XFILLER_24_998 VPWR VGND sg13g2_decap_8
XFILLER_10_125 VPWR VGND sg13g2_fill_1
XFILLER_10_114 VPWR VGND sg13g2_fill_1
X_6759_ net69 VGND VPWR _0269_ s0.data_out\[2\]\[5\] clknet_leaf_9_clk sg13g2_dfrbpq_2
XFILLER_7_619 VPWR VGND sg13g2_decap_8
XFILLER_6_129 VPWR VGND sg13g2_fill_1
XFILLER_3_803 VPWR VGND sg13g2_decap_8
XFILLER_12_65 VPWR VGND sg13g2_decap_8
XFILLER_2_324 VPWR VGND sg13g2_fill_2
Xhold170 _0169_ VPWR VGND net490 sg13g2_dlygate4sd3_1
Xhold192 s0.data_out\[2\]\[7\] VPWR VGND net512 sg13g2_dlygate4sd3_1
Xhold181 s0.data_out\[6\]\[1\] VPWR VGND net501 sg13g2_dlygate4sd3_1
XFILLER_19_704 VPWR VGND sg13g2_decap_4
XFILLER_37_40 VPWR VGND sg13g2_fill_2
XFILLER_18_225 VPWR VGND sg13g2_fill_2
XFILLER_19_737 VPWR VGND sg13g2_decap_8
XFILLER_18_236 VPWR VGND sg13g2_decap_8
XFILLER_15_921 VPWR VGND sg13g2_fill_2
XFILLER_18_1015 VPWR VGND sg13g2_decap_8
XFILLER_30_935 VPWR VGND sg13g2_fill_1
XFILLER_30_968 VPWR VGND sg13g2_decap_8
X_6508__44 VPWR VGND net44 sg13g2_tiehi
XFILLER_5_140 VPWR VGND sg13g2_fill_1
XFILLER_10_692 VPWR VGND sg13g2_fill_2
X_5090_ _2535_ VPWR _2541_ VGND _2528_ _2538_ sg13g2_o21ai_1
XFILLER_25_1008 VPWR VGND sg13g2_decap_8
X_4110_ net1385 _1573_ _1655_ VPWR VGND sg13g2_nor2_1
X_4041_ _1588_ net1014 _1587_ VPWR VGND sg13g2_nand2_1
X_5992_ VGND VPWR net1003 _0445_ _0556_ _0555_ sg13g2_a21oi_1
X_4943_ _2406_ net580 net1058 VPWR VGND sg13g2_nand2b_1
XFILLER_24_239 VPWR VGND sg13g2_fill_1
XFILLER_21_957 VPWR VGND sg13g2_decap_8
X_6613_ net226 VGND VPWR _0123_ s0.genblk1\[12\].modules.bubble clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_4874_ VPWR _0244_ _2343_ VGND sg13g2_inv_1
X_3825_ s0.data_out\[11\]\[5\] s0.data_out\[12\]\[5\] net1199 _1404_ VPWR VGND sg13g2_mux2_1
X_6544_ net301 VGND VPWR net696 s0.data_out\[19\]\[1\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3756_ net1485 VPWR _1337_ VGND _1334_ _1336_ sg13g2_o21ai_1
X_6475_ net1241 VPWR _0992_ VGND _0934_ _0991_ sg13g2_o21ai_1
X_5426_ VPWR _2844_ net589 VGND sg13g2_inv_1
X_3687_ net1194 net1154 _1277_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_817 VPWR VGND sg13g2_decap_8
X_5357_ VPWR _2775_ net640 VGND sg13g2_inv_1
X_5288_ net361 net1025 net1023 _2715_ VPWR VGND sg13g2_a21o_1
X_4308_ _1831_ _1830_ net1441 _1806_ net1446 VPWR VGND sg13g2_a22oi_1
X_4239_ net1000 _2852_ _1771_ VPWR VGND sg13g2_nor2_1
XFILLER_15_228 VPWR VGND sg13g2_decap_8
XFILLER_24_740 VPWR VGND sg13g2_fill_2
XFILLER_12_913 VPWR VGND sg13g2_decap_8
XFILLER_11_434 VPWR VGND sg13g2_fill_2
XFILLER_11_456 VPWR VGND sg13g2_decap_8
XFILLER_12_968 VPWR VGND sg13g2_decap_8
XFILLER_20_990 VPWR VGND sg13g2_decap_8
XFILLER_3_600 VPWR VGND sg13g2_fill_1
X_6505__47 VPWR VGND net47 sg13g2_tiehi
XFILLER_48_1019 VPWR VGND sg13g2_decap_8
X_6728__102 VPWR VGND net102 sg13g2_tiehi
XFILLER_3_677 VPWR VGND sg13g2_decap_8
XFILLER_2_132 VPWR VGND sg13g2_fill_1
Xfanout1412 net1415 net1412 VPWR VGND sg13g2_buf_1
XFILLER_2_176 VPWR VGND sg13g2_fill_1
Xfanout1401 ui_in[7] net1401 VPWR VGND sg13g2_buf_8
Xfanout1423 net1425 net1423 VPWR VGND sg13g2_buf_8
Xfanout1434 ui_in[4] net1434 VPWR VGND sg13g2_buf_8
Xfanout1445 net1446 net1445 VPWR VGND sg13g2_buf_8
Xfanout1456 net1457 net1456 VPWR VGND sg13g2_buf_8
XFILLER_48_94 VPWR VGND sg13g2_fill_2
XFILLER_48_83 VPWR VGND sg13g2_decap_8
Xfanout1489 net1492 net1489 VPWR VGND sg13g2_buf_1
Xfanout1467 net1469 net1467 VPWR VGND sg13g2_buf_8
Xfanout1478 net1483 net1478 VPWR VGND sg13g2_buf_8
XFILLER_47_843 VPWR VGND sg13g2_decap_8
XFILLER_0_79 VPWR VGND sg13g2_fill_1
XFILLER_21_209 VPWR VGND sg13g2_fill_1
X_4590_ VGND VPWR _2077_ _2079_ _2089_ net1430 sg13g2_a21oi_1
X_3610_ VPWR _0117_ net523 VGND sg13g2_inv_1
XFILLER_11_990 VPWR VGND sg13g2_decap_8
X_3541_ _1143_ net532 net1220 VPWR VGND sg13g2_nand2b_1
X_3472_ net1227 VPWR _1084_ VGND _1012_ _1083_ sg13g2_o21ai_1
X_6260_ net1238 net1172 _0797_ VPWR VGND sg13g2_nor2b_1
X_5211_ _2643_ VPWR _2650_ VGND _2644_ _2646_ sg13g2_o21ai_1
X_6191_ _0737_ _0738_ _0739_ _0740_ VPWR VGND sg13g2_nor3_1
X_5142_ net1346 _2577_ _0273_ VPWR VGND sg13g2_nor2_1
XFILLER_9_1024 VPWR VGND sg13g2_decap_4
XFILLER_29_0 VPWR VGND sg13g2_fill_2
XFILLER_38_821 VPWR VGND sg13g2_fill_1
X_5073_ VGND VPWR net1028 _2523_ _2524_ _2522_ sg13g2_a21oi_1
X_4024_ _1569_ net1124 _1570_ _1571_ VPWR VGND sg13g2_a21o_1
XFILLER_40_507 VPWR VGND sg13g2_fill_2
X_5975_ net1352 _0510_ _0543_ VPWR VGND sg13g2_nor2_1
XFILLER_21_721 VPWR VGND sg13g2_fill_1
X_4926_ net1037 net993 _2389_ VPWR VGND sg13g2_nor2_1
XFILLER_20_231 VPWR VGND sg13g2_fill_2
X_4857_ VPWR _0240_ _2330_ VGND sg13g2_inv_1
X_3808_ VGND VPWR net1195 _1384_ _1387_ _1386_ sg13g2_a21oi_1
X_6527_ net24 VGND VPWR _0037_ s0.was_valid_out\[20\][0] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_4788_ _2263_ net400 net1067 VPWR VGND sg13g2_nand2b_1
X_3739_ net1015 _2831_ _1322_ VPWR VGND sg13g2_nor2_1
X_6458_ net1242 VPWR _0979_ VGND _0918_ _0978_ sg13g2_o21ai_1
X_5409_ VPWR _2827_ net532 VGND sg13g2_inv_1
X_6389_ VPWR VGND _0913_ net1459 _0911_ net1456 _0914_ _0907_ sg13g2_a221oi_1
XFILLER_0_614 VPWR VGND sg13g2_decap_8
XFILLER_29_821 VPWR VGND sg13g2_fill_1
XFILLER_16_548 VPWR VGND sg13g2_fill_1
XFILLER_11_253 VPWR VGND sg13g2_fill_1
XFILLER_4_964 VPWR VGND sg13g2_decap_8
XFILLER_3_441 VPWR VGND sg13g2_decap_4
XFILLER_39_607 VPWR VGND sg13g2_decap_8
Xfanout1231 s0.shift_out\[15\][0] net1231 VPWR VGND sg13g2_buf_8
Xfanout1220 s0.valid_out\[14\][0] net1220 VPWR VGND sg13g2_buf_8
Xfanout1264 s0.shift_out\[18\][0] net1264 VPWR VGND sg13g2_buf_2
Xfanout1242 net1243 net1242 VPWR VGND sg13g2_buf_8
Xfanout1253 net1256 net1253 VPWR VGND sg13g2_buf_1
Xfanout1286 net1289 net1286 VPWR VGND sg13g2_buf_2
Xfanout1297 net1299 net1297 VPWR VGND sg13g2_buf_8
Xfanout1275 net1280 net1275 VPWR VGND sg13g2_buf_8
XFILLER_35_802 VPWR VGND sg13g2_decap_4
X_5760_ net1290 net1170 _0345_ VPWR VGND sg13g2_nor2b_1
X_4711_ VGND VPWR net1065 _2196_ _2198_ _2197_ sg13g2_a21oi_1
X_5691_ _3082_ _3084_ net1416 _3085_ VPWR VGND sg13g2_nand3_1
X_4642_ _2129_ VPWR _2132_ VGND net1077 _2131_ sg13g2_o21ai_1
X_4573_ net1403 _2062_ _2072_ VPWR VGND sg13g2_nor2_1
X_6312_ _0847_ _0845_ net1430 _0849_ VPWR VGND sg13g2_a21o_1
X_3524_ net1201 net1169 _1126_ VPWR VGND sg13g2_nor2b_1
X_6243_ net1477 net326 _0075_ VPWR VGND sg13g2_and2_1
X_3455_ _1069_ _1068_ net1230 VPWR VGND sg13g2_nand2b_1
X_6174_ s0.data_out\[18\]\[4\] s0.data_out\[17\]\[4\] net1259 _0723_ VPWR VGND sg13g2_mux2_1
X_5125_ net1041 VPWR _2569_ VGND _2513_ _2568_ sg13g2_o21ai_1
X_5056_ net1030 net1142 _2507_ VPWR VGND sg13g2_nor2b_1
X_4007_ net1491 VPWR _1564_ VGND _1561_ _1563_ sg13g2_o21ai_1
XFILLER_25_367 VPWR VGND sg13g2_decap_8
XFILLER_26_879 VPWR VGND sg13g2_fill_2
X_5958_ _0474_ _0529_ net1472 _0530_ VPWR VGND sg13g2_nand3_1
X_4909_ s0.data_out\[3\]\[1\] s0.data_out\[2\]\[1\] net1044 _2372_ VPWR VGND sg13g2_mux2_1
X_5889_ _0462_ net1284 net695 VPWR VGND sg13g2_nand2_1
XFILLER_4_205 VPWR VGND sg13g2_fill_2
XFILLER_20_21 VPWR VGND sg13g2_fill_1
XFILLER_1_912 VPWR VGND sg13g2_decap_8
XFILLER_0_400 VPWR VGND sg13g2_fill_1
XFILLER_0_422 VPWR VGND sg13g2_decap_4
XFILLER_49_905 VPWR VGND sg13g2_decap_8
Xhold41 s0.data_out\[0\]\[7\] VPWR VGND net361 sg13g2_dlygate4sd3_1
Xhold30 s0.was_valid_out\[10\][0] VPWR VGND net350 sg13g2_dlygate4sd3_1
XFILLER_0_488 VPWR VGND sg13g2_decap_8
XFILLER_1_989 VPWR VGND sg13g2_decap_8
Xhold52 _1731_ VPWR VGND net372 sg13g2_dlygate4sd3_1
Xhold74 s0.data_out\[0\]\[6\] VPWR VGND net394 sg13g2_dlygate4sd3_1
Xhold63 s0.was_valid_out\[17\][0] VPWR VGND net383 sg13g2_dlygate4sd3_1
Xhold85 _2061_ VPWR VGND net405 sg13g2_dlygate4sd3_1
Xhold96 s0.data_out\[23\]\[4\] VPWR VGND net416 sg13g2_dlygate4sd3_1
XFILLER_16_323 VPWR VGND sg13g2_decap_8
XFILLER_17_835 VPWR VGND sg13g2_fill_1
XFILLER_43_131 VPWR VGND sg13g2_fill_2
XFILLER_16_334 VPWR VGND sg13g2_fill_2
XFILLER_16_356 VPWR VGND sg13g2_fill_1
XFILLER_4_783 VPWR VGND sg13g2_decap_8
XFILLER_39_426 VPWR VGND sg13g2_fill_2
XFILLER_6_1005 VPWR VGND sg13g2_decap_8
Xfanout1083 net1084 net1083 VPWR VGND sg13g2_buf_1
Xfanout1072 net1073 net1072 VPWR VGND sg13g2_buf_8
Xfanout1061 net1063 net1061 VPWR VGND sg13g2_buf_8
Xfanout1050 net1055 net1050 VPWR VGND sg13g2_buf_8
Xfanout1094 net1095 net1094 VPWR VGND sg13g2_buf_8
XFILLER_23_805 VPWR VGND sg13g2_fill_2
X_5812_ _0394_ _0396_ net1427 _0397_ VPWR VGND sg13g2_nand3_1
XFILLER_34_153 VPWR VGND sg13g2_decap_4
X_5743_ _0331_ _0330_ net698 VPWR VGND sg13g2_nand2b_1
XFILLER_31_882 VPWR VGND sg13g2_fill_1
X_5674_ net1398 _3058_ _3068_ VPWR VGND sg13g2_nor2_1
X_4625_ _2117_ VPWR _2118_ VGND net1480 net630 sg13g2_o21ai_1
X_4556_ _2052_ _2054_ _2055_ VPWR VGND sg13g2_nor2_1
X_3507_ net1018 VPWR _1112_ VGND net566 net1222 sg13g2_o21ai_1
X_4487_ _0206_ _1993_ _1994_ _2858_ net1371 VPWR VGND sg13g2_a22oi_1
X_6226_ _0767_ net1470 _0768_ VPWR VGND _0716_ sg13g2_nand3b_1
X_3438_ VGND VPWR _1052_ _1042_ net1404 sg13g2_or2_1
X_6157_ net1249 net1143 _0706_ VPWR VGND sg13g2_nor2b_1
X_5108_ _2555_ VPWR _2556_ VGND net1468 net582 sg13g2_o21ai_1
XFILLER_39_982 VPWR VGND sg13g2_decap_8
X_6088_ _0055_ _0644_ _0645_ _2795_ net1355 VPWR VGND sg13g2_a22oi_1
X_5039_ _2490_ net1009 _2489_ VPWR VGND sg13g2_nand2_1
XFILLER_15_98 VPWR VGND sg13g2_fill_2
XFILLER_22_860 VPWR VGND sg13g2_fill_1
Xoutput7 net7 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_49_702 VPWR VGND sg13g2_decap_8
XFILLER_1_786 VPWR VGND sg13g2_decap_8
XFILLER_49_779 VPWR VGND sg13g2_decap_8
XFILLER_45_963 VPWR VGND sg13g2_decap_8
XFILLER_29_492 VPWR VGND sg13g2_decap_4
XFILLER_17_698 VPWR VGND sg13g2_decap_8
XFILLER_16_186 VPWR VGND sg13g2_fill_1
XFILLER_12_381 VPWR VGND sg13g2_decap_8
X_4410_ _1919_ net1085 _1920_ _1921_ VPWR VGND sg13g2_a21o_1
X_5390_ VPWR _2808_ net503 VGND sg13g2_inv_1
X_4341_ _1864_ net639 net1119 VPWR VGND sg13g2_nand2b_1
X_4272_ _1798_ _1795_ _1797_ VPWR VGND sg13g2_nand2_1
X_6011_ net1265 net1167 _0572_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_429 VPWR VGND sg13g2_decap_4
XFILLER_23_624 VPWR VGND sg13g2_fill_2
XFILLER_35_462 VPWR VGND sg13g2_fill_2
XFILLER_22_134 VPWR VGND sg13g2_decap_8
X_6775_ net203 VGND VPWR _0285_ s0.valid_out\[0\][0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3987_ _1509_ _1546_ net1490 _1547_ VPWR VGND sg13g2_nand3_1
X_5726_ VGND VPWR net1012 _3083_ _0317_ net1340 sg13g2_a21oi_1
X_5657_ _3048_ _3050_ _3051_ VPWR VGND sg13g2_nor2_1
X_5588_ net1317 s0.data_out\[22\]\[2\] _2991_ VPWR VGND sg13g2_and2_1
X_4608_ VGND VPWR net1074 net606 _2104_ _2045_ sg13g2_a21oi_1
Xhold330 s0.data_out\[21\]\[6\] VPWR VGND net650 sg13g2_dlygate4sd3_1
Xhold352 s0.data_out\[20\]\[0\] VPWR VGND net672 sg13g2_dlygate4sd3_1
Xhold341 s0.data_out\[11\]\[0\] VPWR VGND net661 sg13g2_dlygate4sd3_1
X_4539_ _2036_ net1075 _2037_ _2038_ VPWR VGND sg13g2_a21o_1
Xhold374 _1102_ VPWR VGND net694 sg13g2_dlygate4sd3_1
Xhold385 s0.data_new_delayed\[0\] VPWR VGND net705 sg13g2_dlygate4sd3_1
Xhold363 s0.data_out\[1\]\[2\] VPWR VGND net683 sg13g2_dlygate4sd3_1
X_6209_ net1268 VPWR _0755_ VGND _0674_ _0754_ sg13g2_o21ai_1
XFILLER_46_705 VPWR VGND sg13g2_fill_2
XFILLER_26_20 VPWR VGND sg13g2_decap_4
XFILLER_42_922 VPWR VGND sg13g2_decap_8
XFILLER_27_985 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_26_495 VPWR VGND sg13g2_decap_8
XFILLER_42_999 VPWR VGND sg13g2_decap_8
XFILLER_14_679 VPWR VGND sg13g2_fill_1
XFILLER_10_841 VPWR VGND sg13g2_fill_1
XFILLER_5_344 VPWR VGND sg13g2_fill_1
XFILLER_5_377 VPWR VGND sg13g2_decap_8
XFILLER_1_561 VPWR VGND sg13g2_decap_8
XFILLER_49_576 VPWR VGND sg13g2_decap_8
XFILLER_45_793 VPWR VGND sg13g2_decap_8
X_4890_ _2356_ _2355_ _2354_ VPWR VGND sg13g2_nand2b_1
X_3910_ _1461_ VPWR _1476_ VGND net1454 _1468_ sg13g2_o21ai_1
XFILLER_32_421 VPWR VGND sg13g2_decap_4
X_3841_ _1346_ _1418_ net1484 _1419_ VPWR VGND sg13g2_nand3_1
X_6560_ net284 VGND VPWR _0070_ s0.data_out\[18\]\[5\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3772_ VPWR VGND _1350_ net1459 _1346_ net1455 _1351_ _1344_ sg13g2_a221oi_1
X_6673__162 VPWR VGND net162 sg13g2_tiehi
X_5511_ net1315 net1166 _2917_ VPWR VGND sg13g2_nor2b_1
X_6491_ net63 VGND VPWR _0001_ s0.was_valid_out\[23\][0] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5442_ VPWR _2860_ net404 VGND sg13g2_inv_1
X_5373_ VPWR _2791_ net506 VGND sg13g2_inv_1
X_4324_ _1847_ _1846_ net1403 _1839_ net1412 VPWR VGND sg13g2_a22oi_1
X_4255_ _1783_ VPWR _1784_ VGND net1489 net680 sg13g2_o21ai_1
X_4186_ net1116 net1149 _1721_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_760 VPWR VGND sg13g2_decap_4
XFILLER_35_270 VPWR VGND sg13g2_fill_1
XFILLER_24_977 VPWR VGND sg13g2_decap_8
X_6758_ net70 VGND VPWR _0268_ s0.data_out\[2\]\[4\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_6537__309 VPWR VGND net309 sg13g2_tiehi
X_6517__34 VPWR VGND net34 sg13g2_tiehi
X_6689_ net145 VGND VPWR _0199_ s0.data_out\[8\]\[7\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_5709_ net1342 _3022_ _0304_ VPWR VGND sg13g2_nor2_1
XFILLER_12_88 VPWR VGND sg13g2_fill_2
XFILLER_3_859 VPWR VGND sg13g2_decap_8
Xhold171 s0.data_out\[13\]\[4\] VPWR VGND net491 sg13g2_dlygate4sd3_1
Xhold160 _0090_ VPWR VGND net480 sg13g2_dlygate4sd3_1
Xhold193 _0271_ VPWR VGND net513 sg13g2_dlygate4sd3_1
Xhold182 _0217_ VPWR VGND net502 sg13g2_dlygate4sd3_1
XFILLER_46_513 VPWR VGND sg13g2_fill_1
XFILLER_19_716 VPWR VGND sg13g2_fill_1
XFILLER_26_270 VPWR VGND sg13g2_decap_4
XFILLER_27_782 VPWR VGND sg13g2_fill_1
XFILLER_15_999 VPWR VGND sg13g2_decap_8
XFILLER_30_947 VPWR VGND sg13g2_decap_8
X_6657__179 VPWR VGND net179 sg13g2_tiehi
XFILLER_6_686 VPWR VGND sg13g2_decap_4
XFILLER_5_174 VPWR VGND sg13g2_fill_2
X_4040_ s0.data_out\[9\]\[2\] s0.data_out\[10\]\[2\] net1174 _1587_ VPWR VGND sg13g2_mux2_1
XFILLER_49_395 VPWR VGND sg13g2_decap_8
X_5991_ _0553_ _0554_ _0555_ VPWR VGND sg13g2_nor2_1
XFILLER_24_218 VPWR VGND sg13g2_decap_8
X_4942_ _2403_ net1041 _2404_ _2405_ VPWR VGND sg13g2_a21o_1
XFILLER_24_229 VPWR VGND sg13g2_fill_1
XFILLER_17_292 VPWR VGND sg13g2_fill_1
XFILLER_21_903 VPWR VGND sg13g2_fill_1
XFILLER_21_914 VPWR VGND sg13g2_fill_2
XFILLER_33_752 VPWR VGND sg13g2_fill_1
X_6612_ net227 VGND VPWR _0122_ s0.valid_out\[13\][0] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_20_424 VPWR VGND sg13g2_fill_1
X_4873_ _2342_ VPWR _2343_ VGND net1473 net569 sg13g2_o21ai_1
X_3824_ _1403_ net1195 _1402_ VPWR VGND sg13g2_nand2b_1
X_6543_ net302 VGND VPWR _0053_ s0.data_out\[19\]\[0\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_3755_ _1336_ _1333_ _1335_ VPWR VGND sg13g2_nand2_1
X_6474_ net1224 s0.data_out\[15\]\[7\] _0991_ VPWR VGND sg13g2_and2_1
X_3686_ s0.data_out\[13\]\[5\] s0.data_out\[12\]\[5\] net1198 _1276_ VPWR VGND sg13g2_mux2_1
X_5425_ VPWR _2843_ net572 VGND sg13g2_inv_1
X_5356_ _2774_ net1443 VPWR VGND sg13g2_inv_2
X_5287_ VGND VPWR _2714_ _2712_ net1408 sg13g2_or2_1
X_4307_ VGND VPWR net1112 _1827_ _1830_ _1829_ sg13g2_a21oi_1
X_4238_ _0181_ _1769_ _1770_ _2843_ net1374 VPWR VGND sg13g2_a22oi_1
X_6543__302 VPWR VGND net302 sg13g2_tiehi
XFILLER_28_535 VPWR VGND sg13g2_fill_1
X_4169_ VGND VPWR net1111 _1702_ _1704_ _1703_ sg13g2_a21oi_1
XFILLER_24_785 VPWR VGND sg13g2_fill_1
Xfanout1402 net1406 net1402 VPWR VGND sg13g2_buf_8
Xfanout1413 net1415 net1413 VPWR VGND sg13g2_buf_8
Xfanout1424 net1425 net1424 VPWR VGND sg13g2_buf_8
Xfanout1446 net1448 net1446 VPWR VGND sg13g2_buf_8
Xfanout1457 ui_in[1] net1457 VPWR VGND sg13g2_buf_8
Xfanout1435 net1438 net1435 VPWR VGND sg13g2_buf_8
XFILLER_47_822 VPWR VGND sg13g2_decap_8
Xfanout1479 net1482 net1479 VPWR VGND sg13g2_buf_8
Xfanout1468 net1469 net1468 VPWR VGND sg13g2_buf_8
XFILLER_46_332 VPWR VGND sg13g2_fill_2
XFILLER_0_25 VPWR VGND sg13g2_decap_8
XFILLER_47_899 VPWR VGND sg13g2_decap_8
XFILLER_0_36 VPWR VGND sg13g2_decap_8
XFILLER_15_730 VPWR VGND sg13g2_fill_1
XFILLER_31_1013 VPWR VGND sg13g2_decap_8
X_3540_ _1140_ net1203 _1141_ _1142_ VPWR VGND sg13g2_a21o_1
XFILLER_7_995 VPWR VGND sg13g2_decap_8
X_6670__165 VPWR VGND net165 sg13g2_tiehi
X_5210_ _2628_ _2636_ _2645_ _2648_ _2649_ VPWR VGND sg13g2_nor4_1
X_3471_ net1018 _2824_ _1083_ VPWR VGND sg13g2_nor2_1
XFILLER_9_1003 VPWR VGND sg13g2_decap_8
X_6190_ net1439 _0702_ _0739_ VPWR VGND sg13g2_nor2_1
X_5141_ _2581_ _2582_ _0272_ VPWR VGND sg13g2_nor2_1
X_5072_ s0.data_out\[2\]\[4\] s0.data_out\[1\]\[4\] net1035 _2523_ VPWR VGND sg13g2_mux2_1
X_4023_ net1124 net1168 _1570_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_192 VPWR VGND sg13g2_fill_2
XFILLER_49_170 VPWR VGND sg13g2_fill_2
XFILLER_25_516 VPWR VGND sg13g2_fill_2
XFILLER_25_549 VPWR VGND sg13g2_fill_1
X_5974_ net1295 VPWR _0542_ VGND _0507_ _0541_ sg13g2_o21ai_1
XFILLER_21_700 VPWR VGND sg13g2_decap_8
X_4925_ _2387_ VPWR _2388_ VGND net1044 _2877_ sg13g2_o21ai_1
X_4856_ _2329_ VPWR _2330_ VGND net1473 net600 sg13g2_o21ai_1
X_3807_ VGND VPWR _1265_ _1385_ _1386_ net1194 sg13g2_a21oi_1
X_6526_ net25 VGND VPWR _0036_ s0.data_out\[21\]\[7\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_4787_ _2260_ net1049 _2261_ _2262_ VPWR VGND sg13g2_a21o_1
X_3738_ VPWR _0130_ _1321_ VGND sg13g2_inv_1
X_6457_ net1225 s0.data_out\[15\]\[3\] _0978_ VPWR VGND sg13g2_and2_1
X_3669_ s0.data_out\[13\]\[7\] s0.data_out\[12\]\[7\] net1198 _1259_ VPWR VGND sg13g2_mux2_1
X_5408_ VPWR _2826_ net491 VGND sg13g2_inv_1
X_6388_ _0913_ _0912_ net1243 VPWR VGND sg13g2_nand2b_1
X_5339_ _2757_ net1254 VPWR VGND sg13g2_inv_2
XFILLER_47_129 VPWR VGND sg13g2_fill_1
XFILLER_43_324 VPWR VGND sg13g2_fill_1
XFILLER_28_387 VPWR VGND sg13g2_decap_4
XFILLER_12_700 VPWR VGND sg13g2_decap_8
XFILLER_11_298 VPWR VGND sg13g2_fill_2
XFILLER_4_943 VPWR VGND sg13g2_decap_8
Xfanout1232 net1233 net1232 VPWR VGND sg13g2_buf_8
Xfanout1221 s0.valid_out\[14\][0] net1221 VPWR VGND sg13g2_buf_8
Xfanout1210 net1212 net1210 VPWR VGND sg13g2_buf_8
Xfanout1254 net1256 net1254 VPWR VGND sg13g2_buf_8
Xfanout1265 net1266 net1265 VPWR VGND sg13g2_buf_8
Xfanout1243 net1244 net1243 VPWR VGND sg13g2_buf_1
Xfanout1287 net1289 net1287 VPWR VGND sg13g2_buf_8
Xfanout1298 net1299 net1298 VPWR VGND sg13g2_buf_1
Xfanout1276 net1277 net1276 VPWR VGND sg13g2_buf_8
XFILLER_47_685 VPWR VGND sg13g2_decap_8
XFILLER_34_324 VPWR VGND sg13g2_fill_2
XFILLER_15_571 VPWR VGND sg13g2_fill_1
XFILLER_42_390 VPWR VGND sg13g2_decap_8
X_4710_ net1065 net1151 _2197_ VPWR VGND sg13g2_nor2b_1
X_5690_ _3084_ net1012 _3083_ VPWR VGND sg13g2_nand2_1
X_4641_ s0.was_valid_out\[4\][0] net1082 _2131_ VPWR VGND sg13g2_nor2_1
X_4572_ VGND VPWR _2071_ _2069_ net1412 sg13g2_or2_1
X_6311_ _0845_ _0847_ net1430 _0848_ VPWR VGND sg13g2_nand3_1
X_3523_ _1124_ VPWR _1125_ VGND net1210 _2824_ sg13g2_o21ai_1
X_6242_ net1478 _0775_ _0074_ VPWR VGND sg13g2_and2_1
X_3454_ _0945_ VPWR _1068_ VGND net1234 _2821_ sg13g2_o21ai_1
XFILLER_41_0 VPWR VGND sg13g2_decap_4
X_6173_ _0722_ net1257 s0.data_out\[17\]\[4\] VPWR VGND sg13g2_nand2_1
X_5124_ net1032 s0.data_out\[1\]\[6\] _2568_ VPWR VGND sg13g2_and2_1
X_5055_ s0.data_out\[2\]\[7\] s0.data_out\[1\]\[7\] net1034 _2506_ VPWR VGND sg13g2_mux2_1
X_4006_ _1563_ _1560_ _1562_ VPWR VGND sg13g2_nand2_1
X_6540__305 VPWR VGND net305 sg13g2_tiehi
XFILLER_26_847 VPWR VGND sg13g2_fill_1
XFILLER_38_1019 VPWR VGND sg13g2_decap_8
XFILLER_26_869 VPWR VGND sg13g2_fill_1
X_5957_ net1293 VPWR _0529_ VGND _0470_ _0528_ sg13g2_o21ai_1
X_6718__113 VPWR VGND net113 sg13g2_tiehi
X_4908_ _2371_ net1043 net514 VPWR VGND sg13g2_nand2_1
XFILLER_33_390 VPWR VGND sg13g2_fill_1
XFILLER_34_891 VPWR VGND sg13g2_fill_2
X_5888_ VGND VPWR _0461_ _0460_ net1444 sg13g2_or2_1
XFILLER_21_541 VPWR VGND sg13g2_decap_4
X_4839_ VGND VPWR net1053 _2312_ _2314_ _2313_ sg13g2_a21oi_1
XFILLER_5_707 VPWR VGND sg13g2_decap_8
X_6509_ net43 VGND VPWR _0019_ s0.data_out\[22\]\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_2
XFILLER_0_412 VPWR VGND sg13g2_decap_4
XFILLER_1_968 VPWR VGND sg13g2_decap_8
X_6725__106 VPWR VGND net106 sg13g2_tiehi
Xhold20 s0.genblk1\[3\].modules.bubble VPWR VGND net340 sg13g2_dlygate4sd3_1
Xhold31 _0157_ VPWR VGND net351 sg13g2_dlygate4sd3_1
XFILLER_0_456 VPWR VGND sg13g2_decap_4
XFILLER_0_467 VPWR VGND sg13g2_decap_8
Xhold64 s0.shift_out\[5\][0] VPWR VGND net384 sg13g2_dlygate4sd3_1
Xhold42 s0.was_valid_out\[15\][0] VPWR VGND net362 sg13g2_dlygate4sd3_1
XFILLER_29_64 VPWR VGND sg13g2_fill_2
Xhold53 s0.data_out\[11\]\[4\] VPWR VGND net373 sg13g2_dlygate4sd3_1
Xhold75 s0.data_out\[0\]\[5\] VPWR VGND net395 sg13g2_dlygate4sd3_1
Xhold97 _0009_ VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold86 s0.data_out\[13\]\[7\] VPWR VGND net406 sg13g2_dlygate4sd3_1
XFILLER_17_825 VPWR VGND sg13g2_decap_4
XFILLER_8_512 VPWR VGND sg13g2_decap_8
XFILLER_12_563 VPWR VGND sg13g2_fill_2
Xfanout1040 net1041 net1040 VPWR VGND sg13g2_buf_8
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
Xfanout1051 net1054 net1051 VPWR VGND sg13g2_buf_8
Xfanout1073 net384 net1073 VPWR VGND sg13g2_buf_8
Xfanout1062 net1063 net1062 VPWR VGND sg13g2_buf_1
Xfanout1084 net711 net1084 VPWR VGND sg13g2_buf_8
Xfanout1095 s0.valid_out\[6\][0] net1095 VPWR VGND sg13g2_buf_8
X_5811_ _0396_ net1007 _0395_ VPWR VGND sg13g2_nand2_1
X_5742_ _0328_ _0329_ _0330_ VPWR VGND sg13g2_nor2_1
XFILLER_31_850 VPWR VGND sg13g2_fill_2
X_5673_ VGND VPWR _3067_ _3065_ net1407 sg13g2_or2_1
X_4624_ _2116_ VPWR _2117_ VGND net999 _2115_ sg13g2_o21ai_1
X_4555_ _2053_ VPWR _2054_ VGND _2042_ _2050_ sg13g2_o21ai_1
X_3506_ VGND VPWR _1111_ net1211 net566 sg13g2_or2_1
X_4486_ net1371 _1915_ _1994_ VPWR VGND sg13g2_nor2_1
X_6225_ net1262 VPWR _0767_ VGND _0713_ _0766_ sg13g2_o21ai_1
X_3437_ VGND VPWR _1051_ _1049_ net1413 sg13g2_or2_1
XFILLER_44_1023 VPWR VGND sg13g2_decap_4
X_6156_ s0.data_out\[18\]\[7\] s0.data_out\[17\]\[7\] net1258 _0705_ VPWR VGND sg13g2_mux2_1
X_5107_ _2490_ _2554_ net1468 _2555_ VPWR VGND sg13g2_nand3_1
XFILLER_39_961 VPWR VGND sg13g2_decap_8
X_6087_ net1355 _0567_ _0645_ VPWR VGND sg13g2_nor2_1
X_5038_ s0.data_out\[1\]\[2\] s0.data_out\[2\]\[2\] net1043 _2489_ VPWR VGND sg13g2_mux2_1
XFILLER_41_647 VPWR VGND sg13g2_fill_1
XFILLER_40_113 VPWR VGND sg13g2_fill_1
XFILLER_15_66 VPWR VGND sg13g2_fill_1
Xoutput8 net8 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_253 VPWR VGND sg13g2_fill_2
XFILLER_0_242 VPWR VGND sg13g2_decap_8
XFILLER_1_765 VPWR VGND sg13g2_decap_8
XFILLER_49_758 VPWR VGND sg13g2_decap_8
XFILLER_0_297 VPWR VGND sg13g2_fill_1
XFILLER_48_257 VPWR VGND sg13g2_fill_2
XFILLER_45_942 VPWR VGND sg13g2_decap_8
XFILLER_44_441 VPWR VGND sg13g2_decap_4
XFILLER_13_872 VPWR VGND sg13g2_decap_8
XFILLER_31_157 VPWR VGND sg13g2_decap_8
XFILLER_31_168 VPWR VGND sg13g2_fill_1
XFILLER_9_865 VPWR VGND sg13g2_fill_2
X_4340_ _1861_ net1102 _1862_ _1863_ VPWR VGND sg13g2_a21o_1
X_4271_ _2759_ VPWR _1797_ VGND s0.was_valid_out\[7\][0] net1120 sg13g2_o21ai_1
XFILLER_28_1018 VPWR VGND sg13g2_decap_8
X_6010_ _0570_ VPWR _0571_ VGND net1270 _2796_ sg13g2_o21ai_1
XFILLER_39_257 VPWR VGND sg13g2_decap_4
XFILLER_39_279 VPWR VGND sg13g2_fill_1
XFILLER_36_986 VPWR VGND sg13g2_decap_8
X_6774_ net228 VGND VPWR _0284_ s0.was_valid_out\[0\][0] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_3986_ net1184 VPWR _1546_ VGND _1505_ _1545_ sg13g2_o21ai_1
X_5725_ VGND VPWR net1300 s0.data_out\[21\]\[5\] _0316_ _3080_ sg13g2_a21oi_1
X_6715__116 VPWR VGND net116 sg13g2_tiehi
X_5656_ _3049_ VPWR _3050_ VGND _3039_ _3046_ sg13g2_o21ai_1
XFILLER_30_190 VPWR VGND sg13g2_decap_8
XFILLER_11_1011 VPWR VGND sg13g2_decap_8
X_4607_ _0217_ _2102_ _2103_ _2863_ net1370 VPWR VGND sg13g2_a22oi_1
X_5587_ _0006_ _2989_ _2990_ _2776_ net1341 VPWR VGND sg13g2_a22oi_1
Xhold320 s0.data_out\[22\]\[1\] VPWR VGND net640 sg13g2_dlygate4sd3_1
Xhold342 s0.data_out\[16\]\[0\] VPWR VGND net662 sg13g2_dlygate4sd3_1
Xhold353 s0.data_out\[8\]\[1\] VPWR VGND net673 sg13g2_dlygate4sd3_1
Xhold331 s0.data_out\[12\]\[2\] VPWR VGND net651 sg13g2_dlygate4sd3_1
X_4538_ net1075 net1161 _2037_ VPWR VGND sg13g2_nor2b_1
Xhold386 s0.valid_out\[4\][0] VPWR VGND net706 sg13g2_dlygate4sd3_1
X_4469_ _1966_ VPWR _1980_ VGND _1973_ _1975_ sg13g2_o21ai_1
Xhold364 s0.data_out\[14\]\[5\] VPWR VGND net684 sg13g2_dlygate4sd3_1
XFILLER_7_9 VPWR VGND sg13g2_decap_8
Xhold375 s0.data_out\[19\]\[1\] VPWR VGND net695 sg13g2_dlygate4sd3_1
X_6208_ _2757_ _2806_ _0754_ VPWR VGND sg13g2_nor2_1
XFILLER_46_717 VPWR VGND sg13g2_decap_4
X_6139_ net1252 net1172 _0688_ VPWR VGND sg13g2_nor2b_1
X_6722__109 VPWR VGND net109 sg13g2_tiehi
XFILLER_18_419 VPWR VGND sg13g2_decap_8
XFILLER_27_964 VPWR VGND sg13g2_decap_8
XFILLER_26_485 VPWR VGND sg13g2_fill_1
XFILLER_42_978 VPWR VGND sg13g2_decap_8
XFILLER_13_146 VPWR VGND sg13g2_decap_8
XFILLER_14_658 VPWR VGND sg13g2_fill_2
XFILLER_13_179 VPWR VGND sg13g2_fill_1
X_6772__254 VPWR VGND net254 sg13g2_tiehi
XFILLER_5_301 VPWR VGND sg13g2_fill_1
XFILLER_10_864 VPWR VGND sg13g2_fill_1
XFILLER_6_879 VPWR VGND sg13g2_decap_8
XFILLER_1_540 VPWR VGND sg13g2_decap_8
XFILLER_49_555 VPWR VGND sg13g2_decap_8
X_6666__170 VPWR VGND net170 sg13g2_tiehi
XFILLER_36_238 VPWR VGND sg13g2_decap_8
XFILLER_36_227 VPWR VGND sg13g2_fill_2
XFILLER_45_772 VPWR VGND sg13g2_decap_8
XFILLER_32_400 VPWR VGND sg13g2_decap_8
X_3840_ net1191 VPWR _1418_ VGND _1347_ _1417_ sg13g2_o21ai_1
XFILLER_13_680 VPWR VGND sg13g2_decap_8
X_3771_ _1350_ net1191 _1349_ VPWR VGND sg13g2_nand2b_1
XFILLER_32_477 VPWR VGND sg13g2_decap_4
X_5510_ _2915_ VPWR _2916_ VGND net1320 _2776_ sg13g2_o21ai_1
X_6490_ net215 VGND VPWR _0000_ s0.module0.bubble clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5441_ VPWR _2859_ net408 VGND sg13g2_inv_1
X_5372_ VPWR _2790_ net633 VGND sg13g2_inv_1
X_4323_ VGND VPWR net1115 _1843_ _1846_ _1845_ sg13g2_a21oi_1
X_4254_ _1743_ _1782_ net1489 _1783_ VPWR VGND sg13g2_nand3_1
X_4185_ s0.data_out\[9\]\[6\] s0.data_out\[8\]\[6\] net1121 _1720_ VPWR VGND sg13g2_mux2_1
XFILLER_41_1015 VPWR VGND sg13g2_decap_8
XFILLER_28_717 VPWR VGND sg13g2_decap_8
XFILLER_42_219 VPWR VGND sg13g2_fill_1
X_6757_ net71 VGND VPWR net464 s0.data_out\[2\]\[3\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_5708_ net1316 VPWR _0303_ VGND _3019_ _0302_ sg13g2_o21ai_1
X_3969_ net1014 _2839_ _1533_ VPWR VGND sg13g2_nor2_1
X_6688_ net146 VGND VPWR _0198_ s0.data_out\[8\]\[6\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_12_23 VPWR VGND sg13g2_fill_2
X_5639_ s0.data_out\[22\]\[3\] s0.data_out\[21\]\[3\] net1307 _3033_ VPWR VGND sg13g2_mux2_1
XFILLER_3_838 VPWR VGND sg13g2_decap_8
Xhold150 s0.data_out\[7\]\[5\] VPWR VGND net470 sg13g2_dlygate4sd3_1
Xhold161 s0.data_out\[13\]\[1\] VPWR VGND net481 sg13g2_dlygate4sd3_1
Xhold172 s0.data_out\[4\]\[7\] VPWR VGND net492 sg13g2_dlygate4sd3_1
Xhold183 s0.data_out\[16\]\[7\] VPWR VGND net503 sg13g2_dlygate4sd3_1
Xhold194 s0.data_out\[2\]\[1\] VPWR VGND net514 sg13g2_dlygate4sd3_1
XFILLER_37_42 VPWR VGND sg13g2_fill_1
XFILLER_37_53 VPWR VGND sg13g2_decap_8
XFILLER_42_720 VPWR VGND sg13g2_fill_1
XFILLER_15_923 VPWR VGND sg13g2_fill_1
XFILLER_15_978 VPWR VGND sg13g2_decap_8
XFILLER_6_676 VPWR VGND sg13g2_decap_4
XFILLER_2_882 VPWR VGND sg13g2_decap_8
X_5990_ net1394 _2756_ _0554_ VPWR VGND sg13g2_nor2_1
X_4941_ net1040 net1147 _2404_ VPWR VGND sg13g2_nor2b_1
X_4872_ _2341_ VPWR _2342_ VGND net995 _2340_ sg13g2_o21ai_1
X_6611_ net229 VGND VPWR net567 s0.was_valid_out\[13\][0] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_3823_ VGND VPWR net1182 _1400_ _1402_ _1401_ sg13g2_a21oi_1
X_6536__310 VPWR VGND net310 sg13g2_tiehi
X_6542_ net303 VGND VPWR _0052_ s0.shift_out\[19\][0] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3754_ net1015 VPWR _1335_ VGND s0.was_valid_out\[11\][0] net1198 sg13g2_o21ai_1
X_6473_ VPWR _0095_ _0990_ VGND sg13g2_inv_1
XFILLER_9_492 VPWR VGND sg13g2_decap_4
X_3685_ _1275_ _1272_ _1273_ _1274_ VPWR VGND sg13g2_and3_1
X_5424_ VPWR _2842_ net636 VGND sg13g2_inv_1
X_6514__38 VPWR VGND net38 sg13g2_tiehi
X_5355_ VPWR _2773_ net412 VGND sg13g2_inv_1
X_5286_ _2713_ _2712_ net1408 _2688_ net1416 VPWR VGND sg13g2_a22oi_1
X_4306_ VGND VPWR _1710_ _1828_ _1829_ net1112 sg13g2_a21oi_1
X_4237_ net1374 _1700_ _1770_ VPWR VGND sg13g2_nor2_1
X_4168_ net1111 net1171 _1703_ VPWR VGND sg13g2_nor2b_1
X_4099_ _1559_ VPWR _1646_ VGND _1619_ _1621_ sg13g2_o21ai_1
XFILLER_24_720 VPWR VGND sg13g2_decap_4
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_8_919 VPWR VGND sg13g2_decap_8
XFILLER_11_436 VPWR VGND sg13g2_fill_1
XFILLER_7_429 VPWR VGND sg13g2_fill_2
XFILLER_11_469 VPWR VGND sg13g2_fill_2
X_6656__180 VPWR VGND net180 sg13g2_tiehi
Xfanout1403 net1406 net1403 VPWR VGND sg13g2_buf_1
Xfanout1414 net1415 net1414 VPWR VGND sg13g2_buf_8
Xfanout1425 ui_in[5] net1425 VPWR VGND sg13g2_buf_8
Xfanout1447 net1448 net1447 VPWR VGND sg13g2_buf_8
Xfanout1436 net1438 net1436 VPWR VGND sg13g2_buf_1
XFILLER_47_801 VPWR VGND sg13g2_decap_8
Xfanout1469 net1476 net1469 VPWR VGND sg13g2_buf_8
Xfanout1458 net1461 net1458 VPWR VGND sg13g2_buf_8
X_6663__173 VPWR VGND net173 sg13g2_tiehi
XFILLER_19_525 VPWR VGND sg13g2_fill_1
XFILLER_47_878 VPWR VGND sg13g2_decap_8
XFILLER_10_480 VPWR VGND sg13g2_decap_8
XFILLER_7_974 VPWR VGND sg13g2_decap_8
XFILLER_6_462 VPWR VGND sg13g2_decap_4
XFILLER_10_491 VPWR VGND sg13g2_fill_1
X_3470_ VPWR _0101_ _1082_ VGND sg13g2_inv_1
X_5140_ net1468 VPWR _2582_ VGND net516 _2577_ sg13g2_o21ai_1
X_6781__117 VPWR VGND net117 sg13g2_tiehi
X_5071_ net1028 net1156 _2522_ VPWR VGND sg13g2_nor2b_1
X_4022_ s0.data_out\[10\]\[1\] s0.data_out\[9\]\[1\] net1133 _1569_ VPWR VGND sg13g2_mux2_1
X_5973_ _2755_ _2793_ _0541_ VPWR VGND sg13g2_nor2_1
XFILLER_25_539 VPWR VGND sg13g2_fill_1
X_4924_ _2387_ net1044 net463 VPWR VGND sg13g2_nand2_1
X_4855_ _2328_ VPWR _2329_ VGND net995 _2327_ sg13g2_o21ai_1
XFILLER_21_767 VPWR VGND sg13g2_fill_2
X_3806_ _1385_ s0.data_out\[11\]\[6\] net1199 VPWR VGND sg13g2_nand2b_1
X_4786_ net1049 net1167 _2261_ VPWR VGND sg13g2_nor2b_1
X_6525_ net26 VGND VPWR _0035_ s0.data_out\[21\]\[6\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_3737_ _1320_ VPWR _1321_ VGND net1486 net686 sg13g2_o21ai_1
X_6456_ _0091_ _0976_ _0977_ _2812_ net1367 VPWR VGND sg13g2_a22oi_1
X_3668_ _1258_ net1199 net595 VPWR VGND sg13g2_nand2_1
X_3599_ net1216 VPWR _1198_ VGND _1118_ _1197_ sg13g2_o21ai_1
X_5407_ VPWR _2825_ net406 VGND sg13g2_inv_1
X_6387_ s0.data_out\[15\]\[0\] s0.data_out\[16\]\[0\] net1248 _0912_ VPWR VGND sg13g2_mux2_1
X_5338_ VPWR _2756_ net1272 VGND sg13g2_inv_1
XFILLER_0_649 VPWR VGND sg13g2_decap_8
X_5269_ _2695_ VPWR _2696_ VGND net1001 net1162 sg13g2_o21ai_1
XFILLER_28_355 VPWR VGND sg13g2_fill_1
XFILLER_18_88 VPWR VGND sg13g2_fill_1
XFILLER_43_358 VPWR VGND sg13g2_decap_4
XFILLER_12_723 VPWR VGND sg13g2_fill_1
XFILLER_12_745 VPWR VGND sg13g2_fill_1
XFILLER_12_778 VPWR VGND sg13g2_fill_1
XFILLER_4_922 VPWR VGND sg13g2_decap_8
XFILLER_4_999 VPWR VGND sg13g2_decap_8
X_6501__52 VPWR VGND net52 sg13g2_tiehi
Xfanout1222 s0.valid_out\[14\][0] net1222 VPWR VGND sg13g2_buf_1
Xfanout1211 net1212 net1211 VPWR VGND sg13g2_buf_8
Xfanout1200 s0.valid_out\[12\][0] net1200 VPWR VGND sg13g2_buf_8
Xfanout1233 net1235 net1233 VPWR VGND sg13g2_buf_8
Xfanout1244 net703 net1244 VPWR VGND sg13g2_buf_8
Xfanout1255 net1256 net1255 VPWR VGND sg13g2_buf_1
Xfanout1288 net1289 net1288 VPWR VGND sg13g2_buf_1
Xfanout1299 s0.valid_out\[20\][0] net1299 VPWR VGND sg13g2_buf_2
Xfanout1266 net472 net1266 VPWR VGND sg13g2_buf_8
Xfanout1277 net1280 net1277 VPWR VGND sg13g2_buf_2
XFILLER_47_664 VPWR VGND sg13g2_decap_8
XFILLER_47_642 VPWR VGND sg13g2_decap_8
XFILLER_15_583 VPWR VGND sg13g2_fill_2
X_4640_ net1065 _2125_ _2130_ VPWR VGND sg13g2_nor2_1
XFILLER_30_564 VPWR VGND sg13g2_decap_8
X_4571_ _2070_ _2069_ net1412 _2062_ net1403 VPWR VGND sg13g2_a22oi_1
X_6310_ _0847_ net1002 _0846_ VPWR VGND sg13g2_nand2_1
X_6533__313 VPWR VGND net313 sg13g2_tiehi
X_3522_ _1124_ net1210 net481 VPWR VGND sg13g2_nand2_1
X_6241_ VGND VPWR _2737_ _0775_ _0073_ _0780_ sg13g2_a21oi_1
X_3453_ _1067_ net1230 _1066_ VPWR VGND sg13g2_nand2b_1
X_6172_ _0720_ _0718_ _0721_ VPWR VGND _0719_ sg13g2_nand3b_1
X_5123_ VPWR _0269_ net577 VGND sg13g2_inv_1
XFILLER_34_0 VPWR VGND sg13g2_decap_8
X_5054_ _2502_ _2504_ _2505_ VPWR VGND sg13g2_nor2_1
X_4005_ net1014 VPWR _1562_ VGND s0.was_valid_out\[9\][0] net1174 sg13g2_o21ai_1
X_5956_ net1276 s0.data_out\[19\]\[0\] _0528_ VPWR VGND sg13g2_and2_1
XFILLER_34_870 VPWR VGND sg13g2_decap_8
X_5887_ VGND VPWR net1293 _0457_ _0460_ _0459_ sg13g2_a21oi_1
XFILLER_21_520 VPWR VGND sg13g2_fill_2
X_4907_ net1444 _2369_ _2370_ VPWR VGND sg13g2_nor2_1
X_4838_ net1053 net1152 _2313_ VPWR VGND sg13g2_nor2b_1
XFILLER_14_1020 VPWR VGND sg13g2_decap_8
X_4769_ _2243_ VPWR _2247_ VGND net524 net1059 sg13g2_o21ai_1
X_6508_ net44 VGND VPWR net641 s0.data_out\[22\]\[1\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_6653__183 VPWR VGND net183 sg13g2_tiehi
X_6439_ _0944_ _0960_ _0962_ _0963_ _0964_ VPWR VGND sg13g2_nor4_1
XFILLER_20_89 VPWR VGND sg13g2_fill_2
XFILLER_1_947 VPWR VGND sg13g2_decap_8
Xhold32 s0.data_out\[19\]\[5\] VPWR VGND net352 sg13g2_dlygate4sd3_1
Xhold10 s0.genblk1\[22\].modules.bubble VPWR VGND net330 sg13g2_dlygate4sd3_1
Xhold21 s0.genblk1\[11\].modules.bubble VPWR VGND net341 sg13g2_dlygate4sd3_1
Xhold43 _0097_ VPWR VGND net363 sg13g2_dlygate4sd3_1
Xhold54 _1515_ VPWR VGND net374 sg13g2_dlygate4sd3_1
Xhold65 s0.data_out\[0\]\[4\] VPWR VGND net385 sg13g2_dlygate4sd3_1
Xhold76 s0.valid_out\[2\][0] VPWR VGND net396 sg13g2_dlygate4sd3_1
Xhold87 _0132_ VPWR VGND net407 sg13g2_dlygate4sd3_1
Xhold98 s0.data_out\[18\]\[1\] VPWR VGND net418 sg13g2_dlygate4sd3_1
XFILLER_21_1013 VPWR VGND sg13g2_decap_8
XFILLER_43_100 VPWR VGND sg13g2_decap_4
XFILLER_43_122 VPWR VGND sg13g2_fill_1
X_6660__176 VPWR VGND net176 sg13g2_tiehi
XFILLER_28_196 VPWR VGND sg13g2_fill_2
XFILLER_43_144 VPWR VGND sg13g2_fill_2
XFILLER_31_339 VPWR VGND sg13g2_decap_8
XFILLER_40_851 VPWR VGND sg13g2_decap_8
XFILLER_4_796 VPWR VGND sg13g2_decap_8
Xfanout1030 net1032 net1030 VPWR VGND sg13g2_buf_8
XFILLER_39_417 VPWR VGND sg13g2_decap_4
XFILLER_39_406 VPWR VGND sg13g2_decap_8
Xfanout1052 net1054 net1052 VPWR VGND sg13g2_buf_1
Xfanout1041 net1042 net1041 VPWR VGND sg13g2_buf_8
Xfanout1063 net608 net1063 VPWR VGND sg13g2_buf_8
Xfanout1074 net1075 net1074 VPWR VGND sg13g2_buf_2
Xfanout1085 net1087 net1085 VPWR VGND sg13g2_buf_8
Xfanout1096 net1097 net1096 VPWR VGND sg13g2_buf_8
XFILLER_48_984 VPWR VGND sg13g2_decap_8
XFILLER_34_100 VPWR VGND sg13g2_fill_2
XFILLER_47_494 VPWR VGND sg13g2_fill_1
XFILLER_34_122 VPWR VGND sg13g2_decap_4
X_5810_ _3071_ VPWR _0395_ VGND net1309 _2787_ sg13g2_o21ai_1
XFILLER_16_870 VPWR VGND sg13g2_fill_1
XFILLER_23_818 VPWR VGND sg13g2_fill_2
X_5741_ VGND VPWR net1336 net1308 _0329_ net1301 sg13g2_a21oi_1
X_5672_ _3066_ _3065_ net1407 _3058_ net1398 VPWR VGND sg13g2_a22oi_1
XFILLER_30_372 VPWR VGND sg13g2_fill_1
X_4623_ VGND VPWR net999 _2085_ _2116_ net1372 sg13g2_a21oi_1
X_4554_ _2053_ net1439 _2041_ VPWR VGND sg13g2_nand2_1
X_3505_ _1109_ VPWR _1110_ VGND net1217 _0995_ sg13g2_o21ai_1
X_6224_ net1249 s0.data_out\[17\]\[6\] _0766_ VPWR VGND sg13g2_and2_1
X_4485_ net1096 VPWR _1993_ VGND _1912_ _1992_ sg13g2_o21ai_1
XFILLER_44_1002 VPWR VGND sg13g2_decap_8
X_3436_ _1050_ _1049_ net1413 _1042_ net1404 VPWR VGND sg13g2_a22oi_1
X_6155_ _0704_ net1257 net560 VPWR VGND sg13g2_nand2_1
X_6086_ net1278 VPWR _0644_ VGND _0564_ _0643_ sg13g2_o21ai_1
X_5106_ net1038 VPWR _2554_ VGND _2487_ _2553_ sg13g2_o21ai_1
XFILLER_39_940 VPWR VGND sg13g2_decap_8
X_5037_ VGND VPWR net1027 _2486_ _2488_ _2487_ sg13g2_a21oi_1
XFILLER_26_623 VPWR VGND sg13g2_decap_4
XFILLER_26_656 VPWR VGND sg13g2_fill_2
XFILLER_41_637 VPWR VGND sg13g2_fill_2
XFILLER_25_199 VPWR VGND sg13g2_decap_8
X_5939_ _0512_ net1281 net352 VPWR VGND sg13g2_nand2_1
XFILLER_31_44 VPWR VGND sg13g2_fill_2
XFILLER_31_88 VPWR VGND sg13g2_fill_2
Xoutput9 net9 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_0_221 VPWR VGND sg13g2_decap_8
XFILLER_1_744 VPWR VGND sg13g2_decap_8
XFILLER_49_737 VPWR VGND sg13g2_decap_8
XFILLER_48_247 VPWR VGND sg13g2_fill_1
XFILLER_45_921 VPWR VGND sg13g2_decap_8
XFILLER_45_998 VPWR VGND sg13g2_decap_8
XFILLER_44_464 VPWR VGND sg13g2_fill_1
XFILLER_16_133 VPWR VGND sg13g2_fill_2
XFILLER_44_486 VPWR VGND sg13g2_fill_2
XFILLER_13_851 VPWR VGND sg13g2_decap_4
XFILLER_40_681 VPWR VGND sg13g2_fill_2
XFILLER_12_361 VPWR VGND sg13g2_fill_2
X_6530__316 VPWR VGND net316 sg13g2_tiehi
X_4270_ net1103 _1791_ _1796_ VPWR VGND sg13g2_nor2_1
X_6708__124 VPWR VGND net124 sg13g2_tiehi
XFILLER_39_236 VPWR VGND sg13g2_decap_8
XFILLER_48_781 VPWR VGND sg13g2_decap_8
XFILLER_36_965 VPWR VGND sg13g2_decap_8
XFILLER_35_464 VPWR VGND sg13g2_fill_1
X_6773_ net241 VGND VPWR _0283_ s0.data_out\[1\]\[7\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_3985_ net1140 s0.data_out\[10\]\[5\] _1545_ VPWR VGND sg13g2_and2_1
X_5724_ VPWR _0021_ _0315_ VGND sg13g2_inv_1
X_5655_ _3049_ net1435 _3038_ VPWR VGND sg13g2_nand2_1
X_4606_ net1370 _2025_ _2103_ VPWR VGND sg13g2_nor2_1
Xhold310 s0.data_out\[6\]\[5\] VPWR VGND net630 sg13g2_dlygate4sd3_1
X_5586_ net1341 _2914_ _2990_ VPWR VGND sg13g2_nor2_1
Xhold321 _0018_ VPWR VGND net641 sg13g2_dlygate4sd3_1
Xhold343 s0.data_out\[2\]\[0\] VPWR VGND net663 sg13g2_dlygate4sd3_1
Xhold332 s0.data_out\[1\]\[0\] VPWR VGND net652 sg13g2_dlygate4sd3_1
X_4537_ s0.data_out\[6\]\[3\] s0.data_out\[5\]\[3\] net1081 _2036_ VPWR VGND sg13g2_mux2_1
X_4468_ _1941_ _1959_ _1976_ _1978_ _1979_ VPWR VGND sg13g2_or4_1
Xhold354 s0.data_out\[10\]\[2\] VPWR VGND net674 sg13g2_dlygate4sd3_1
Xhold365 _1210_ VPWR VGND net685 sg13g2_dlygate4sd3_1
Xhold376 _0054_ VPWR VGND net696 sg13g2_dlygate4sd3_1
Xhold387 s0.data_new_delayed\[7\] VPWR VGND net707 sg13g2_dlygate4sd3_1
X_6650__186 VPWR VGND net186 sg13g2_tiehi
X_3419_ VGND VPWR net1227 _1030_ _1033_ _1032_ sg13g2_a21oi_1
X_6207_ _0066_ _0752_ _0753_ _2802_ net1366 VPWR VGND sg13g2_a22oi_1
X_4399_ net1475 net339 _0202_ VPWR VGND sg13g2_and2_1
X_6138_ s0.data_out\[18\]\[0\] s0.data_out\[17\]\[0\] net1259 _0687_ VPWR VGND sg13g2_mux2_1
XFILLER_45_217 VPWR VGND sg13g2_decap_4
X_6069_ net1418 _0626_ _0630_ VPWR VGND sg13g2_nor2_1
XFILLER_27_921 VPWR VGND sg13g2_decap_4
XFILLER_26_55 VPWR VGND sg13g2_fill_2
XFILLER_26_66 VPWR VGND sg13g2_decap_8
XFILLER_42_957 VPWR VGND sg13g2_decap_8
XFILLER_42_32 VPWR VGND sg13g2_fill_2
XFILLER_41_478 VPWR VGND sg13g2_fill_2
XFILLER_6_803 VPWR VGND sg13g2_fill_2
XFILLER_21_191 VPWR VGND sg13g2_decap_8
XFILLER_3_15 VPWR VGND sg13g2_fill_2
XFILLER_49_501 VPWR VGND sg13g2_fill_1
XFILLER_3_59 VPWR VGND sg13g2_fill_2
XFILLER_1_596 VPWR VGND sg13g2_decap_4
XFILLER_49_534 VPWR VGND sg13g2_decap_8
XFILLER_37_707 VPWR VGND sg13g2_decap_4
XFILLER_36_206 VPWR VGND sg13g2_decap_8
XFILLER_18_987 VPWR VGND sg13g2_decap_8
XFILLER_32_445 VPWR VGND sg13g2_fill_1
XFILLER_33_979 VPWR VGND sg13g2_decap_8
X_3770_ VGND VPWR net1178 _1348_ _1349_ _1347_ sg13g2_a21oi_1
XFILLER_34_1012 VPWR VGND sg13g2_decap_8
X_6526__25 VPWR VGND net25 sg13g2_tiehi
XFILLER_8_162 VPWR VGND sg13g2_decap_8
XFILLER_8_140 VPWR VGND sg13g2_decap_8
X_5440_ VPWR _2858_ net453 VGND sg13g2_inv_1
X_5371_ VPWR _2789_ net424 VGND sg13g2_inv_1
X_4322_ VGND VPWR _1726_ _1844_ _1845_ net1115 sg13g2_a21oi_1
X_4253_ net1125 VPWR _1782_ VGND _1739_ _1781_ sg13g2_o21ai_1
X_4184_ _1719_ net1120 net654 VPWR VGND sg13g2_nand2_1
X_6721__110 VPWR VGND net110 sg13g2_tiehi
X_6756_ net72 VGND VPWR _0266_ s0.data_out\[2\]\[2\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_3968_ VPWR _0149_ _1532_ VGND sg13g2_inv_1
X_5707_ net1007 _2782_ _0302_ VPWR VGND sg13g2_nor2_1
X_6687_ net147 VGND VPWR net688 s0.data_out\[8\]\[5\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_12_13 VPWR VGND sg13g2_fill_2
X_3899_ _1463_ net1136 _1464_ _1465_ VPWR VGND sg13g2_a21o_1
X_5638_ _3032_ net1309 net519 VPWR VGND sg13g2_nand2_1
XFILLER_3_817 VPWR VGND sg13g2_decap_8
X_5569_ net1435 _2937_ _2975_ VPWR VGND sg13g2_nor2_1
Xhold151 _0209_ VPWR VGND net471 sg13g2_dlygate4sd3_1
Xhold140 _0010_ VPWR VGND net460 sg13g2_dlygate4sd3_1
XFILLER_2_338 VPWR VGND sg13g2_fill_1
Xhold162 s0.data_out\[16\]\[3\] VPWR VGND net482 sg13g2_dlygate4sd3_1
Xhold173 _0247_ VPWR VGND net493 sg13g2_dlygate4sd3_1
Xhold184 _0096_ VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold195 _0265_ VPWR VGND net515 sg13g2_dlygate4sd3_1
XFILLER_46_537 VPWR VGND sg13g2_fill_1
XFILLER_42_743 VPWR VGND sg13g2_fill_2
XFILLER_15_957 VPWR VGND sg13g2_decap_8
XFILLER_26_294 VPWR VGND sg13g2_decap_4
XFILLER_30_905 VPWR VGND sg13g2_fill_1
X_6523__28 VPWR VGND net28 sg13g2_tiehi
XFILLER_5_176 VPWR VGND sg13g2_fill_1
XFILLER_2_861 VPWR VGND sg13g2_decap_8
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_49_353 VPWR VGND sg13g2_decap_8
X_6705__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_18_762 VPWR VGND sg13g2_fill_1
X_4940_ s0.data_out\[3\]\[6\] s0.data_out\[2\]\[6\] net1046 _2403_ VPWR VGND sg13g2_mux2_1
X_4871_ VGND VPWR net995 _2307_ _2341_ net1359 sg13g2_a21oi_1
X_6610_ net230 VGND VPWR _0120_ s0.data_out\[14\]\[7\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_3822_ net1186 net1153 _1401_ VPWR VGND sg13g2_nor2b_1
X_6541_ net304 VGND VPWR _0051_ s0.genblk1\[18\].modules.bubble clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_3753_ net1183 _1329_ _1334_ VPWR VGND sg13g2_nor2_1
X_6472_ _0989_ VPWR _0990_ VGND net1477 net599 sg13g2_o21ai_1
X_3684_ VGND VPWR _1274_ _1264_ net1404 sg13g2_or2_1
X_5423_ VPWR _2841_ net536 VGND sg13g2_inv_1
X_5354_ _2772_ net712 VPWR VGND sg13g2_inv_2
X_4305_ _1828_ net632 net1118 VPWR VGND sg13g2_nand2b_1
X_5285_ _2711_ VPWR _2712_ VGND net1001 net1147 sg13g2_o21ai_1
X_4236_ net1122 VPWR _1769_ VGND _1695_ _1768_ sg13g2_o21ai_1
X_4167_ s0.data_out\[9\]\[0\] s0.data_out\[8\]\[0\] net1118 _1702_ VPWR VGND sg13g2_mux2_1
X_4098_ _1622_ _1644_ _1645_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_242 VPWR VGND sg13g2_fill_2
XFILLER_23_275 VPWR VGND sg13g2_fill_2
X_6739_ net90 VGND VPWR _0249_ s0.valid_out\[3\][0] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_23_89 VPWR VGND sg13g2_fill_1
Xfanout1404 net1406 net1404 VPWR VGND sg13g2_buf_8
Xfanout1426 net1429 net1426 VPWR VGND sg13g2_buf_8
Xfanout1448 ui_in[2] net1448 VPWR VGND sg13g2_buf_8
Xfanout1415 ui_in[6] net1415 VPWR VGND sg13g2_buf_8
Xfanout1437 net1438 net1437 VPWR VGND sg13g2_buf_8
Xfanout1459 net1460 net1459 VPWR VGND sg13g2_buf_8
XFILLER_47_857 VPWR VGND sg13g2_decap_8
XFILLER_46_367 VPWR VGND sg13g2_fill_2
XFILLER_46_378 VPWR VGND sg13g2_fill_1
XFILLER_30_779 VPWR VGND sg13g2_decap_8
XFILLER_7_953 VPWR VGND sg13g2_decap_8
XFILLER_6_496 VPWR VGND sg13g2_fill_2
X_5070_ _2518_ _2519_ _2521_ VPWR VGND _2520_ sg13g2_nand3b_1
XFILLER_49_150 VPWR VGND sg13g2_fill_1
X_4021_ _1568_ net1131 net572 VPWR VGND sg13g2_nand2_1
XFILLER_49_194 VPWR VGND sg13g2_fill_1
X_5972_ _0044_ _0539_ _0540_ _2788_ net1354 VPWR VGND sg13g2_a22oi_1
XFILLER_25_529 VPWR VGND sg13g2_fill_2
XFILLER_46_890 VPWR VGND sg13g2_decap_8
X_4923_ _2370_ _2384_ _2385_ _2386_ VPWR VGND sg13g2_nor3_1
XFILLER_33_573 VPWR VGND sg13g2_fill_2
XFILLER_20_201 VPWR VGND sg13g2_decap_8
X_4854_ VGND VPWR net995 _2270_ _2328_ net1358 sg13g2_a21oi_1
X_3805_ _1382_ net1182 _1383_ _1384_ VPWR VGND sg13g2_a21o_1
X_4785_ _2259_ VPWR _2260_ VGND net1057 _2873_ sg13g2_o21ai_1
X_6524_ net27 VGND VPWR _0034_ s0.data_out\[21\]\[5\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_3736_ _1281_ _1319_ net1486 _1320_ VPWR VGND sg13g2_nand3_1
XFILLER_20_278 VPWR VGND sg13g2_fill_2
X_6455_ net1367 _0898_ _0977_ VPWR VGND sg13g2_nor2_1
X_3667_ _1256_ VPWR _1257_ VGND _1247_ _1248_ sg13g2_o21ai_1
XFILLER_47_1011 VPWR VGND sg13g2_decap_8
X_3598_ net1203 net457 _1197_ VPWR VGND sg13g2_and2_1
X_5406_ VPWR _2824_ net647 VGND sg13g2_inv_1
X_6386_ _0911_ net1243 _0910_ VPWR VGND sg13g2_nand2b_1
XFILLER_0_628 VPWR VGND sg13g2_decap_8
X_5337_ _2755_ net1275 VPWR VGND sg13g2_inv_2
X_6510__42 VPWR VGND net42 sg13g2_tiehi
X_5268_ net386 net1024 net1019 _2695_ VPWR VGND sg13g2_a21o_1
X_4219_ VGND VPWR _1750_ _1752_ _1754_ net1433 sg13g2_a21oi_1
X_5199_ _2638_ net1006 _2637_ VPWR VGND sg13g2_nand2_1
XFILLER_29_835 VPWR VGND sg13g2_decap_8
XFILLER_16_518 VPWR VGND sg13g2_fill_2
XFILLER_34_66 VPWR VGND sg13g2_fill_2
XFILLER_4_901 VPWR VGND sg13g2_decap_8
XFILLER_4_978 VPWR VGND sg13g2_decap_8
Xfanout1223 net1231 net1223 VPWR VGND sg13g2_buf_2
Xfanout1201 net1202 net1201 VPWR VGND sg13g2_buf_2
Xfanout1212 s0.valid_out\[13\][0] net1212 VPWR VGND sg13g2_buf_8
Xfanout1234 net1235 net1234 VPWR VGND sg13g2_buf_8
Xfanout1256 net498 net1256 VPWR VGND sg13g2_buf_2
Xfanout1245 s0.valid_out\[16\][0] net1245 VPWR VGND sg13g2_buf_8
Xfanout1289 s0.shift_out\[20\][0] net1289 VPWR VGND sg13g2_buf_2
Xfanout1278 net1280 net1278 VPWR VGND sg13g2_buf_8
XFILLER_19_312 VPWR VGND sg13g2_decap_4
Xfanout1267 net1268 net1267 VPWR VGND sg13g2_buf_8
XFILLER_34_326 VPWR VGND sg13g2_fill_1
XFILLER_43_893 VPWR VGND sg13g2_fill_2
XFILLER_30_543 VPWR VGND sg13g2_decap_8
X_4570_ VGND VPWR net1088 _2066_ _2069_ _2068_ sg13g2_a21oi_1
X_3521_ VGND VPWR _1123_ _1122_ net1445 sg13g2_or2_1
X_6240_ net1478 VPWR _0780_ VGND _0777_ _0779_ sg13g2_o21ai_1
X_3452_ VGND VPWR net1216 _1064_ _1066_ _1065_ sg13g2_a21oi_1
X_6171_ VGND VPWR _0720_ _0710_ net1402 sg13g2_or2_1
X_5122_ _2566_ VPWR _2567_ VGND net1468 net576 sg13g2_o21ai_1
XFILLER_27_0 VPWR VGND sg13g2_fill_1
XFILLER_38_632 VPWR VGND sg13g2_fill_2
XFILLER_38_610 VPWR VGND sg13g2_fill_2
X_5053_ _2503_ VPWR _2504_ VGND _2492_ _2500_ sg13g2_o21ai_1
X_6646__191 VPWR VGND net191 sg13g2_tiehi
X_4004_ net1129 _1556_ _1561_ VPWR VGND sg13g2_nor2_1
XFILLER_37_186 VPWR VGND sg13g2_fill_2
X_5955_ VGND VPWR _0524_ _0526_ _0040_ _0527_ sg13g2_a21oi_1
X_5886_ VGND VPWR _0351_ _0458_ _0459_ net1293 sg13g2_a21oi_1
X_4906_ VGND VPWR net1048 _2366_ _2369_ _2368_ sg13g2_a21oi_1
XFILLER_34_893 VPWR VGND sg13g2_fill_1
X_4837_ s0.data_out\[4\]\[5\] s0.data_out\[3\]\[5\] net1059 _2312_ VPWR VGND sg13g2_mux2_1
X_4768_ _2246_ _2245_ net699 VPWR VGND sg13g2_nand2b_1
X_4699_ _2183_ _2184_ _2186_ VPWR VGND _2185_ sg13g2_nand3b_1
X_3719_ net1202 VPWR _1307_ VGND _1236_ _1306_ sg13g2_o21ai_1
X_6507_ net45 VGND VPWR net604 s0.data_out\[22\]\[0\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_6438_ _0963_ net1430 _0951_ VPWR VGND sg13g2_xnor2_1
XFILLER_1_926 VPWR VGND sg13g2_decap_8
X_6369_ s0.data_out\[16\]\[2\] s0.data_out\[15\]\[2\] net1232 _0894_ VPWR VGND sg13g2_mux2_1
XFILLER_49_919 VPWR VGND sg13g2_decap_8
Xhold11 s0.genblk1\[5\].modules.bubble VPWR VGND net331 sg13g2_dlygate4sd3_1
Xhold22 s0.genblk1\[12\].modules.bubble VPWR VGND net342 sg13g2_dlygate4sd3_1
Xhold44 s0.was_valid_out\[6\][0] VPWR VGND net364 sg13g2_dlygate4sd3_1
Xhold33 _0517_ VPWR VGND net353 sg13g2_dlygate4sd3_1
Xhold55 s0.data_out\[0\]\[1\] VPWR VGND net375 sg13g2_dlygate4sd3_1
XFILLER_29_66 VPWR VGND sg13g2_fill_1
Xhold77 s0.shift_out\[0\][0] VPWR VGND net397 sg13g2_dlygate4sd3_1
Xhold99 _0066_ VPWR VGND net419 sg13g2_dlygate4sd3_1
Xhold88 s0.data_out\[7\]\[1\] VPWR VGND net408 sg13g2_dlygate4sd3_1
Xhold66 s0.data_out\[0\]\[2\] VPWR VGND net386 sg13g2_dlygate4sd3_1
XFILLER_45_54 VPWR VGND sg13g2_fill_1
XFILLER_17_849 VPWR VGND sg13g2_fill_2
XFILLER_45_98 VPWR VGND sg13g2_decap_4
XFILLER_43_156 VPWR VGND sg13g2_fill_1
XFILLER_40_885 VPWR VGND sg13g2_decap_8
XFILLER_6_48 VPWR VGND sg13g2_fill_2
Xfanout1031 net710 net1031 VPWR VGND sg13g2_buf_8
XFILLER_6_1019 VPWR VGND sg13g2_decap_8
Xfanout1020 net1021 net1020 VPWR VGND sg13g2_buf_8
Xfanout1053 net1054 net1053 VPWR VGND sg13g2_buf_8
Xfanout1064 net1066 net1064 VPWR VGND sg13g2_buf_8
Xfanout1042 s0.shift_out\[2\][0] net1042 VPWR VGND sg13g2_buf_2
XFILLER_0_992 VPWR VGND sg13g2_decap_8
XFILLER_48_963 VPWR VGND sg13g2_decap_8
Xfanout1075 net384 net1075 VPWR VGND sg13g2_buf_8
Xfanout1097 net1104 net1097 VPWR VGND sg13g2_buf_8
XFILLER_19_120 VPWR VGND sg13g2_decap_4
Xfanout1086 net1087 net1086 VPWR VGND sg13g2_buf_1
X_5740_ _0326_ _0327_ _0328_ VPWR VGND sg13g2_nor2_1
X_5671_ VGND VPWR net1313 _3062_ _3065_ _3064_ sg13g2_a21oi_1
X_4622_ VGND VPWR net1078 net568 _2115_ _2082_ sg13g2_a21oi_1
X_4553_ _2033_ _2034_ _2042_ _2051_ _2052_ VPWR VGND sg13g2_nor4_1
XFILLER_7_591 VPWR VGND sg13g2_decap_4
X_3504_ VPWR _1109_ _1108_ VGND sg13g2_inv_1
X_4484_ net1086 s0.data_out\[6\]\[2\] _1992_ VPWR VGND sg13g2_and2_1
X_6223_ _0070_ _0764_ _0765_ _2798_ net1356 VPWR VGND sg13g2_a22oi_1
X_3435_ VGND VPWR net1229 _1046_ _1049_ _1048_ sg13g2_a21oi_1
X_6154_ VPWR VGND net1439 _0695_ _0702_ net1447 _0703_ _0678_ sg13g2_a221oi_1
X_6085_ net1266 net428 _0643_ VPWR VGND sg13g2_and2_1
X_5105_ net1027 s0.data_out\[1\]\[2\] _2553_ VPWR VGND sg13g2_and2_1
X_5036_ net1027 net1162 _2487_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_996 VPWR VGND sg13g2_decap_8
XFILLER_26_602 VPWR VGND sg13g2_fill_2
XFILLER_38_495 VPWR VGND sg13g2_fill_1
XFILLER_41_605 VPWR VGND sg13g2_decap_8
X_5938_ VGND VPWR net1295 _0508_ _0511_ _0510_ sg13g2_a21oi_1
XFILLER_13_329 VPWR VGND sg13g2_decap_8
XFILLER_15_57 VPWR VGND sg13g2_fill_2
XFILLER_22_830 VPWR VGND sg13g2_decap_4
X_5869_ _0445_ net1336 net1282 VPWR VGND sg13g2_nand2_1
XFILLER_31_56 VPWR VGND sg13g2_decap_4
XFILLER_1_723 VPWR VGND sg13g2_decap_8
XFILLER_49_716 VPWR VGND sg13g2_decap_8
XFILLER_45_900 VPWR VGND sg13g2_decap_8
XFILLER_45_977 VPWR VGND sg13g2_decap_8
XFILLER_9_867 VPWR VGND sg13g2_fill_1
XFILLER_48_760 VPWR VGND sg13g2_decap_8
X_6643__194 VPWR VGND net194 sg13g2_tiehi
X_6772_ net254 VGND VPWR _0282_ s0.data_out\[1\]\[6\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_3984_ _0153_ net611 _1544_ _2835_ net1386 VPWR VGND sg13g2_a22oi_1
X_5723_ _0314_ VPWR _0315_ VGND net1462 net635 sg13g2_o21ai_1
X_5654_ _3030_ _3031_ _3039_ _3047_ _3048_ VPWR VGND sg13g2_nor4_1
X_4605_ net1085 VPWR _2102_ VGND _2022_ _2101_ sg13g2_o21ai_1
X_5585_ net1325 VPWR _2989_ VGND _2917_ _2988_ sg13g2_o21ai_1
Xhold300 _0142_ VPWR VGND net620 sg13g2_dlygate4sd3_1
Xhold311 s0.data_out\[12\]\[4\] VPWR VGND net631 sg13g2_dlygate4sd3_1
Xhold344 s0.data_out\[17\]\[6\] VPWR VGND net664 sg13g2_dlygate4sd3_1
Xhold333 s0.data_out\[17\]\[0\] VPWR VGND net653 sg13g2_dlygate4sd3_1
Xhold322 s0.data_out\[4\]\[1\] VPWR VGND net642 sg13g2_dlygate4sd3_1
X_4536_ _2035_ net1080 net549 VPWR VGND sg13g2_nand2_1
Xhold355 s0.data_out\[9\]\[4\] VPWR VGND net675 sg13g2_dlygate4sd3_1
Xhold377 s0.data_out\[11\]\[6\] VPWR VGND net697 sg13g2_dlygate4sd3_1
X_4467_ _1978_ _1973_ _1977_ VPWR VGND sg13g2_nand2_1
Xhold366 s0.data_out\[13\]\[5\] VPWR VGND net686 sg13g2_dlygate4sd3_1
X_4398_ net1375 _1904_ _0201_ VPWR VGND sg13g2_nor2_1
X_3418_ VGND VPWR _0916_ _1031_ _1032_ net1227 sg13g2_a21oi_1
Xhold388 s0.data_new_delayed\[5\] VPWR VGND net708 sg13g2_dlygate4sd3_1
X_6206_ net1366 _0685_ _0753_ VPWR VGND sg13g2_nor2_1
X_6137_ VGND VPWR net1267 _0683_ _0686_ _0685_ sg13g2_a21oi_1
X_6068_ VGND VPWR _0629_ _0591_ net1437 sg13g2_or2_1
X_5019_ net1469 _2466_ _0261_ VPWR VGND sg13g2_and2_1
XFILLER_14_605 VPWR VGND sg13g2_fill_1
XFILLER_26_45 VPWR VGND sg13g2_fill_1
XFILLER_42_936 VPWR VGND sg13g2_decap_8
XFILLER_41_424 VPWR VGND sg13g2_fill_1
XFILLER_27_999 VPWR VGND sg13g2_decap_8
XFILLER_27_1020 VPWR VGND sg13g2_decap_8
XFILLER_49_513 VPWR VGND sg13g2_decap_8
XFILLER_1_575 VPWR VGND sg13g2_decap_8
XFILLER_17_454 VPWR VGND sg13g2_decap_8
XFILLER_18_966 VPWR VGND sg13g2_decap_8
X_6597__244 VPWR VGND net244 sg13g2_tiehi
XFILLER_33_958 VPWR VGND sg13g2_decap_8
XFILLER_41_980 VPWR VGND sg13g2_decap_8
X_5370_ VPWR _2788_ net628 VGND sg13g2_inv_1
X_4321_ _1844_ net555 net1120 VPWR VGND sg13g2_nand2b_1
XFILLER_5_892 VPWR VGND sg13g2_decap_8
X_4252_ net1000 _2849_ _1781_ VPWR VGND sg13g2_nor2_1
X_4183_ _1717_ VPWR _1718_ VGND _1708_ _1709_ sg13g2_o21ai_1
XFILLER_48_590 VPWR VGND sg13g2_decap_8
XFILLER_23_413 VPWR VGND sg13g2_fill_2
XFILLER_24_925 VPWR VGND sg13g2_decap_8
XFILLER_23_446 VPWR VGND sg13g2_decap_8
X_3967_ _1531_ VPWR _1532_ VGND net1488 net661 sg13g2_o21ai_1
X_6755_ net73 VGND VPWR net515 s0.data_out\[2\]\[1\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_5706_ _0017_ _0300_ _0301_ _2777_ net1342 VPWR VGND sg13g2_a22oi_1
X_6686_ net148 VGND VPWR net671 s0.data_out\[8\]\[4\] clknet_leaf_17_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_30_clk clknet_3_5__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_3898_ net1135 net1168 _1464_ VPWR VGND sg13g2_nor2b_1
X_5637_ net1449 _3023_ _3031_ VPWR VGND sg13g2_nor2_1
X_5568_ _2974_ _2973_ net1416 _2966_ net1426 VPWR VGND sg13g2_a22oi_1
Xhold130 _0234_ VPWR VGND net450 sg13g2_dlygate4sd3_1
X_4519_ net1479 _2014_ _0213_ VPWR VGND sg13g2_and2_1
Xhold152 s0.shift_out\[18\][0] VPWR VGND net472 sg13g2_dlygate4sd3_1
Xhold141 s0.data_out\[11\]\[3\] VPWR VGND net461 sg13g2_dlygate4sd3_1
Xhold185 s0.data_out\[9\]\[7\] VPWR VGND net505 sg13g2_dlygate4sd3_1
Xhold163 _0092_ VPWR VGND net483 sg13g2_dlygate4sd3_1
X_5499_ net412 net1328 _2905_ VPWR VGND sg13g2_nor2b_1
Xhold174 s0.data_out\[1\]\[1\] VPWR VGND net494 sg13g2_dlygate4sd3_1
Xhold196 s0.was_valid_out\[1\][0] VPWR VGND net516 sg13g2_dlygate4sd3_1
XFILLER_2_1022 VPWR VGND sg13g2_decap_8
XFILLER_42_733 VPWR VGND sg13g2_fill_1
XFILLER_18_1008 VPWR VGND sg13g2_decap_8
XFILLER_42_788 VPWR VGND sg13g2_decap_4
XFILLER_23_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_21_clk clknet_3_7__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_10_630 VPWR VGND sg13g2_fill_1
XFILLER_10_674 VPWR VGND sg13g2_fill_2
XFILLER_6_656 VPWR VGND sg13g2_fill_2
XFILLER_2_840 VPWR VGND sg13g2_decap_8
XFILLER_45_560 VPWR VGND sg13g2_decap_8
XFILLER_17_251 VPWR VGND sg13g2_fill_1
X_6640__197 VPWR VGND net197 sg13g2_tiehi
XFILLER_32_221 VPWR VGND sg13g2_fill_1
XFILLER_32_232 VPWR VGND sg13g2_fill_1
X_4870_ VGND VPWR net1050 net387 _2340_ _2302_ sg13g2_a21oi_1
X_3821_ s0.data_out\[12\]\[5\] s0.data_out\[11\]\[5\] net1188 _1400_ VPWR VGND sg13g2_mux2_1
X_6540_ net305 VGND VPWR _0050_ s0.valid_out\[19\][0] clknet_leaf_36_clk sg13g2_dfrbpq_1
XFILLER_20_449 VPWR VGND sg13g2_fill_1
XFILLER_32_298 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_12_clk clknet_3_3__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_3752_ _1331_ VPWR _1333_ VGND s0.was_valid_out\[11\][0] net1188 sg13g2_o21ai_1
X_6471_ _0988_ net1477 _0989_ VPWR VGND _0930_ sg13g2_nand3b_1
X_3683_ VGND VPWR _1273_ _1271_ net1413 sg13g2_or2_1
X_5422_ VPWR _2840_ net477 VGND sg13g2_inv_1
X_5353_ _2771_ net354 VPWR VGND sg13g2_inv_2
X_4304_ _1825_ net1099 _1826_ _1827_ VPWR VGND sg13g2_a21o_1
X_5284_ net394 net1025 net1023 _2711_ VPWR VGND sg13g2_a21o_1
X_4235_ net1000 _2853_ _1768_ VPWR VGND sg13g2_nor2_1
XFILLER_28_505 VPWR VGND sg13g2_fill_1
X_4166_ VGND VPWR net1122 _1698_ _1701_ _1700_ sg13g2_a21oi_1
X_4097_ _1638_ VPWR _1644_ VGND _1630_ _1641_ sg13g2_o21ai_1
X_4999_ _0257_ _2454_ _2455_ _2875_ net1360 VPWR VGND sg13g2_a22oi_1
XFILLER_11_416 VPWR VGND sg13g2_fill_1
X_6738_ net92 VGND VPWR _0248_ s0.was_valid_out\[3\][0] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_11_449 VPWR VGND sg13g2_decap_8
X_6669_ net166 VGND VPWR _0179_ s0.shift_out\[9\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_20_983 VPWR VGND sg13g2_decap_8
XFILLER_3_637 VPWR VGND sg13g2_decap_4
Xfanout1405 net1406 net1405 VPWR VGND sg13g2_buf_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
Xfanout1416 net1420 net1416 VPWR VGND sg13g2_buf_8
Xfanout1427 net1429 net1427 VPWR VGND sg13g2_buf_8
XFILLER_24_1012 VPWR VGND sg13g2_decap_8
Xfanout1438 ui_in[3] net1438 VPWR VGND sg13g2_buf_8
Xfanout1449 net1451 net1449 VPWR VGND sg13g2_buf_8
XFILLER_47_836 VPWR VGND sg13g2_decap_8
XFILLER_46_357 VPWR VGND sg13g2_fill_1
XFILLER_27_560 VPWR VGND sg13g2_decap_4
XFILLER_34_519 VPWR VGND sg13g2_fill_2
XFILLER_14_221 VPWR VGND sg13g2_decap_8
XFILLER_30_747 VPWR VGND sg13g2_fill_1
X_6594__247 VPWR VGND net247 sg13g2_tiehi
XFILLER_7_932 VPWR VGND sg13g2_decap_8
XFILLER_11_983 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_6_442 VPWR VGND sg13g2_fill_2
X_6711__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_9_1017 VPWR VGND sg13g2_decap_8
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_4020_ net1142 net1398 net1391 _0166_ VPWR VGND sg13g2_mux2_1
XFILLER_38_836 VPWR VGND sg13g2_fill_2
XFILLER_37_357 VPWR VGND sg13g2_decap_8
X_5971_ net1354 _0482_ _0540_ VPWR VGND sg13g2_nor2_1
X_4922_ VPWR VGND _2383_ net1461 _2381_ net1457 _2385_ _2377_ sg13g2_a221oi_1
XFILLER_20_224 VPWR VGND sg13g2_decap_8
X_4853_ VGND VPWR net1049 net540 _2327_ _2267_ sg13g2_a21oi_1
X_3804_ net1182 net1149 _1383_ VPWR VGND sg13g2_nor2b_1
X_4784_ _2259_ net1056 net400 VPWR VGND sg13g2_nand2_1
X_6523_ net28 VGND VPWR _0033_ s0.data_out\[21\]\[4\] clknet_leaf_1_clk sg13g2_dfrbpq_2
X_3735_ net1207 VPWR _1319_ VGND _1277_ _1318_ sg13g2_o21ai_1
X_6454_ net1242 VPWR _0976_ VGND _0895_ _0975_ sg13g2_o21ai_1
X_5405_ VPWR _2823_ net548 VGND sg13g2_inv_1
X_3666_ _1256_ _1255_ net1440 _1232_ net1445 VPWR VGND sg13g2_a22oi_1
X_3597_ _0114_ _1195_ _1196_ _2824_ net1378 VPWR VGND sg13g2_a22oi_1
X_6385_ VGND VPWR net1225 _0908_ _0910_ _0909_ sg13g2_a21oi_1
X_5336_ _2754_ net1031 VPWR VGND sg13g2_inv_2
XFILLER_0_607 VPWR VGND sg13g2_decap_8
X_5267_ VPWR VGND _2693_ net1458 _2692_ net1449 _2694_ _2691_ sg13g2_a221oi_1
X_4218_ _1750_ _1752_ net1433 _1753_ VPWR VGND sg13g2_nand3_1
XFILLER_29_814 VPWR VGND sg13g2_decap_8
X_5198_ s0.data_out\[0\]\[5\] s0.data_out\[1\]\[5\] net1034 _2637_ VPWR VGND sg13g2_mux2_1
X_4149_ VGND VPWR _1682_ _1685_ _0176_ _1686_ sg13g2_a21oi_1
XFILLER_18_46 VPWR VGND sg13g2_fill_2
Xclkload0 clknet_leaf_2_clk clkload0/Y VPWR VGND sg13g2_inv_4
XFILLER_4_957 VPWR VGND sg13g2_decap_8
XFILLER_3_445 VPWR VGND sg13g2_fill_1
XFILLER_3_434 VPWR VGND sg13g2_decap_8
XFILLER_3_423 VPWR VGND sg13g2_decap_4
Xfanout1213 net1215 net1213 VPWR VGND sg13g2_buf_8
Xfanout1202 net1203 net1202 VPWR VGND sg13g2_buf_1
Xfanout1224 net1231 net1224 VPWR VGND sg13g2_buf_1
Xfanout1235 net701 net1235 VPWR VGND sg13g2_buf_8
Xfanout1246 s0.valid_out\[16\][0] net1246 VPWR VGND sg13g2_buf_1
Xfanout1257 net1258 net1257 VPWR VGND sg13g2_buf_8
Xfanout1268 s0.shift_out\[18\][0] net1268 VPWR VGND sg13g2_buf_8
Xfanout1279 net1280 net1279 VPWR VGND sg13g2_buf_1
X_6780__130 VPWR VGND net130 sg13g2_tiehi
XFILLER_47_699 VPWR VGND sg13g2_fill_2
XFILLER_34_305 VPWR VGND sg13g2_fill_1
XFILLER_43_883 VPWR VGND sg13g2_decap_4
XFILLER_30_522 VPWR VGND sg13g2_fill_1
X_3520_ VGND VPWR net1216 _1119_ _1122_ _1121_ sg13g2_a21oi_1
XFILLER_7_795 VPWR VGND sg13g2_fill_1
X_3451_ net1216 net1159 _1065_ VPWR VGND sg13g2_nor2b_1
X_6170_ net1411 _0717_ _0719_ VPWR VGND sg13g2_nor2_1
X_5121_ _2565_ VPWR _2566_ VGND net1010 _2564_ sg13g2_o21ai_1
X_5052_ _2503_ net1436 _2499_ VPWR VGND sg13g2_nand2_1
X_4003_ _1558_ VPWR _1560_ VGND s0.was_valid_out\[9\][0] net1134 sg13g2_o21ai_1
XFILLER_26_806 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_20 VPWR VGND uio_out[5] sg13g2_tielo
X_5954_ VGND VPWR _0527_ net1329 net338 sg13g2_or2_1
X_5885_ _0458_ s0.data_out\[19\]\[2\] net1298 VPWR VGND sg13g2_nand2b_1
XFILLER_21_500 VPWR VGND sg13g2_fill_1
X_4905_ VGND VPWR _2251_ _2367_ _2368_ net1047 sg13g2_a21oi_1
X_4836_ _2311_ net1058 net601 VPWR VGND sg13g2_nand2_1
X_4767_ _2243_ _2244_ _2245_ VPWR VGND sg13g2_nor2_1
X_6506_ net46 VGND VPWR _0016_ s0.shift_out\[22\][0] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_21_599 VPWR VGND sg13g2_decap_8
X_4698_ net1400 _2182_ _2185_ VPWR VGND sg13g2_nor2_1
X_3718_ net1016 _2833_ _1306_ VPWR VGND sg13g2_nor2_1
X_6437_ _0961_ VPWR _0962_ VGND net1440 _0922_ sg13g2_o21ai_1
X_3649_ VGND VPWR _1124_ _1238_ _1239_ net1202 sg13g2_a21oi_1
XFILLER_20_58 VPWR VGND sg13g2_fill_1
XFILLER_1_905 VPWR VGND sg13g2_decap_8
X_6368_ _0893_ net1235 net420 VPWR VGND sg13g2_nand2_1
X_5319_ VPWR _2737_ net383 VGND sg13g2_inv_1
XFILLER_0_426 VPWR VGND sg13g2_fill_1
X_6299_ _0834_ net1236 _0835_ _0836_ VPWR VGND sg13g2_a21o_1
Xhold12 s0.genblk1\[21\].modules.bubble VPWR VGND net332 sg13g2_dlygate4sd3_1
Xhold23 s0.genblk1\[13\].modules.bubble VPWR VGND net343 sg13g2_dlygate4sd3_1
Xhold45 s0.shift_out\[14\][0] VPWR VGND net365 sg13g2_dlygate4sd3_1
Xhold34 s0.data_out\[23\]\[3\] VPWR VGND net354 sg13g2_dlygate4sd3_1
Xhold56 _0289_ VPWR VGND net376 sg13g2_dlygate4sd3_1
Xhold78 s0.shift_out\[23\][0] VPWR VGND net398 sg13g2_dlygate4sd3_1
Xhold89 _0205_ VPWR VGND net409 sg13g2_dlygate4sd3_1
XFILLER_28_121 VPWR VGND sg13g2_decap_4
XFILLER_28_132 VPWR VGND sg13g2_decap_4
Xhold67 s0.data_out\[3\]\[4\] VPWR VGND net387 sg13g2_dlygate4sd3_1
XFILLER_28_154 VPWR VGND sg13g2_fill_1
XFILLER_16_316 VPWR VGND sg13g2_decap_8
XFILLER_16_349 VPWR VGND sg13g2_fill_2
XFILLER_28_198 VPWR VGND sg13g2_fill_1
XFILLER_43_146 VPWR VGND sg13g2_fill_1
XFILLER_8_526 VPWR VGND sg13g2_fill_2
XFILLER_4_732 VPWR VGND sg13g2_decap_8
XFILLER_4_776 VPWR VGND sg13g2_decap_8
XFILLER_3_275 VPWR VGND sg13g2_decap_4
Xfanout1010 _2751_ net1010 VPWR VGND sg13g2_buf_8
Xfanout1021 net397 net1021 VPWR VGND sg13g2_buf_8
Xfanout1032 s0.shift_out\[1\][0] net1032 VPWR VGND sg13g2_buf_1
Xfanout1054 net1055 net1054 VPWR VGND sg13g2_buf_8
Xfanout1065 net1066 net1065 VPWR VGND sg13g2_buf_8
XFILLER_0_971 VPWR VGND sg13g2_decap_8
XFILLER_20_8 VPWR VGND sg13g2_fill_2
Xfanout1043 net1046 net1043 VPWR VGND sg13g2_buf_8
XFILLER_48_942 VPWR VGND sg13g2_decap_8
Xfanout1076 net1077 net1076 VPWR VGND sg13g2_buf_8
Xfanout1098 net1099 net1098 VPWR VGND sg13g2_buf_2
Xfanout1087 net1091 net1087 VPWR VGND sg13g2_buf_8
XFILLER_19_176 VPWR VGND sg13g2_fill_1
XFILLER_34_146 VPWR VGND sg13g2_decap_8
XFILLER_37_1022 VPWR VGND sg13g2_decap_8
X_5670_ VGND VPWR _2951_ _3063_ _3064_ net1313 sg13g2_a21oi_1
X_4621_ VPWR _0220_ _2114_ VGND sg13g2_inv_1
X_4552_ _2051_ net1335 _2049_ VPWR VGND sg13g2_xnor2_1
X_3503_ _1106_ _1107_ _1108_ VPWR VGND sg13g2_nor2_1
X_4483_ _0205_ _1990_ _1991_ _2859_ net1371 VPWR VGND sg13g2_a22oi_1
X_3434_ VGND VPWR _0925_ _1047_ _1048_ net1230 sg13g2_a21oi_1
X_6222_ net1356 net369 _0765_ VPWR VGND sg13g2_nor2_1
X_6153_ VGND VPWR net1267 _0699_ _0702_ _0701_ sg13g2_a21oi_1
X_6084_ _0054_ _0641_ _0642_ _2796_ net1355 VPWR VGND sg13g2_a22oi_1
X_5104_ _0265_ _2551_ _2552_ _2883_ net1348 VPWR VGND sg13g2_a22oi_1
X_5035_ s0.data_out\[2\]\[2\] s0.data_out\[1\]\[2\] net1033 _2486_ VPWR VGND sg13g2_mux2_1
XFILLER_39_975 VPWR VGND sg13g2_decap_8
XFILLER_25_113 VPWR VGND sg13g2_fill_1
XFILLER_14_809 VPWR VGND sg13g2_fill_2
XFILLER_26_658 VPWR VGND sg13g2_fill_1
XFILLER_41_639 VPWR VGND sg13g2_fill_1
XFILLER_40_105 VPWR VGND sg13g2_fill_1
X_5937_ VGND VPWR _0391_ _0509_ _0510_ net1295 sg13g2_a21oi_1
X_5868_ net1287 VPWR _0444_ VGND net1393 net1273 sg13g2_o21ai_1
X_4819_ _2294_ s0.data_out\[3\]\[6\] net1069 VPWR VGND sg13g2_nand2b_1
X_5799_ VGND VPWR _3059_ _0383_ _0384_ net1301 sg13g2_a21oi_1
XFILLER_5_529 VPWR VGND sg13g2_fill_1
XFILLER_1_702 VPWR VGND sg13g2_decap_8
XFILLER_1_779 VPWR VGND sg13g2_decap_8
XFILLER_45_956 VPWR VGND sg13g2_decap_8
XFILLER_29_496 VPWR VGND sg13g2_fill_2
XFILLER_16_146 VPWR VGND sg13g2_fill_2
XFILLER_32_628 VPWR VGND sg13g2_decap_4
XFILLER_9_802 VPWR VGND sg13g2_fill_1
XFILLER_12_363 VPWR VGND sg13g2_fill_1
XFILLER_40_683 VPWR VGND sg13g2_fill_1
XFILLER_12_374 VPWR VGND sg13g2_decap_8
XFILLER_8_367 VPWR VGND sg13g2_fill_1
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_39_205 VPWR VGND sg13g2_decap_8
X_6771_ net267 VGND VPWR _0281_ s0.data_out\[1\]\[5\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_5722_ _0313_ VPWR _0314_ VGND net1011 _0312_ sg13g2_o21ai_1
X_3983_ net1386 net374 _1544_ VPWR VGND sg13g2_nor2_1
XFILLER_31_672 VPWR VGND sg13g2_decap_8
X_5653_ _3047_ net1334 _3045_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_683 VPWR VGND sg13g2_fill_1
X_5584_ net1011 _2775_ _2988_ VPWR VGND sg13g2_nor2_1
X_4604_ net1074 s0.data_out\[5\]\[1\] _2101_ VPWR VGND sg13g2_and2_1
XFILLER_11_1025 VPWR VGND sg13g2_decap_4
Xhold301 s0.data_out\[12\]\[0\] VPWR VGND net621 sg13g2_dlygate4sd3_1
X_4535_ net1452 _2026_ _2034_ VPWR VGND sg13g2_nor2_1
Xhold334 s0.data_out\[8\]\[6\] VPWR VGND net654 sg13g2_dlygate4sd3_1
Xhold323 s0.data_out\[15\]\[4\] VPWR VGND net643 sg13g2_dlygate4sd3_1
Xhold312 s0.data_out\[7\]\[3\] VPWR VGND net632 sg13g2_dlygate4sd3_1
Xhold367 s0.data_out\[8\]\[5\] VPWR VGND net687 sg13g2_dlygate4sd3_1
X_4466_ _1974_ _1975_ _1977_ VPWR VGND sg13g2_nor2_1
Xhold378 s0.was_valid_out\[21\][0] VPWR VGND net698 sg13g2_dlygate4sd3_1
Xhold345 _0880_ VPWR VGND net665 sg13g2_dlygate4sd3_1
Xhold356 s0.data_out\[4\]\[2\] VPWR VGND net676 sg13g2_dlygate4sd3_1
X_4397_ VGND VPWR _1906_ _1909_ _0200_ _1910_ sg13g2_a21oi_1
X_3417_ _1031_ s0.data_out\[14\]\[3\] net1235 VPWR VGND sg13g2_nand2b_1
X_6205_ net1268 VPWR _0752_ VGND _0682_ _0751_ sg13g2_o21ai_1
Xhold389 s0.data_new_delayed\[6\] VPWR VGND net709 sg13g2_dlygate4sd3_1
X_6136_ VGND VPWR _0570_ _0684_ _0685_ net1267 sg13g2_a21oi_1
X_6067_ net1427 _0619_ _0628_ VPWR VGND sg13g2_nor2_1
X_5018_ VGND VPWR _2729_ _2466_ _0260_ _2471_ sg13g2_a21oi_1
XFILLER_26_13 VPWR VGND sg13g2_decap_8
XFILLER_27_978 VPWR VGND sg13g2_decap_8
XFILLER_42_915 VPWR VGND sg13g2_decap_8
XFILLER_13_127 VPWR VGND sg13g2_decap_4
XFILLER_10_889 VPWR VGND sg13g2_fill_2
XFILLER_3_17 VPWR VGND sg13g2_fill_1
XFILLER_1_554 VPWR VGND sg13g2_decap_8
XFILLER_49_569 VPWR VGND sg13g2_decap_8
XFILLER_44_241 VPWR VGND sg13g2_fill_2
XFILLER_45_786 VPWR VGND sg13g2_decap_8
XFILLER_32_414 VPWR VGND sg13g2_decap_8
XFILLER_32_425 VPWR VGND sg13g2_fill_2
XFILLER_32_458 VPWR VGND sg13g2_fill_1
XFILLER_40_480 VPWR VGND sg13g2_fill_1
X_4320_ _1841_ net1103 _1842_ _1843_ VPWR VGND sg13g2_a21o_1
XFILLER_4_370 VPWR VGND sg13g2_decap_8
X_4251_ VPWR _0184_ _1780_ VGND sg13g2_inv_1
X_4182_ _1717_ _1716_ net1442 _1693_ net1446 VPWR VGND sg13g2_a22oi_1
XFILLER_36_742 VPWR VGND sg13g2_decap_4
XFILLER_35_263 VPWR VGND sg13g2_decap_8
X_6765__49 VPWR VGND net49 sg13g2_tiehi
X_6754_ net74 VGND VPWR _0264_ s0.data_out\[2\]\[0\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_3966_ _1474_ _1530_ net1488 _1531_ VPWR VGND sg13g2_nand3_1
X_6685_ net149 VGND VPWR net638 s0.data_out\[8\]\[3\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5705_ VGND VPWR net1011 _3024_ _0301_ net1341 sg13g2_a21oi_1
XFILLER_32_992 VPWR VGND sg13g2_decap_8
X_5636_ VPWR VGND _3029_ net1458 _3025_ net1449 _3030_ _3023_ sg13g2_a221oi_1
X_3897_ _1462_ VPWR _1463_ VGND net1174 _2838_ sg13g2_o21ai_1
X_5567_ VGND VPWR net1323 _2972_ _2973_ _2969_ sg13g2_a21oi_1
X_4518_ VGND VPWR _2731_ _2014_ _0212_ _2019_ sg13g2_a21oi_1
Xhold131 s0.data_out\[11\]\[7\] VPWR VGND net451 sg13g2_dlygate4sd3_1
Xhold153 s0.data_out\[20\]\[7\] VPWR VGND net473 sg13g2_dlygate4sd3_1
X_5498_ net1462 net330 _0003_ VPWR VGND sg13g2_and2_1
Xhold120 s0.data_out\[18\]\[4\] VPWR VGND net440 sg13g2_dlygate4sd3_1
Xhold142 _0152_ VPWR VGND net462 sg13g2_dlygate4sd3_1
Xhold164 s0.data_out\[3\]\[7\] VPWR VGND net484 sg13g2_dlygate4sd3_1
X_4449_ s0.data_out\[7\]\[5\] s0.data_out\[6\]\[5\] net1095 _1960_ VPWR VGND sg13g2_mux2_1
Xhold186 s0.data_out\[19\]\[7\] VPWR VGND net506 sg13g2_dlygate4sd3_1
Xhold175 _0277_ VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold197 _0272_ VPWR VGND net517 sg13g2_dlygate4sd3_1
XFILLER_46_506 VPWR VGND sg13g2_decap_8
XFILLER_37_12 VPWR VGND sg13g2_fill_1
X_6119_ net1470 VPWR _0671_ VGND net543 _0665_ sg13g2_o21ai_1
XFILLER_2_1001 VPWR VGND sg13g2_decap_8
XFILLER_39_591 VPWR VGND sg13g2_fill_2
XFILLER_27_764 VPWR VGND sg13g2_fill_2
XFILLER_42_767 VPWR VGND sg13g2_fill_1
XFILLER_1_362 VPWR VGND sg13g2_fill_1
XFILLER_49_322 VPWR VGND sg13g2_decap_8
XFILLER_2_896 VPWR VGND sg13g2_decap_8
XFILLER_1_395 VPWR VGND sg13g2_fill_1
XFILLER_49_344 VPWR VGND sg13g2_decap_4
XFILLER_49_388 VPWR VGND sg13g2_decap_8
X_3820_ _1396_ _1398_ net1432 _1399_ VPWR VGND sg13g2_nand3_1
XFILLER_14_992 VPWR VGND sg13g2_decap_8
X_3751_ VGND VPWR net1015 _1218_ _1332_ _1331_ sg13g2_a21oi_1
X_6470_ net1240 VPWR _0988_ VGND _0927_ _0987_ sg13g2_o21ai_1
X_3682_ _1272_ _1271_ net1413 _1264_ net1404 VPWR VGND sg13g2_a22oi_1
X_5421_ VPWR _2839_ net489 VGND sg13g2_inv_1
X_5352_ VPWR _2770_ net586 VGND sg13g2_inv_1
X_4303_ net1099 net994 _1826_ VPWR VGND sg13g2_nor2_1
X_5283_ _2689_ VPWR _2710_ VGND _2708_ _2709_ sg13g2_o21ai_1
X_4234_ VPWR _0180_ _1767_ VGND sg13g2_inv_1
X_4165_ VGND VPWR _1568_ _1699_ _1700_ net1122 sg13g2_a21oi_1
X_4096_ _1604_ _1622_ _1639_ _1642_ _1643_ VPWR VGND sg13g2_or4_1
XFILLER_23_200 VPWR VGND sg13g2_fill_2
XFILLER_23_244 VPWR VGND sg13g2_fill_1
X_4998_ net1360 _2417_ _2455_ VPWR VGND sg13g2_nor2_1
XFILLER_17_1020 VPWR VGND sg13g2_decap_8
XFILLER_23_25 VPWR VGND sg13g2_decap_4
XFILLER_23_277 VPWR VGND sg13g2_fill_1
X_6737_ net93 VGND VPWR net493 s0.data_out\[4\]\[7\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_20_962 VPWR VGND sg13g2_decap_8
XFILLER_23_47 VPWR VGND sg13g2_decap_4
X_3949_ VGND VPWR _1393_ _1514_ _1515_ net1183 sg13g2_a21oi_1
X_6668_ net167 VGND VPWR _0178_ s0.genblk1\[8\].modules.bubble clknet_leaf_18_clk
+ sg13g2_dfrbpq_1
X_5619_ net1463 VPWR _3016_ VGND _3013_ _3015_ sg13g2_o21ai_1
X_6599_ net242 VGND VPWR _0109_ s0.was_valid_out\[14\][0] clknet_leaf_30_clk sg13g2_dfrbpq_1
Xfanout1417 net1420 net1417 VPWR VGND sg13g2_buf_1
Xfanout1428 net1429 net1428 VPWR VGND sg13g2_buf_1
X_6587__255 VPWR VGND net255 sg13g2_tiehi
Xfanout1406 ui_in[7] net1406 VPWR VGND sg13g2_buf_8
Xfanout1439 net1442 net1439 VPWR VGND sg13g2_buf_8
XFILLER_47_815 VPWR VGND sg13g2_decap_8
XFILLER_46_325 VPWR VGND sg13g2_decap_8
XFILLER_19_517 VPWR VGND sg13g2_fill_2
XFILLER_0_18 VPWR VGND sg13g2_decap_8
XFILLER_46_369 VPWR VGND sg13g2_fill_1
XFILLER_31_1006 VPWR VGND sg13g2_decap_8
X_6737__93 VPWR VGND net93 sg13g2_tiehi
XFILLER_7_911 VPWR VGND sg13g2_decap_8
XFILLER_11_962 VPWR VGND sg13g2_decap_8
XFILLER_6_432 VPWR VGND sg13g2_decap_4
XFILLER_7_988 VPWR VGND sg13g2_decap_8
XFILLER_2_693 VPWR VGND sg13g2_decap_8
XFILLER_49_185 VPWR VGND sg13g2_decap_8
XFILLER_37_325 VPWR VGND sg13g2_decap_4
X_5970_ net1293 VPWR _0539_ VGND _0479_ _0538_ sg13g2_o21ai_1
XFILLER_45_380 VPWR VGND sg13g2_decap_8
X_4921_ net1457 _2377_ _2384_ VPWR VGND sg13g2_nor2_1
X_4852_ net321 net1330 _2326_ _0239_ VPWR VGND sg13g2_nor3_1
XFILLER_33_542 VPWR VGND sg13g2_decap_8
X_3803_ s0.data_out\[12\]\[6\] s0.data_out\[11\]\[6\] net1188 _1382_ VPWR VGND sg13g2_mux2_1
XFILLER_33_575 VPWR VGND sg13g2_fill_1
X_4783_ VGND VPWR _2258_ _2257_ net1444 sg13g2_or2_1
X_6522_ net29 VGND VPWR net520 s0.data_out\[21\]\[3\] clknet_leaf_1_clk sg13g2_dfrbpq_2
X_3734_ net1194 s0.data_out\[12\]\[5\] _1318_ VPWR VGND sg13g2_and2_1
X_6453_ net1225 net420 _0975_ VPWR VGND sg13g2_and2_1
X_3665_ VGND VPWR net1204 _1252_ _1255_ _1254_ sg13g2_a21oi_1
X_5404_ VPWR _2822_ net602 VGND sg13g2_inv_1
X_3596_ net1378 _1129_ _1196_ VPWR VGND sg13g2_nor2_1
X_6384_ net1226 net1171 _0909_ VPWR VGND sg13g2_nor2b_1
X_5335_ _2753_ net1297 VPWR VGND sg13g2_inv_2
X_5266_ net1001 net547 net1024 _2693_ VPWR VGND sg13g2_nand3_1
X_4217_ _1752_ _1751_ net1125 VPWR VGND sg13g2_nand2b_1
X_5197_ VGND VPWR _2630_ _2635_ _2636_ net1426 sg13g2_a21oi_1
X_4148_ net1488 VPWR _1686_ VGND net666 _1680_ sg13g2_o21ai_1
XFILLER_18_58 VPWR VGND sg13g2_decap_8
X_4079_ VGND VPWR net1130 _1625_ _1626_ _1623_ sg13g2_a21oi_1
XFILLER_18_69 VPWR VGND sg13g2_decap_4
Xclkload1 VPWR clkload1/Y clknet_leaf_4_clk VGND sg13g2_inv_1
X_6734__96 VPWR VGND net96 sg13g2_tiehi
XFILLER_4_936 VPWR VGND sg13g2_decap_8
Xfanout1214 net1215 net1214 VPWR VGND sg13g2_buf_1
Xfanout1203 net1209 net1203 VPWR VGND sg13g2_buf_1
Xfanout1247 net1248 net1247 VPWR VGND sg13g2_buf_2
Xfanout1236 net1244 net1236 VPWR VGND sg13g2_buf_2
Xfanout1225 net1228 net1225 VPWR VGND sg13g2_buf_8
Xfanout1258 s0.valid_out\[17\][0] net1258 VPWR VGND sg13g2_buf_8
Xfanout1269 net1272 net1269 VPWR VGND sg13g2_buf_8
XFILLER_47_678 VPWR VGND sg13g2_decap_8
XFILLER_19_369 VPWR VGND sg13g2_fill_1
XFILLER_28_870 VPWR VGND sg13g2_decap_8
XFILLER_46_188 VPWR VGND sg13g2_decap_4
XFILLER_15_531 VPWR VGND sg13g2_decap_8
XFILLER_15_542 VPWR VGND sg13g2_fill_1
XFILLER_42_383 VPWR VGND sg13g2_decap_8
X_3450_ s0.data_out\[15\]\[4\] s0.data_out\[14\]\[4\] net1220 _1064_ VPWR VGND sg13g2_mux2_1
XFILLER_41_4 VPWR VGND sg13g2_fill_2
X_5120_ VGND VPWR net1010 _2533_ _2565_ net1349 sg13g2_a21oi_1
X_5051_ _2485_ _2493_ _2500_ _2501_ _2502_ VPWR VGND sg13g2_nor4_1
X_4002_ VGND VPWR net1013 _1446_ _1559_ _1558_ sg13g2_a21oi_1
XFILLER_38_634 VPWR VGND sg13g2_fill_1
Xheichips25_top_sorter_21 VPWR VGND uio_out[6] sg13g2_tielo
Xheichips25_top_sorter_10 VPWR VGND uio_oe[0] sg13g2_tielo
X_5953_ VPWR VGND _0525_ _0447_ _0504_ _0501_ _0526_ _0502_ sg13g2_a221oi_1
XFILLER_34_840 VPWR VGND sg13g2_fill_1
X_5884_ _0455_ net1276 _0456_ _0457_ VPWR VGND sg13g2_a21o_1
X_4904_ _2367_ s0.data_out\[2\]\[2\] net1056 VPWR VGND sg13g2_nand2b_1
XFILLER_34_884 VPWR VGND sg13g2_fill_2
XFILLER_21_534 VPWR VGND sg13g2_decap_8
XFILLER_21_545 VPWR VGND sg13g2_fill_1
X_4835_ net1437 _2280_ _2310_ VPWR VGND sg13g2_nor2_1
X_4766_ VGND VPWR net1338 net1069 _2244_ net1064 sg13g2_a21oi_1
X_6577__265 VPWR VGND net265 sg13g2_tiehi
X_6505_ net47 VGND VPWR _0015_ s0.genblk1\[21\].modules.bubble clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3717_ VPWR _0125_ _1305_ VGND sg13g2_inv_1
X_4697_ VGND VPWR _2184_ _2175_ net1410 sg13g2_or2_1
X_6436_ _0961_ net1421 _0959_ VPWR VGND sg13g2_nand2_1
X_3648_ _1238_ _2740_ net442 VPWR VGND sg13g2_nand2_1
X_6367_ net1484 net323 _0087_ VPWR VGND sg13g2_and2_1
X_3579_ _1181_ net1017 _1180_ VPWR VGND sg13g2_nand2_1
X_6731__99 VPWR VGND net99 sg13g2_tiehi
X_5318_ VPWR _2736_ net370 VGND sg13g2_inv_1
XFILLER_0_405 VPWR VGND sg13g2_decap_8
XFILLER_0_416 VPWR VGND sg13g2_fill_1
Xhold13 s0.module0.bubble VPWR VGND net333 sg13g2_dlygate4sd3_1
X_6298_ net1236 net1153 _0835_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_438 VPWR VGND sg13g2_decap_4
Xhold24 s0.genblk1\[7\].modules.bubble VPWR VGND net344 sg13g2_dlygate4sd3_1
X_5249_ VPWR _0282_ _2680_ VGND sg13g2_inv_1
X_6584__258 VPWR VGND net258 sg13g2_tiehi
Xhold46 s0.was_valid_out\[19\][0] VPWR VGND net366 sg13g2_dlygate4sd3_1
Xhold35 _2932_ VPWR VGND net355 sg13g2_dlygate4sd3_1
Xhold57 s0.data_out\[22\]\[7\] VPWR VGND net377 sg13g2_dlygate4sd3_1
Xhold79 _2995_ VPWR VGND net399 sg13g2_dlygate4sd3_1
XFILLER_21_1027 VPWR VGND sg13g2_fill_2
XFILLER_29_79 VPWR VGND sg13g2_decap_4
Xhold68 _2426_ VPWR VGND net388 sg13g2_dlygate4sd3_1
XFILLER_29_667 VPWR VGND sg13g2_fill_1
XFILLER_45_34 VPWR VGND sg13g2_fill_2
XFILLER_28_177 VPWR VGND sg13g2_decap_4
X_6701__132 VPWR VGND net132 sg13g2_tiehi
XFILLER_12_556 VPWR VGND sg13g2_decap_8
XFILLER_4_711 VPWR VGND sg13g2_decap_8
XFILLER_10_70 VPWR VGND sg13g2_fill_2
Xfanout1022 net1023 net1022 VPWR VGND sg13g2_buf_8
Xfanout1000 _2759_ net1000 VPWR VGND sg13g2_buf_8
XFILLER_0_950 VPWR VGND sg13g2_decap_8
Xfanout1011 _2749_ net1011 VPWR VGND sg13g2_buf_8
XFILLER_48_921 VPWR VGND sg13g2_decap_8
Xfanout1055 net585 net1055 VPWR VGND sg13g2_buf_8
Xfanout1044 net1046 net1044 VPWR VGND sg13g2_buf_1
Xfanout1033 net1035 net1033 VPWR VGND sg13g2_buf_8
Xfanout1088 net1090 net1088 VPWR VGND sg13g2_buf_8
Xfanout1077 net1079 net1077 VPWR VGND sg13g2_buf_2
Xfanout1066 net608 net1066 VPWR VGND sg13g2_buf_8
XFILLER_48_998 VPWR VGND sg13g2_decap_8
Xfanout1099 net1104 net1099 VPWR VGND sg13g2_buf_1
XFILLER_19_144 VPWR VGND sg13g2_fill_2
XFILLER_19_155 VPWR VGND sg13g2_fill_2
XFILLER_35_626 VPWR VGND sg13g2_decap_4
XFILLER_37_1001 VPWR VGND sg13g2_decap_8
XFILLER_43_670 VPWR VGND sg13g2_decap_4
XFILLER_31_810 VPWR VGND sg13g2_fill_2
XFILLER_34_169 VPWR VGND sg13g2_decap_8
X_4620_ _2113_ VPWR _2114_ VGND net1479 net669 sg13g2_o21ai_1
XFILLER_30_353 VPWR VGND sg13g2_fill_1
XFILLER_31_887 VPWR VGND sg13g2_fill_1
X_4551_ VGND VPWR _2050_ _2049_ net1335 sg13g2_or2_1
X_3502_ _2740_ net1395 _1107_ VPWR VGND sg13g2_nor2_1
X_4482_ net1371 _1923_ _1991_ VPWR VGND sg13g2_nor2_1
X_6221_ net1263 VPWR _0764_ VGND _0731_ _0763_ sg13g2_o21ai_1
X_3433_ _1047_ net545 net1234 VPWR VGND sg13g2_nand2b_1
X_6152_ VGND VPWR _0585_ _0700_ _0701_ net1267 sg13g2_a21oi_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_44_1016 VPWR VGND sg13g2_decap_8
X_5103_ net1348 _2477_ _2552_ VPWR VGND sg13g2_nor2_1
XFILLER_32_0 VPWR VGND sg13g2_decap_8
X_6083_ net1355 _0575_ _0642_ VPWR VGND sg13g2_nor2_1
XFILLER_39_954 VPWR VGND sg13g2_decap_8
X_5034_ VPWR VGND _2484_ net1458 _2480_ net1450 _2485_ _2478_ sg13g2_a221oi_1
XFILLER_25_147 VPWR VGND sg13g2_decap_4
X_5936_ _0509_ _2753_ net486 VPWR VGND sg13g2_nand2_1
XFILLER_25_169 VPWR VGND sg13g2_decap_4
X_5867_ _0036_ _0442_ _0443_ _2779_ net1344 VPWR VGND sg13g2_a22oi_1
X_4818_ _2291_ net1053 _2292_ _2293_ VPWR VGND sg13g2_a21o_1
X_5798_ _0383_ net432 net1308 VPWR VGND sg13g2_nand2b_1
XFILLER_22_898 VPWR VGND sg13g2_decap_8
X_4749_ VPWR _0232_ _2230_ VGND sg13g2_inv_1
X_6590__251 VPWR VGND net251 sg13g2_tiehi
X_6419_ _0940_ _0941_ _0939_ _0944_ VPWR VGND sg13g2_nand3_1
XFILLER_0_235 VPWR VGND sg13g2_decap_8
XFILLER_1_758 VPWR VGND sg13g2_decap_8
XFILLER_29_442 VPWR VGND sg13g2_decap_4
XFILLER_45_935 VPWR VGND sg13g2_decap_8
XFILLER_44_423 VPWR VGND sg13g2_fill_1
XFILLER_29_475 VPWR VGND sg13g2_decap_4
XFILLER_44_445 VPWR VGND sg13g2_fill_2
XFILLER_44_434 VPWR VGND sg13g2_fill_2
XFILLER_31_139 VPWR VGND sg13g2_fill_2
XFILLER_9_825 VPWR VGND sg13g2_fill_1
XFILLER_13_887 VPWR VGND sg13g2_fill_1
XFILLER_40_673 VPWR VGND sg13g2_decap_4
XFILLER_48_795 VPWR VGND sg13g2_decap_8
XFILLER_36_979 VPWR VGND sg13g2_decap_8
XFILLER_35_434 VPWR VGND sg13g2_fill_2
X_3982_ net1183 VPWR _1543_ VGND _1512_ _1542_ sg13g2_o21ai_1
X_6770_ net280 VGND VPWR _0280_ s0.data_out\[1\]\[4\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_5721_ VGND VPWR net1011 _3075_ _0313_ net1344 sg13g2_a21oi_1
X_5652_ VGND VPWR _3046_ _3045_ net1334 sg13g2_or2_1
XFILLER_11_1004 VPWR VGND sg13g2_decap_8
X_5583_ _0005_ _2986_ _2987_ _2778_ net1341 VPWR VGND sg13g2_a22oi_1
X_4603_ _0216_ _2099_ _2100_ _2864_ net1370 VPWR VGND sg13g2_a22oi_1
Xhold302 s0.data_out\[19\]\[6\] VPWR VGND net622 sg13g2_dlygate4sd3_1
X_4534_ VPWR VGND _2032_ net1460 _2028_ net1452 _2033_ _2026_ sg13g2_a221oi_1
Xhold335 _1897_ VPWR VGND net655 sg13g2_dlygate4sd3_1
Xhold313 s0.data_out\[20\]\[1\] VPWR VGND net633 sg13g2_dlygate4sd3_1
Xhold324 s0.was_valid_out\[11\][0] VPWR VGND net644 sg13g2_dlygate4sd3_1
Xhold346 s0.was_valid_out\[9\][0] VPWR VGND net666 sg13g2_dlygate4sd3_1
Xhold368 _0197_ VPWR VGND net688 sg13g2_dlygate4sd3_1
X_4465_ _1966_ VPWR _1976_ VGND net1442 _1940_ sg13g2_o21ai_1
Xhold357 s0.data_out\[1\]\[4\] VPWR VGND net677 sg13g2_dlygate4sd3_1
Xhold379 s0.was_valid_out\[4\][0] VPWR VGND net699 sg13g2_dlygate4sd3_1
X_4396_ net1482 VPWR _1910_ VGND net552 _1904_ sg13g2_o21ai_1
X_3416_ _1028_ net1213 _1029_ _1030_ VPWR VGND sg13g2_a21o_1
X_6204_ net1002 _2807_ _0751_ VPWR VGND sg13g2_nor2_1
X_6135_ _0684_ s0.data_out\[17\]\[1\] net1271 VPWR VGND sg13g2_nand2b_1
X_6066_ _0627_ _0626_ net1418 _0619_ net1427 VPWR VGND sg13g2_a22oi_1
X_5017_ net1468 VPWR _2471_ VGND _2468_ _2470_ sg13g2_o21ai_1
XFILLER_39_751 VPWR VGND sg13g2_decap_4
XFILLER_39_795 VPWR VGND sg13g2_fill_2
XFILLER_27_957 VPWR VGND sg13g2_decap_8
X_5919_ VGND VPWR net1287 _0489_ _0492_ _0491_ sg13g2_a21oi_1
XFILLER_42_57 VPWR VGND sg13g2_fill_1
XFILLER_22_684 VPWR VGND sg13g2_fill_2
XFILLER_1_533 VPWR VGND sg13g2_decap_8
XFILLER_49_548 VPWR VGND sg13g2_decap_8
XFILLER_18_902 VPWR VGND sg13g2_fill_2
XFILLER_29_272 VPWR VGND sg13g2_decap_8
XFILLER_45_765 VPWR VGND sg13g2_decap_8
X_6759__69 VPWR VGND net69 sg13g2_tiehi
X_6777__169 VPWR VGND net169 sg13g2_tiehi
XFILLER_13_673 VPWR VGND sg13g2_decap_8
XFILLER_34_1026 VPWR VGND sg13g2_fill_2
XFILLER_8_154 VPWR VGND sg13g2_decap_4
XFILLER_9_655 VPWR VGND sg13g2_fill_2
XFILLER_8_176 VPWR VGND sg13g2_decap_8
XFILLER_5_850 VPWR VGND sg13g2_fill_1
X_4250_ _1779_ VPWR _1780_ VGND net1489 net675 sg13g2_o21ai_1
XFILLER_4_382 VPWR VGND sg13g2_decap_8
X_4181_ VGND VPWR net1123 _1713_ _1716_ _1715_ sg13g2_a21oi_1
XFILLER_41_1008 VPWR VGND sg13g2_decap_8
XFILLER_35_242 VPWR VGND sg13g2_fill_1
X_6753_ net75 VGND VPWR _0263_ s0.shift_out\[2\][0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3965_ net1179 VPWR _1530_ VGND _1470_ _1529_ sg13g2_o21ai_1
X_5704_ net1317 VPWR _0300_ VGND _3026_ _0299_ sg13g2_o21ai_1
X_3896_ _1462_ net1174 net489 VPWR VGND sg13g2_nand2_1
X_6684_ net150 VGND VPWR _0194_ s0.data_out\[8\]\[2\] clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_32_971 VPWR VGND sg13g2_decap_8
X_5635_ _3029_ net1316 _3028_ VPWR VGND sg13g2_nand2b_1
XFILLER_12_38 VPWR VGND sg13g2_fill_2
Xhold110 s0.data_out\[15\]\[5\] VPWR VGND net430 sg13g2_dlygate4sd3_1
X_5566_ _2970_ net1311 _2971_ _2972_ VPWR VGND sg13g2_a21o_1
X_4517_ net1479 VPWR _2019_ VGND _2016_ _2018_ sg13g2_o21ai_1
Xhold132 _0156_ VPWR VGND net452 sg13g2_dlygate4sd3_1
X_5497_ net1340 _2898_ _0002_ VPWR VGND sg13g2_nor2_1
Xhold121 _0069_ VPWR VGND net441 sg13g2_dlygate4sd3_1
Xhold143 s0.data_out\[2\]\[3\] VPWR VGND net463 sg13g2_dlygate4sd3_1
Xhold165 _0259_ VPWR VGND net485 sg13g2_dlygate4sd3_1
X_4448_ _1958_ _1956_ _1959_ VPWR VGND _1957_ sg13g2_nand3b_1
Xhold154 _0048_ VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold176 s0.data_out\[20\]\[4\] VPWR VGND net496 sg13g2_dlygate4sd3_1
Xhold187 s0.data_out\[4\]\[6\] VPWR VGND net507 sg13g2_dlygate4sd3_1
Xhold198 s0.data_out\[8\]\[2\] VPWR VGND net518 sg13g2_dlygate4sd3_1
X_4379_ net1115 VPWR _1895_ VGND _1835_ _1894_ sg13g2_o21ai_1
X_6118_ _0668_ _0669_ _0670_ VPWR VGND sg13g2_nor2_1
X_6049_ VGND VPWR _0610_ _0600_ net1400 sg13g2_or2_1
XFILLER_18_209 VPWR VGND sg13g2_fill_1
XFILLER_15_927 VPWR VGND sg13g2_fill_2
X_6749__80 VPWR VGND net80 sg13g2_tiehi
XFILLER_10_654 VPWR VGND sg13g2_fill_2
XFILLER_6_636 VPWR VGND sg13g2_fill_1
XFILLER_6_658 VPWR VGND sg13g2_fill_1
XFILLER_6_647 VPWR VGND sg13g2_fill_2
XFILLER_2_875 VPWR VGND sg13g2_decap_8
X_6629__209 VPWR VGND net209 sg13g2_tiehi
XFILLER_49_301 VPWR VGND sg13g2_fill_1
XFILLER_49_367 VPWR VGND sg13g2_decap_4
XFILLER_45_540 VPWR VGND sg13g2_fill_2
XFILLER_17_242 VPWR VGND sg13g2_fill_2
XFILLER_14_971 VPWR VGND sg13g2_decap_8
X_3750_ _1329_ _1330_ _1331_ VPWR VGND sg13g2_nor2_1
X_3681_ VGND VPWR net1207 _1268_ _1271_ _1270_ sg13g2_a21oi_1
XFILLER_9_496 VPWR VGND sg13g2_fill_1
X_5420_ VPWR _2838_ net588 VGND sg13g2_inv_1
X_5351_ VPWR _2769_ net416 VGND sg13g2_inv_1
X_5282_ net1429 _2705_ _2709_ VPWR VGND sg13g2_and2_1
X_4302_ _1824_ VPWR _1825_ VGND net1106 _2851_ sg13g2_o21ai_1
XFILLER_4_61 VPWR VGND sg13g2_fill_1
X_4233_ _1766_ VPWR _1767_ VGND net1481 net596 sg13g2_o21ai_1
X_4164_ _1699_ _2747_ s0.data_out\[8\]\[1\] VPWR VGND sg13g2_nand2_1
X_4095_ VGND VPWR _1642_ _1641_ _1640_ sg13g2_or2_1
XFILLER_36_551 VPWR VGND sg13g2_fill_2
XFILLER_24_724 VPWR VGND sg13g2_fill_1
XFILLER_24_779 VPWR VGND sg13g2_fill_1
X_6736_ net94 VGND VPWR net508 s0.data_out\[4\]\[6\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_4997_ net1051 VPWR _2454_ VGND _2414_ _2453_ sg13g2_o21ai_1
X_3948_ _1514_ s0.data_out\[10\]\[4\] net1189 VPWR VGND sg13g2_nand2b_1
X_6746__83 VPWR VGND net83 sg13g2_tiehi
X_6667_ net168 VGND VPWR _0177_ s0.valid_out\[9\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3879_ net350 net1176 _1449_ VPWR VGND sg13g2_nor2_1
X_5618_ _3015_ _3012_ _3014_ VPWR VGND sg13g2_nand2_1
X_6598_ net243 VGND VPWR net562 s0.data_out\[15\]\[7\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_5549_ VGND VPWR net1323 _2954_ _2955_ _2950_ sg13g2_a21oi_1
Xfanout1418 net1420 net1418 VPWR VGND sg13g2_buf_8
Xfanout1429 ui_in[4] net1429 VPWR VGND sg13g2_buf_8
Xfanout1407 net1410 net1407 VPWR VGND sg13g2_buf_8
XFILLER_42_576 VPWR VGND sg13g2_decap_4
X_6635__202 VPWR VGND net202 sg13g2_tiehi
XFILLER_6_411 VPWR VGND sg13g2_fill_1
XFILLER_7_967 VPWR VGND sg13g2_decap_8
XFILLER_10_473 VPWR VGND sg13g2_decap_8
XFILLER_6_466 VPWR VGND sg13g2_fill_2
XFILLER_36_7 VPWR VGND sg13g2_fill_1
XFILLER_2_672 VPWR VGND sg13g2_decap_8
XFILLER_38_838 VPWR VGND sg13g2_fill_1
X_4920_ _2383_ _2382_ net1047 VPWR VGND sg13g2_nand2b_1
X_4851_ VPWR VGND _2301_ _2325_ _2324_ _2282_ _2326_ _2323_ sg13g2_a221oi_1
XFILLER_33_554 VPWR VGND sg13g2_fill_2
X_3802_ _1381_ net1188 s0.data_out\[11\]\[6\] VPWR VGND sg13g2_nand2_1
X_4782_ VGND VPWR net1060 _2254_ _2257_ _2256_ sg13g2_a21oi_1
X_6521_ net30 VGND VPWR _0031_ s0.data_out\[21\]\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_2
X_3733_ _0129_ _1316_ _1317_ _2826_ net1381 VPWR VGND sg13g2_a22oi_1
X_6452_ _0090_ _0973_ _0974_ _2813_ net1369 VPWR VGND sg13g2_a22oi_1
X_3664_ VGND VPWR _1139_ _1253_ _1254_ net1204 sg13g2_a21oi_1
X_5403_ _2821_ s0.data_out\[14\]\[4\] VPWR VGND sg13g2_inv_2
X_6743__86 VPWR VGND net86 sg13g2_tiehi
X_3595_ net1214 VPWR _1195_ VGND _1126_ _1194_ sg13g2_o21ai_1
X_6383_ s0.data_out\[16\]\[0\] s0.data_out\[15\]\[0\] net1232 _0908_ VPWR VGND sg13g2_mux2_1
XFILLER_47_1025 VPWR VGND sg13g2_decap_4
X_5334_ VPWR _2752_ net1305 VGND sg13g2_inv_1
X_5265_ _2692_ net1019 net1170 VPWR VGND sg13g2_nand2_1
X_4216_ _1624_ VPWR _1751_ VGND net1132 _2850_ sg13g2_o21ai_1
X_5196_ net1029 VPWR _2635_ VGND _2633_ _2634_ sg13g2_o21ai_1
X_4147_ _1683_ _1684_ _1685_ VPWR VGND sg13g2_nor2_1
XFILLER_44_808 VPWR VGND sg13g2_fill_1
X_4078_ s0.data_out\[10\]\[4\] s0.data_out\[9\]\[4\] net1134 _1625_ VPWR VGND sg13g2_mux2_1
XFILLER_37_871 VPWR VGND sg13g2_fill_2
XFILLER_43_329 VPWR VGND sg13g2_decap_4
XFILLER_37_893 VPWR VGND sg13g2_fill_1
XFILLER_12_716 VPWR VGND sg13g2_decap_8
XFILLER_12_738 VPWR VGND sg13g2_decap_8
XFILLER_24_576 VPWR VGND sg13g2_decap_4
XFILLER_11_226 VPWR VGND sg13g2_decap_8
XFILLER_11_237 VPWR VGND sg13g2_fill_1
XFILLER_7_219 VPWR VGND sg13g2_fill_1
X_6719_ net112 VGND VPWR _0229_ s0.data_out\[5\]\[1\] clknet_leaf_6_clk sg13g2_dfrbpq_2
Xclkload2 clknet_leaf_7_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_20_793 VPWR VGND sg13g2_decap_4
XFILLER_4_915 VPWR VGND sg13g2_decap_8
Xfanout1204 net1209 net1204 VPWR VGND sg13g2_buf_8
Xfanout1237 net1244 net1237 VPWR VGND sg13g2_buf_1
Xfanout1215 net1216 net1215 VPWR VGND sg13g2_buf_2
Xfanout1226 net1228 net1226 VPWR VGND sg13g2_buf_1
Xfanout1248 s0.valid_out\[16\][0] net1248 VPWR VGND sg13g2_buf_8
Xfanout1259 s0.valid_out\[17\][0] net1259 VPWR VGND sg13g2_buf_8
XFILLER_47_657 VPWR VGND sg13g2_decap_8
XFILLER_47_635 VPWR VGND sg13g2_decap_8
XFILLER_19_326 VPWR VGND sg13g2_decap_4
XFILLER_43_852 VPWR VGND sg13g2_fill_1
XFILLER_43_841 VPWR VGND sg13g2_decap_8
XFILLER_30_557 VPWR VGND sg13g2_decap_8
XFILLER_10_270 VPWR VGND sg13g2_decap_4
XFILLER_11_782 VPWR VGND sg13g2_decap_8
X_6740__89 VPWR VGND net89 sg13g2_tiehi
XFILLER_3_992 VPWR VGND sg13g2_decap_8
X_5050_ net1450 _2478_ _2501_ VPWR VGND sg13g2_nor2_1
X_4001_ _1556_ _1557_ _1558_ VPWR VGND sg13g2_nor2_1
XFILLER_37_101 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_22 VPWR VGND uio_out[7] sg13g2_tielo
Xheichips25_top_sorter_11 VPWR VGND uio_oe[1] sg13g2_tielo
X_5952_ _0519_ _0521_ _0525_ VPWR VGND sg13g2_nor2_1
X_4903_ _2364_ net1036 _2365_ _2366_ VPWR VGND sg13g2_a21o_1
X_5883_ net1276 net1162 _0456_ VPWR VGND sg13g2_nor2b_1
X_4834_ _2306_ _2308_ net1428 _2309_ VPWR VGND sg13g2_nand3_1
X_4765_ _2241_ _2242_ _2243_ VPWR VGND sg13g2_nor2_1
XFILLER_14_1013 VPWR VGND sg13g2_decap_8
X_6504_ net48 VGND VPWR _0014_ s0.valid_out\[22\][0] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3716_ _1304_ VPWR _1305_ VGND net1487 net679 sg13g2_o21ai_1
X_4696_ _2183_ _2182_ net1400 _2175_ net1409 VPWR VGND sg13g2_a22oi_1
X_6435_ net1421 _0959_ _0960_ VPWR VGND sg13g2_nor2_1
X_3647_ _1235_ net1191 _1236_ _1237_ VPWR VGND sg13g2_a21o_1
X_6366_ net1367 _0885_ _0886_ _0086_ VPWR VGND sg13g2_nor3_1
X_3578_ _1063_ VPWR _1180_ VGND net1221 _2826_ sg13g2_o21ai_1
X_5317_ VPWR _2735_ net362 VGND sg13g2_inv_1
Xhold14 s0.genblk1\[2\].modules.bubble VPWR VGND net334 sg13g2_dlygate4sd3_1
X_6297_ s0.data_out\[17\]\[5\] s0.data_out\[16\]\[5\] net1245 _0834_ VPWR VGND sg13g2_mux2_1
X_5248_ _2679_ VPWR _2680_ VGND net1467 net605 sg13g2_o21ai_1
Xhold25 s0.was_valid_out\[5\][0] VPWR VGND net345 sg13g2_dlygate4sd3_1
Xhold36 s0.was_valid_out\[2\][0] VPWR VGND net356 sg13g2_dlygate4sd3_1
Xhold47 _0049_ VPWR VGND net367 sg13g2_dlygate4sd3_1
X_5179_ s0.data_out\[0\]\[6\] s0.data_out\[1\]\[6\] net1034 _2618_ VPWR VGND sg13g2_mux2_1
Xhold58 _3057_ VPWR VGND net378 sg13g2_dlygate4sd3_1
XFILLER_21_1006 VPWR VGND sg13g2_decap_8
Xhold69 s0.data_out\[6\]\[3\] VPWR VGND net389 sg13g2_dlygate4sd3_1
XFILLER_28_145 VPWR VGND sg13g2_fill_2
XFILLER_29_679 VPWR VGND sg13g2_decap_8
XFILLER_43_115 VPWR VGND sg13g2_decap_8
XFILLER_24_351 VPWR VGND sg13g2_fill_2
XFILLER_8_528 VPWR VGND sg13g2_fill_1
XFILLER_3_211 VPWR VGND sg13g2_decap_8
XFILLER_3_244 VPWR VGND sg13g2_decap_4
XFILLER_3_233 VPWR VGND sg13g2_decap_8
Xfanout1001 _2758_ net1001 VPWR VGND sg13g2_buf_8
Xfanout1012 _2749_ net1012 VPWR VGND sg13g2_buf_8
XFILLER_48_900 VPWR VGND sg13g2_decap_8
Xfanout1045 net1046 net1045 VPWR VGND sg13g2_buf_8
Xfanout1034 net1035 net1034 VPWR VGND sg13g2_buf_8
Xfanout1023 net397 net1023 VPWR VGND sg13g2_buf_8
Xfanout1056 net1059 net1056 VPWR VGND sg13g2_buf_8
Xfanout1089 net1090 net1089 VPWR VGND sg13g2_buf_1
Xfanout1078 net1079 net1078 VPWR VGND sg13g2_buf_8
Xfanout1067 net1071 net1067 VPWR VGND sg13g2_buf_8
XFILLER_48_977 VPWR VGND sg13g2_decap_8
XFILLER_34_115 VPWR VGND sg13g2_decap_8
XFILLER_30_321 VPWR VGND sg13g2_decap_8
XFILLER_30_332 VPWR VGND sg13g2_decap_4
XFILLER_7_550 VPWR VGND sg13g2_fill_1
X_4550_ _2048_ VPWR _2049_ VGND net997 _2046_ sg13g2_o21ai_1
X_3501_ net1218 VPWR _1106_ VGND net1205 net1395 sg13g2_o21ai_1
X_4481_ net1096 VPWR _1990_ VGND _1920_ _1989_ sg13g2_o21ai_1
X_6220_ net1002 _2804_ _0763_ VPWR VGND sg13g2_nor2_1
X_3432_ _1044_ net1217 _1045_ _1046_ VPWR VGND sg13g2_a21o_1
X_6151_ _0700_ s0.data_out\[17\]\[3\] net1270 VPWR VGND sg13g2_nand2b_1
X_5102_ net1038 VPWR _2551_ VGND _2474_ _2550_ sg13g2_o21ai_1
X_6082_ net1279 VPWR _0641_ VGND _0572_ _0640_ sg13g2_o21ai_1
XFILLER_39_933 VPWR VGND sg13g2_decap_8
X_5033_ _2484_ net1038 _2483_ VPWR VGND sg13g2_nand2b_1
XFILLER_26_627 VPWR VGND sg13g2_fill_1
X_5935_ _0506_ net1277 _0507_ _0508_ VPWR VGND sg13g2_a21o_1
X_5866_ net1344 _0377_ _0443_ VPWR VGND sg13g2_nor2_1
X_4817_ net1053 net1148 _2292_ VPWR VGND sg13g2_nor2b_1
X_5797_ _0380_ net1286 _0381_ _0382_ VPWR VGND sg13g2_a21o_1
X_4748_ _2229_ VPWR _2230_ VGND net1474 net570 sg13g2_o21ai_1
X_4679_ _2147_ _2155_ _2163_ _2165_ _2166_ VPWR VGND sg13g2_nor4_1
X_6418_ _0943_ _0939_ _0940_ _0941_ VPWR VGND sg13g2_and3_1
X_6349_ _0878_ net1478 _0879_ VPWR VGND _0825_ sg13g2_nand3b_1
XFILLER_1_737 VPWR VGND sg13g2_decap_8
XFILLER_5_1011 VPWR VGND sg13g2_decap_8
XFILLER_45_914 VPWR VGND sg13g2_decap_8
XFILLER_16_148 VPWR VGND sg13g2_fill_1
XFILLER_25_671 VPWR VGND sg13g2_decap_8
XFILLER_24_170 VPWR VGND sg13g2_decap_8
XFILLER_25_682 VPWR VGND sg13g2_fill_2
XFILLER_9_815 VPWR VGND sg13g2_fill_1
XFILLER_12_354 VPWR VGND sg13g2_decap_8
XFILLER_13_855 VPWR VGND sg13g2_fill_1
XFILLER_13_866 VPWR VGND sg13g2_fill_1
XFILLER_9_859 VPWR VGND sg13g2_fill_2
XFILLER_8_347 VPWR VGND sg13g2_fill_2
XFILLER_4_531 VPWR VGND sg13g2_fill_2
XFILLER_21_81 VPWR VGND sg13g2_fill_1
X_6567__276 VPWR VGND net276 sg13g2_tiehi
XFILLER_48_774 VPWR VGND sg13g2_decap_8
XFILLER_36_958 VPWR VGND sg13g2_decap_8
XFILLER_16_660 VPWR VGND sg13g2_fill_1
X_3981_ net1140 net610 _1542_ VPWR VGND sg13g2_and2_1
X_5720_ VGND VPWR net1304 net609 _0312_ _3070_ sg13g2_a21oi_1
XFILLER_31_630 VPWR VGND sg13g2_decap_8
XFILLER_31_663 VPWR VGND sg13g2_decap_4
X_5651_ _3044_ VPWR _3045_ VGND net1011 _3042_ sg13g2_o21ai_1
XFILLER_30_162 VPWR VGND sg13g2_fill_1
X_6574__269 VPWR VGND net269 sg13g2_tiehi
X_5582_ net1341 _2922_ _2987_ VPWR VGND sg13g2_nor2_1
X_4602_ VGND VPWR net997 _2027_ _2100_ net1370 sg13g2_a21oi_1
X_4533_ _2032_ net1085 _2031_ VPWR VGND sg13g2_nand2b_1
Xhold303 _0658_ VPWR VGND net623 sg13g2_dlygate4sd3_1
Xhold314 _0042_ VPWR VGND net634 sg13g2_dlygate4sd3_1
Xhold325 _0144_ VPWR VGND net645 sg13g2_dlygate4sd3_1
Xhold358 s0.data_out\[3\]\[6\] VPWR VGND net678 sg13g2_dlygate4sd3_1
Xhold347 _0176_ VPWR VGND net667 sg13g2_dlygate4sd3_1
X_4464_ net1421 _1965_ _1975_ VPWR VGND sg13g2_nor2_1
Xhold369 s0.data_out\[17\]\[3\] VPWR VGND net689 sg13g2_dlygate4sd3_1
X_6203_ VPWR _0065_ _0750_ VGND sg13g2_inv_1
Xhold336 s0.data_out\[5\]\[1\] VPWR VGND net656 sg13g2_dlygate4sd3_1
X_4395_ _1907_ _1908_ _1909_ VPWR VGND sg13g2_nor2_1
X_3415_ net1213 net993 _1029_ VPWR VGND sg13g2_nor2_1
X_6134_ _0681_ net1253 _0682_ _0683_ VPWR VGND sg13g2_a21o_1
X_6065_ VGND VPWR net1274 _0623_ _0626_ _0625_ sg13g2_a21oi_1
X_5016_ _2470_ _2467_ _2469_ VPWR VGND sg13g2_nand2_1
XFILLER_39_785 VPWR VGND sg13g2_decap_4
XFILLER_41_438 VPWR VGND sg13g2_fill_2
X_5918_ VGND VPWR _0372_ _0490_ _0491_ net1287 sg13g2_a21oi_1
Xclkbuf_leaf_33_clk clknet_3_4__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
X_5849_ _0032_ _0428_ _0429_ _2781_ net1345 VPWR VGND sg13g2_a22oi_1
XFILLER_5_306 VPWR VGND sg13g2_fill_2
XFILLER_1_501 VPWR VGND sg13g2_fill_2
XFILLER_1_512 VPWR VGND sg13g2_decap_8
XFILLER_49_527 VPWR VGND sg13g2_decap_8
XFILLER_1_589 VPWR VGND sg13g2_decap_8
XFILLER_45_744 VPWR VGND sg13g2_fill_1
XFILLER_16_70 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_24_clk clknet_3_6__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_34_1005 VPWR VGND sg13g2_decap_8
XFILLER_41_994 VPWR VGND sg13g2_decap_8
XFILLER_9_634 VPWR VGND sg13g2_fill_2
X_4180_ VGND VPWR _1592_ _1714_ _1715_ net1123 sg13g2_a21oi_1
XFILLER_48_571 VPWR VGND sg13g2_fill_1
X_6580__262 VPWR VGND net262 sg13g2_tiehi
XFILLER_36_777 VPWR VGND sg13g2_fill_1
XFILLER_35_298 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_15_clk clknet_3_3__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_6752_ net76 VGND VPWR _0262_ s0.genblk1\[23\].modules.bubble clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3964_ net1135 s0.data_out\[10\]\[0\] _1529_ VPWR VGND sg13g2_and2_1
XFILLER_32_950 VPWR VGND sg13g2_decap_8
X_6758__70 VPWR VGND net70 sg13g2_tiehi
X_5703_ net1303 s0.data_out\[21\]\[0\] _0299_ VPWR VGND sg13g2_and2_1
X_6683_ net151 VGND VPWR _0193_ s0.data_out\[8\]\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3895_ VGND VPWR _1461_ _1460_ net1445 sg13g2_or2_1
X_5634_ VGND VPWR net1303 _3027_ _3028_ _3026_ sg13g2_a21oi_1
X_5565_ net1311 net1151 _2971_ VPWR VGND sg13g2_nor2b_1
Xhold100 s0.data_out\[15\]\[2\] VPWR VGND net420 sg13g2_dlygate4sd3_1
X_4516_ _2018_ _2015_ _2017_ VPWR VGND sg13g2_nand2_1
Xhold111 _0106_ VPWR VGND net431 sg13g2_dlygate4sd3_1
X_5496_ VGND VPWR _2900_ _2903_ _0001_ _2904_ sg13g2_a21oi_1
Xhold122 s0.data_out\[12\]\[1\] VPWR VGND net442 sg13g2_dlygate4sd3_1
Xhold133 s0.data_out\[7\]\[2\] VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold144 _0267_ VPWR VGND net464 sg13g2_dlygate4sd3_1
X_4447_ VGND VPWR _1958_ _1955_ net1402 sg13g2_or2_1
Xhold155 s0.data_out\[16\]\[5\] VPWR VGND net475 sg13g2_dlygate4sd3_1
Xhold177 _0045_ VPWR VGND net497 sg13g2_dlygate4sd3_1
Xhold166 s0.data_out\[19\]\[4\] VPWR VGND net486 sg13g2_dlygate4sd3_1
Xhold188 _0246_ VPWR VGND net508 sg13g2_dlygate4sd3_1
Xhold199 s0.data_out\[21\]\[3\] VPWR VGND net519 sg13g2_dlygate4sd3_1
X_4378_ net1103 s0.data_out\[7\]\[6\] _1894_ VPWR VGND sg13g2_and2_1
X_6117_ VGND VPWR _2737_ _2756_ _0669_ net1262 sg13g2_a21oi_1
X_7097_ s0.was_valid_out\[23\][0] net1 VPWR VGND sg13g2_buf_1
X_6048_ VGND VPWR _0609_ _0607_ net1409 sg13g2_or2_1
XFILLER_39_593 VPWR VGND sg13g2_fill_1
XFILLER_27_766 VPWR VGND sg13g2_fill_1
XFILLER_26_298 VPWR VGND sg13g2_fill_2
XFILLER_42_758 VPWR VGND sg13g2_decap_4
XFILLER_23_994 VPWR VGND sg13g2_decap_8
X_6764__62 VPWR VGND net62 sg13g2_tiehi
XFILLER_5_158 VPWR VGND sg13g2_fill_2
XFILLER_2_854 VPWR VGND sg13g2_decap_8
X_6564__279 VPWR VGND net279 sg13g2_tiehi
XFILLER_45_574 VPWR VGND sg13g2_fill_2
XFILLER_14_950 VPWR VGND sg13g2_decap_8
XFILLER_32_268 VPWR VGND sg13g2_decap_8
X_6755__73 VPWR VGND net73 sg13g2_tiehi
X_3680_ VGND VPWR _1155_ _1269_ _1270_ net1206 sg13g2_a21oi_1
X_5350_ _2768_ net1426 VPWR VGND sg13g2_inv_8
X_5281_ VGND VPWR _2699_ _2703_ _2708_ _2707_ sg13g2_a21oi_1
X_4301_ _1824_ net1106 s0.data_out\[7\]\[3\] VPWR VGND sg13g2_nand2_1
X_4232_ _1707_ _1765_ net1481 _1766_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_4_clk clknet_3_1__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ _1697_ net1111 _1695_ _1698_ VPWR VGND sg13g2_a21o_1
X_4094_ VGND VPWR _1635_ _1637_ _1641_ net1424 sg13g2_a21oi_1
XFILLER_28_519 VPWR VGND sg13g2_fill_1
XFILLER_49_891 VPWR VGND sg13g2_decap_8
XFILLER_36_541 VPWR VGND sg13g2_fill_1
XFILLER_24_736 VPWR VGND sg13g2_decap_4
X_4996_ net1040 net576 _2453_ VPWR VGND sg13g2_and2_1
X_6735_ net95 VGND VPWR _0245_ s0.data_out\[4\]\[5\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_3947_ _1511_ net1140 _1512_ _1513_ VPWR VGND sg13g2_a21o_1
X_6666_ net170 VGND VPWR net667 s0.was_valid_out\[9\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3878_ _1447_ VPWR _1448_ VGND net1185 _1330_ sg13g2_o21ai_1
X_5617_ net1012 VPWR _3014_ VGND s0.was_valid_out\[21\][0] net1318 sg13g2_o21ai_1
X_6597_ net244 VGND VPWR _0107_ s0.data_out\[15\]\[6\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_20_997 VPWR VGND sg13g2_decap_8
X_5548_ _2952_ net1311 _2953_ _2954_ VPWR VGND sg13g2_a21o_1
XFILLER_2_106 VPWR VGND sg13g2_fill_2
X_5479_ _2891_ VPWR net7 VGND _2767_ net991 sg13g2_o21ai_1
XFILLER_3_8 VPWR VGND sg13g2_fill_2
Xfanout1408 net1410 net1408 VPWR VGND sg13g2_buf_1
Xfanout1419 net1420 net1419 VPWR VGND sg13g2_buf_1
XFILLER_48_35 VPWR VGND sg13g2_decap_8
X_6628__210 VPWR VGND net210 sg13g2_tiehi
XFILLER_24_1026 VPWR VGND sg13g2_fill_2
XFILLER_19_519 VPWR VGND sg13g2_fill_1
XFILLER_15_736 VPWR VGND sg13g2_fill_2
XFILLER_30_717 VPWR VGND sg13g2_fill_2
XFILLER_22_290 VPWR VGND sg13g2_decap_8
X_6490__215 VPWR VGND net215 sg13g2_tiehi
XFILLER_7_946 VPWR VGND sg13g2_decap_8
XFILLER_11_997 VPWR VGND sg13g2_decap_8
X_6752__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_2_651 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_46_883 VPWR VGND sg13g2_decap_8
X_4850_ _2245_ VPWR _2325_ VGND _2297_ _2299_ sg13g2_o21ai_1
X_3801_ VGND VPWR net1195 _1377_ _1380_ _1379_ sg13g2_a21oi_1
X_6520_ net31 VGND VPWR net558 s0.data_out\[21\]\[1\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_4781_ VGND VPWR _2148_ _2255_ _2256_ net1060 sg13g2_a21oi_1
X_3732_ net1382 net415 _1317_ VPWR VGND sg13g2_nor2_1
X_6451_ net1369 _0906_ _0974_ VPWR VGND sg13g2_nor2_1
X_3663_ _1253_ _2740_ net467 VPWR VGND sg13g2_nand2_1
X_5402_ _2820_ net545 VPWR VGND sg13g2_inv_2
X_6382_ VGND VPWR net1242 _0904_ _0907_ _0906_ sg13g2_a21oi_1
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
X_5333_ _2751_ net1039 VPWR VGND sg13g2_inv_2
X_3594_ net1201 net481 _1194_ VPWR VGND sg13g2_and2_1
X_5264_ _2690_ VPWR _2691_ VGND net1001 net1166 sg13g2_o21ai_1
X_4215_ _1750_ net1125 _1749_ VPWR VGND sg13g2_nand2b_1
X_5195_ net1019 net1156 _2634_ VPWR VGND sg13g2_nor2b_1
X_4146_ VGND VPWR _2732_ _2747_ _1684_ net1125 sg13g2_a21oi_1
X_4077_ _1624_ net1132 s0.data_out\[9\]\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_34_37 VPWR VGND sg13g2_fill_2
X_4979_ VPWR _0252_ _2440_ VGND sg13g2_inv_1
X_6718_ net113 VGND VPWR _0228_ s0.data_out\[5\]\[0\] clknet_leaf_5_clk sg13g2_dfrbpq_2
Xclkload3 VPWR clkload3/Y clknet_leaf_6_clk VGND sg13g2_inv_1
XFILLER_20_772 VPWR VGND sg13g2_decap_8
XFILLER_20_783 VPWR VGND sg13g2_decap_8
X_6649_ net187 VGND VPWR _0159_ s0.data_new_delayed\[0\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_3_415 VPWR VGND sg13g2_fill_2
Xfanout1205 net1208 net1205 VPWR VGND sg13g2_buf_8
Xfanout1227 net1228 net1227 VPWR VGND sg13g2_buf_8
Xfanout1216 net365 net1216 VPWR VGND sg13g2_buf_8
Xfanout1238 net1239 net1238 VPWR VGND sg13g2_buf_2
Xfanout1249 net1251 net1249 VPWR VGND sg13g2_buf_8
XFILLER_46_102 VPWR VGND sg13g2_fill_2
XFILLER_19_316 VPWR VGND sg13g2_fill_2
XFILLER_43_820 VPWR VGND sg13g2_fill_2
XFILLER_27_382 VPWR VGND sg13g2_fill_2
XFILLER_7_765 VPWR VGND sg13g2_fill_2
XFILLER_3_971 VPWR VGND sg13g2_decap_8
X_4000_ net1396 _2747_ _1557_ VPWR VGND sg13g2_nor2_1
Xheichips25_top_sorter_12 VPWR VGND uio_oe[3] sg13g2_tielo
X_5951_ _0504_ _0519_ _0485_ _0524_ VPWR VGND _0523_ sg13g2_nand4_1
X_4902_ net1036 net1163 _2365_ VPWR VGND sg13g2_nor2b_1
X_5882_ s0.data_out\[20\]\[2\] s0.data_out\[19\]\[2\] net1283 _0455_ VPWR VGND sg13g2_mux2_1
X_4833_ _2308_ net996 _2307_ VPWR VGND sg13g2_nand2_1
X_4764_ net1397 _2748_ _2242_ VPWR VGND sg13g2_nor2_1
X_6503_ net50 VGND VPWR net393 s0.was_valid_out\[22\][0] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3715_ _1246_ _1303_ net1484 _1304_ VPWR VGND sg13g2_nand3_1
X_4695_ VGND VPWR net1076 _2179_ _2182_ _2181_ sg13g2_a21oi_1
X_6434_ VGND VPWR net1241 _0956_ _0959_ _0958_ sg13g2_a21oi_1
X_3646_ net1191 net1168 _1236_ VPWR VGND sg13g2_nor2b_1
X_6365_ VGND VPWR _2736_ _0887_ _0085_ _0892_ sg13g2_a21oi_1
X_3577_ VGND VPWR net1204 _1178_ _1179_ _1176_ sg13g2_a21oi_1
X_6296_ _0833_ net1248 net475 VPWR VGND sg13g2_nand2_1
XFILLER_1_919 VPWR VGND sg13g2_decap_8
X_5316_ VPWR _2734_ net348 VGND sg13g2_inv_1
X_5247_ _2678_ VPWR _2679_ VGND net1006 _2677_ sg13g2_o21ai_1
Xhold26 _0224_ VPWR VGND net346 sg13g2_dlygate4sd3_1
Xhold37 _0260_ VPWR VGND net357 sg13g2_dlygate4sd3_1
Xhold15 s0.genblk1\[23\].modules.bubble VPWR VGND net335 sg13g2_dlygate4sd3_1
X_5178_ _2615_ net1031 _2616_ _2617_ VPWR VGND sg13g2_a21o_1
Xhold48 s0.data_out\[17\]\[5\] VPWR VGND net368 sg13g2_dlygate4sd3_1
Xhold59 s0.data_out\[23\]\[0\] VPWR VGND net379 sg13g2_dlygate4sd3_1
X_6625__213 VPWR VGND net213 sg13g2_tiehi
X_4129_ _1669_ VPWR _1670_ VGND net1491 net613 sg13g2_o21ai_1
XFILLER_43_138 VPWR VGND sg13g2_fill_1
XFILLER_25_831 VPWR VGND sg13g2_decap_8
X_6632__206 VPWR VGND net206 sg13g2_tiehi
XFILLER_4_746 VPWR VGND sg13g2_decap_8
XFILLER_3_267 VPWR VGND sg13g2_decap_4
Xfanout1013 _2746_ net1013 VPWR VGND sg13g2_buf_8
XFILLER_3_289 VPWR VGND sg13g2_fill_2
Xfanout1002 _2757_ net1002 VPWR VGND sg13g2_buf_8
Xfanout1046 net396 net1046 VPWR VGND sg13g2_buf_8
Xfanout1024 net1026 net1024 VPWR VGND sg13g2_buf_8
Xfanout1035 s0.valid_out\[1\][0] net1035 VPWR VGND sg13g2_buf_8
Xfanout1079 s0.shift_out\[5\][0] net1079 VPWR VGND sg13g2_buf_1
XFILLER_0_985 VPWR VGND sg13g2_decap_8
Xfanout1057 net1059 net1057 VPWR VGND sg13g2_buf_8
Xfanout1068 net1071 net1068 VPWR VGND sg13g2_buf_8
XFILLER_48_956 VPWR VGND sg13g2_decap_8
XFILLER_19_146 VPWR VGND sg13g2_fill_1
XFILLER_47_499 VPWR VGND sg13g2_decap_4
XFILLER_31_812 VPWR VGND sg13g2_fill_1
XFILLER_35_91 VPWR VGND sg13g2_fill_2
X_3500_ _0108_ _1104_ _1105_ _2814_ net1380 VPWR VGND sg13g2_a22oi_1
XFILLER_11_591 VPWR VGND sg13g2_fill_1
X_4480_ net997 _2863_ _1989_ VPWR VGND sg13g2_nor2_1
X_3431_ net1217 net1150 _1045_ VPWR VGND sg13g2_nor2b_1
X_6150_ _0697_ net1253 _0698_ _0699_ VPWR VGND sg13g2_a21o_1
X_5101_ net1004 _2884_ _2550_ VPWR VGND sg13g2_nor2_1
X_6081_ net1266 net418 _0640_ VPWR VGND sg13g2_and2_1
X_5032_ VGND VPWR net1027 _2482_ _2483_ _2481_ sg13g2_a21oi_1
XFILLER_39_989 VPWR VGND sg13g2_decap_8
XFILLER_38_466 VPWR VGND sg13g2_fill_1
XFILLER_26_617 VPWR VGND sg13g2_fill_1
X_5934_ net1277 net1156 _0507_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_801 VPWR VGND sg13g2_fill_1
X_5865_ net1301 VPWR _0442_ VGND _0374_ _0441_ sg13g2_o21ai_1
XFILLER_22_834 VPWR VGND sg13g2_fill_1
XFILLER_34_672 VPWR VGND sg13g2_fill_1
X_4816_ s0.data_out\[4\]\[6\] s0.data_out\[3\]\[6\] net1058 _2291_ VPWR VGND sg13g2_mux2_1
X_5796_ net1286 net1147 _0381_ VPWR VGND sg13g2_nor2b_1
X_4747_ _2193_ _2228_ net1474 _2229_ VPWR VGND sg13g2_nand3_1
X_4678_ _2164_ VPWR _2165_ VGND net1452 _2140_ sg13g2_o21ai_1
X_6417_ VPWR _0942_ _0941_ VGND sg13g2_inv_1
X_3629_ VGND VPWR _1222_ _1221_ _1219_ sg13g2_or2_1
X_6348_ net1250 VPWR _0878_ VGND _0822_ _0877_ sg13g2_o21ai_1
XFILLER_1_716 VPWR VGND sg13g2_decap_8
XFILLER_49_709 VPWR VGND sg13g2_decap_8
X_6279_ _0814_ net1236 _0815_ _0816_ VPWR VGND sg13g2_a21o_1
XFILLER_13_845 VPWR VGND sg13g2_fill_1
XFILLER_12_388 VPWR VGND sg13g2_fill_2
XFILLER_0_782 VPWR VGND sg13g2_decap_8
XFILLER_48_753 VPWR VGND sg13g2_decap_8
XFILLER_35_436 VPWR VGND sg13g2_fill_1
X_3980_ _0152_ _1540_ _1541_ _2836_ net1384 VPWR VGND sg13g2_a22oi_1
XFILLER_44_981 VPWR VGND sg13g2_decap_8
X_5650_ _3044_ _2749_ _3043_ VPWR VGND sg13g2_nand2_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_4601_ net1085 VPWR _2099_ VGND _2029_ _2098_ sg13g2_o21ai_1
X_5581_ net1326 VPWR _2986_ VGND _2925_ _2985_ sg13g2_o21ai_1
X_4532_ VGND VPWR net1075 _2030_ _2031_ _2029_ sg13g2_a21oi_1
X_4463_ VGND VPWR _1970_ _1972_ _1974_ net1431 sg13g2_a21oi_1
Xhold315 s0.data_out\[22\]\[4\] VPWR VGND net635 sg13g2_dlygate4sd3_1
Xhold326 s0.data_out\[22\]\[2\] VPWR VGND net646 sg13g2_dlygate4sd3_1
Xhold304 s0.data_out\[21\]\[2\] VPWR VGND net624 sg13g2_dlygate4sd3_1
Xhold348 s0.data_out\[17\]\[4\] VPWR VGND net668 sg13g2_dlygate4sd3_1
X_3414_ _1027_ VPWR _1028_ VGND net1219 _2816_ sg13g2_o21ai_1
Xhold337 s0.data_out\[19\]\[2\] VPWR VGND net657 sg13g2_dlygate4sd3_1
X_6202_ _0749_ VPWR _0750_ VGND net1471 net660 sg13g2_o21ai_1
Xhold359 s0.data_out\[13\]\[0\] VPWR VGND net679 sg13g2_dlygate4sd3_1
X_4394_ VGND VPWR _2731_ _2760_ _1908_ net1100 sg13g2_a21oi_1
X_6133_ net1253 net1169 _0682_ VPWR VGND sg13g2_nor2b_1
X_6064_ VGND VPWR _0512_ _0624_ _0625_ net1275 sg13g2_a21oi_1
X_5015_ net1010 VPWR _2469_ VGND s0.was_valid_out\[1\][0] net1045 sg13g2_o21ai_1
XFILLER_39_797 VPWR VGND sg13g2_fill_1
XFILLER_38_285 VPWR VGND sg13g2_fill_1
XFILLER_42_929 VPWR VGND sg13g2_decap_8
XFILLER_35_981 VPWR VGND sg13g2_decap_8
X_5917_ _0490_ s0.data_out\[19\]\[7\] net1296 VPWR VGND sg13g2_nand2b_1
X_5848_ net1345 _0364_ _0429_ VPWR VGND sg13g2_nor2_1
X_5779_ VGND VPWR _3032_ _0363_ _0364_ net1305 sg13g2_a21oi_1
XFILLER_49_506 VPWR VGND sg13g2_decap_8
XFILLER_1_568 VPWR VGND sg13g2_decap_8
XFILLER_27_1013 VPWR VGND sg13g2_decap_8
XFILLER_29_263 VPWR VGND sg13g2_decap_4
XFILLER_17_425 VPWR VGND sg13g2_fill_2
XFILLER_18_959 VPWR VGND sg13g2_decap_8
XFILLER_26_992 VPWR VGND sg13g2_decap_8
XFILLER_41_973 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_9_646 VPWR VGND sg13g2_fill_2
XFILLER_5_841 VPWR VGND sg13g2_decap_8
X_6573__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_5_885 VPWR VGND sg13g2_decap_8
XFILLER_48_583 VPWR VGND sg13g2_decap_8
XFILLER_17_992 VPWR VGND sg13g2_decap_8
X_6751_ net77 VGND VPWR _0261_ s0.valid_out\[2\][0] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_3963_ VGND VPWR _1523_ _1527_ _0148_ _1528_ sg13g2_a21oi_1
X_5702_ VGND VPWR _3090_ _0297_ _0016_ _0298_ sg13g2_a21oi_1
X_6682_ net152 VGND VPWR _0192_ s0.data_out\[8\]\[0\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3894_ VGND VPWR net1181 _1457_ _1460_ _1459_ sg13g2_a21oi_1
X_5633_ s0.data_out\[22\]\[0\] s0.data_out\[21\]\[0\] net1310 _3027_ VPWR VGND sg13g2_mux2_1
X_5564_ s0.data_out\[23\]\[5\] s0.data_out\[22\]\[5\] net1318 _2970_ VPWR VGND sg13g2_mux2_1
X_4515_ net998 VPWR _2017_ VGND net345 net1094 sg13g2_o21ai_1
Xhold101 _0103_ VPWR VGND net421 sg13g2_dlygate4sd3_1
Xhold112 s0.data_out\[20\]\[6\] VPWR VGND net432 sg13g2_dlygate4sd3_1
X_5495_ net1463 VPWR _2904_ VGND net559 _2898_ sg13g2_o21ai_1
Xhold123 _0137_ VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold134 _0206_ VPWR VGND net454 sg13g2_dlygate4sd3_1
X_4446_ net1411 _1948_ _1957_ VPWR VGND sg13g2_nor2_1
Xhold156 _0094_ VPWR VGND net476 sg13g2_dlygate4sd3_1
Xhold167 _0057_ VPWR VGND net487 sg13g2_dlygate4sd3_1
Xhold145 s0.data_out\[9\]\[2\] VPWR VGND net465 sg13g2_dlygate4sd3_1
Xhold189 s0.data_out\[9\]\[6\] VPWR VGND net509 sg13g2_dlygate4sd3_1
X_4377_ _0197_ _1892_ _1893_ _2849_ net1375 VPWR VGND sg13g2_a22oi_1
Xhold178 s0.shift_out\[17\][0] VPWR VGND net498 sg13g2_dlygate4sd3_1
X_6116_ net1249 _0662_ _0668_ VPWR VGND sg13g2_nor2_1
X_6047_ _0608_ _0607_ net1409 _0600_ net1400 VPWR VGND sg13g2_a22oi_1
XFILLER_39_583 VPWR VGND sg13g2_fill_1
XFILLER_2_1015 VPWR VGND sg13g2_decap_8
XFILLER_27_756 VPWR VGND sg13g2_fill_2
XFILLER_27_778 VPWR VGND sg13g2_decap_4
XFILLER_23_940 VPWR VGND sg13g2_decap_8
XFILLER_23_951 VPWR VGND sg13g2_fill_2
XFILLER_22_450 VPWR VGND sg13g2_fill_1
XFILLER_23_973 VPWR VGND sg13g2_decap_8
X_6557__287 VPWR VGND net287 sg13g2_tiehi
XFILLER_5_126 VPWR VGND sg13g2_fill_2
XFILLER_2_833 VPWR VGND sg13g2_decap_8
XFILLER_49_336 VPWR VGND sg13g2_decap_4
XFILLER_18_723 VPWR VGND sg13g2_fill_2
XFILLER_45_553 VPWR VGND sg13g2_decap_8
XFILLER_45_542 VPWR VGND sg13g2_fill_1
XFILLER_17_244 VPWR VGND sg13g2_fill_1
XFILLER_13_483 VPWR VGND sg13g2_decap_4
XFILLER_40_291 VPWR VGND sg13g2_fill_1
X_4300_ _1807_ VPWR _1823_ VGND net1456 _1814_ sg13g2_o21ai_1
X_5280_ _2706_ VPWR _2707_ VGND net1435 _2702_ sg13g2_o21ai_1
X_4231_ net1122 VPWR _1765_ VGND _1703_ _1764_ sg13g2_o21ai_1
X_4162_ _1696_ VPWR _1697_ VGND net1118 _2843_ sg13g2_o21ai_1
XFILLER_49_870 VPWR VGND sg13g2_decap_8
X_4093_ VGND VPWR _1627_ _1629_ _1640_ net1433 sg13g2_a21oi_1
XFILLER_36_553 VPWR VGND sg13g2_fill_1
X_4995_ _0256_ _2451_ _2452_ _2876_ net1360 VPWR VGND sg13g2_a22oi_1
X_3946_ net1140 net1158 _1512_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_770 VPWR VGND sg13g2_decap_8
X_6734_ net96 VGND VPWR _0244_ s0.data_out\[4\]\[4\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_6665_ net171 VGND VPWR _0175_ s0.data_out\[10\]\[7\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_20_976 VPWR VGND sg13g2_decap_8
X_3877_ _1447_ _1446_ _1445_ VPWR VGND sg13g2_nand2b_1
X_5616_ net1302 _3009_ _3013_ VPWR VGND sg13g2_nor2_1
X_6596_ net245 VGND VPWR net431 s0.data_out\[15\]\[5\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_5547_ net1311 net1147 _2953_ VPWR VGND sg13g2_nor2b_1
X_5478_ _2891_ net1416 net991 VPWR VGND sg13g2_nand2_1
X_4429_ VGND VPWR net1097 _1937_ _1940_ _1939_ sg13g2_a21oi_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
Xfanout1409 net1410 net1409 VPWR VGND sg13g2_buf_8
XFILLER_24_1005 VPWR VGND sg13g2_decap_8
XFILLER_47_829 VPWR VGND sg13g2_decap_8
XFILLER_39_391 VPWR VGND sg13g2_decap_4
XFILLER_15_748 VPWR VGND sg13g2_fill_2
XFILLER_23_781 VPWR VGND sg13g2_fill_1
XFILLER_7_925 VPWR VGND sg13g2_decap_8
XFILLER_6_402 VPWR VGND sg13g2_decap_8
XFILLER_11_976 VPWR VGND sg13g2_decap_8
X_6570__273 VPWR VGND net273 sg13g2_tiehi
XFILLER_38_807 VPWR VGND sg13g2_fill_2
XFILLER_37_306 VPWR VGND sg13g2_fill_2
XFILLER_46_862 VPWR VGND sg13g2_decap_8
XFILLER_45_394 VPWR VGND sg13g2_decap_8
XFILLER_21_707 VPWR VGND sg13g2_fill_1
X_3800_ VGND VPWR _1258_ _1378_ _1379_ net1195 sg13g2_a21oi_1
X_4780_ _2255_ net434 net1067 VPWR VGND sg13g2_nand2b_1
XFILLER_14_770 VPWR VGND sg13g2_fill_1
X_3731_ net1205 VPWR _1316_ VGND _1285_ _1315_ sg13g2_o21ai_1
Xclkload10 clkload10/Y clknet_leaf_21_clk VPWR VGND sg13g2_inv_2
X_6450_ net1242 VPWR _0973_ VGND _0903_ _0972_ sg13g2_o21ai_1
X_3662_ _1250_ net1193 _1251_ _1252_ VPWR VGND sg13g2_a21o_1
X_5401_ _2819_ net612 VPWR VGND sg13g2_inv_2
X_6381_ VGND VPWR _0790_ _0905_ _0906_ net1239 sg13g2_a21oi_1
X_3593_ VPWR _0113_ net592 VGND sg13g2_inv_1
XFILLER_6_991 VPWR VGND sg13g2_decap_8
X_5332_ _2750_ net1328 VPWR VGND sg13g2_inv_2
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_5263_ net375 net1024 net1019 _2690_ VPWR VGND sg13g2_a21o_1
X_4214_ VGND VPWR net1116 _1747_ _1749_ _1748_ sg13g2_a21oi_1
X_5194_ VGND VPWR _2631_ _2632_ _2633_ net1001 sg13g2_a21oi_1
X_4145_ net1116 _1677_ _1683_ VPWR VGND sg13g2_nor2_1
X_4076_ net1130 net1159 _1623_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_350 VPWR VGND sg13g2_fill_1
XFILLER_24_545 VPWR VGND sg13g2_decap_4
XFILLER_12_707 VPWR VGND sg13g2_decap_4
X_4978_ _2439_ VPWR _2440_ VGND net1473 net540 sg13g2_o21ai_1
Xclkload4 VPWR clkload4/Y clknet_leaf_14_clk VGND sg13g2_inv_1
X_3929_ net1138 net1149 _1495_ VPWR VGND sg13g2_nor2b_1
X_6717_ net114 VGND VPWR _0227_ s0.shift_out\[5\][0] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_6648_ net188 VGND VPWR _0158_ s0.valid_out\[10\][0] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_6579_ net263 VGND VPWR _0089_ s0.data_out\[16\]\[0\] clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_8_1010 VPWR VGND sg13g2_decap_8
Xfanout1217 net1218 net1217 VPWR VGND sg13g2_buf_8
Xfanout1228 net1231 net1228 VPWR VGND sg13g2_buf_8
Xfanout1206 net1208 net1206 VPWR VGND sg13g2_buf_2
Xfanout1239 net1244 net1239 VPWR VGND sg13g2_buf_1
XFILLER_27_350 VPWR VGND sg13g2_fill_2
XFILLER_27_361 VPWR VGND sg13g2_decap_8
XFILLER_28_884 VPWR VGND sg13g2_fill_2
XFILLER_43_887 VPWR VGND sg13g2_fill_1
XFILLER_43_876 VPWR VGND sg13g2_decap_8
XFILLER_42_397 VPWR VGND sg13g2_decap_4
XFILLER_24_71 VPWR VGND sg13g2_decap_8
XFILLER_3_950 VPWR VGND sg13g2_decap_8
XFILLER_37_147 VPWR VGND sg13g2_decap_4
Xheichips25_top_sorter_13 VPWR VGND uio_oe[4] sg13g2_tielo
X_5950_ _0520_ _0521_ _0522_ _0523_ VPWR VGND sg13g2_nor3_1
XFILLER_19_862 VPWR VGND sg13g2_decap_8
X_4901_ s0.data_out\[3\]\[2\] s0.data_out\[2\]\[2\] net1043 _2364_ VPWR VGND sg13g2_mux2_1
XFILLER_34_854 VPWR VGND sg13g2_decap_4
X_5881_ _0454_ net1284 net657 VPWR VGND sg13g2_nand2_1
X_4832_ _2188_ VPWR _2307_ VGND net1067 _2876_ sg13g2_o21ai_1
X_4763_ net1064 VPWR _2241_ VGND net1393 net1054 sg13g2_o21ai_1
X_4694_ VGND VPWR _2056_ _2180_ _2181_ net1076 sg13g2_a21oi_1
X_6502_ net51 VGND VPWR net439 s0.data_out\[23\]\[7\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_6618__221 VPWR VGND net221 sg13g2_tiehi
X_3714_ net1202 VPWR _1303_ VGND _1242_ _1302_ sg13g2_o21ai_1
X_6433_ VGND VPWR _0833_ _0957_ _0958_ net1241 sg13g2_a21oi_1
X_3645_ _1234_ VPWR _1235_ VGND net1197 _2829_ sg13g2_o21ai_1
X_6364_ net1477 VPWR _0892_ VGND _0889_ _0891_ sg13g2_o21ai_1
X_3576_ _1177_ VPWR _1178_ VGND net1210 _2821_ sg13g2_o21ai_1
X_6295_ _0828_ _0829_ _0827_ _0832_ VPWR VGND sg13g2_nand3_1
X_5315_ VPWR _2733_ net350 VGND sg13g2_inv_1
X_5246_ VGND VPWR _2754_ _2618_ _2678_ net1347 sg13g2_a21oi_1
Xhold38 s0.was_valid_out\[8\][0] VPWR VGND net358 sg13g2_dlygate4sd3_1
Xhold16 s0.genblk1\[9\].modules.bubble VPWR VGND net336 sg13g2_dlygate4sd3_1
Xhold27 s0.shift_out\[21\][0] VPWR VGND net347 sg13g2_dlygate4sd3_1
X_5177_ net1031 _2612_ _2616_ VPWR VGND sg13g2_nor2_1
Xhold49 _0734_ VPWR VGND net369 sg13g2_dlygate4sd3_1
XFILLER_28_114 VPWR VGND sg13g2_decap_8
X_4128_ _1668_ VPWR _1669_ VGND net1013 _1667_ sg13g2_o21ai_1
XFILLER_28_125 VPWR VGND sg13g2_fill_2
XFILLER_28_136 VPWR VGND sg13g2_fill_1
XFILLER_28_147 VPWR VGND sg13g2_fill_1
X_4059_ s0.data_out\[10\]\[7\] s0.data_out\[9\]\[7\] net1134 _1606_ VPWR VGND sg13g2_mux2_1
XFILLER_37_692 VPWR VGND sg13g2_fill_2
XFILLER_25_843 VPWR VGND sg13g2_fill_2
X_6775__203 VPWR VGND net203 sg13g2_tiehi
XFILLER_24_331 VPWR VGND sg13g2_fill_2
XFILLER_40_824 VPWR VGND sg13g2_decap_4
XFILLER_12_526 VPWR VGND sg13g2_fill_2
XFILLER_25_898 VPWR VGND sg13g2_fill_2
XFILLER_8_519 VPWR VGND sg13g2_decap_8
XFILLER_20_570 VPWR VGND sg13g2_fill_2
XFILLER_4_725 VPWR VGND sg13g2_decap_8
XFILLER_3_279 VPWR VGND sg13g2_fill_1
Xfanout1003 _2755_ net1003 VPWR VGND sg13g2_buf_8
Xfanout1025 net1026 net1025 VPWR VGND sg13g2_buf_8
Xfanout1014 _2746_ net1014 VPWR VGND sg13g2_buf_8
XFILLER_0_964 VPWR VGND sg13g2_decap_8
Xfanout1036 net1042 net1036 VPWR VGND sg13g2_buf_2
Xfanout1047 net1055 net1047 VPWR VGND sg13g2_buf_8
XFILLER_48_935 VPWR VGND sg13g2_decap_8
Xfanout1058 net1059 net1058 VPWR VGND sg13g2_buf_8
Xfanout1069 net1071 net1069 VPWR VGND sg13g2_buf_8
XFILLER_37_1015 VPWR VGND sg13g2_decap_8
XFILLER_30_301 VPWR VGND sg13g2_decap_8
XFILLER_30_378 VPWR VGND sg13g2_fill_1
XFILLER_7_530 VPWR VGND sg13g2_fill_2
X_3430_ s0.data_out\[15\]\[6\] s0.data_out\[14\]\[6\] net1221 _1044_ VPWR VGND sg13g2_mux2_1
X_6080_ VPWR _0053_ net598 VGND sg13g2_inv_1
X_5100_ VPWR _0264_ _2549_ VGND sg13g2_inv_1
X_5031_ s0.data_out\[2\]\[0\] s0.data_out\[1\]\[0\] net1035 _2482_ VPWR VGND sg13g2_mux2_1
XFILLER_39_968 VPWR VGND sg13g2_decap_8
XFILLER_47_990 VPWR VGND sg13g2_decap_8
X_5933_ _0505_ VPWR _0506_ VGND net1283 _2787_ sg13g2_o21ai_1
XFILLER_18_180 VPWR VGND sg13g2_fill_1
X_5864_ net1286 net473 _0441_ VPWR VGND sg13g2_and2_1
XFILLER_33_150 VPWR VGND sg13g2_fill_2
XFILLER_34_695 VPWR VGND sg13g2_decap_8
X_4815_ _2290_ net1058 net678 VPWR VGND sg13g2_nand2_1
X_5795_ s0.data_out\[21\]\[6\] s0.data_out\[20\]\[6\] net1296 _0380_ VPWR VGND sg13g2_mux2_1
X_4746_ net1073 VPWR _2228_ VGND _2187_ _2227_ sg13g2_o21ai_1
X_4677_ _2152_ _2154_ net1447 _2164_ VPWR VGND sg13g2_nand3_1
X_6416_ VGND VPWR _0941_ _0938_ net1402 sg13g2_or2_1
X_3628_ net348 net1198 _1221_ VPWR VGND sg13g2_nor2_1
X_6347_ net1237 s0.data_out\[16\]\[6\] _0877_ VPWR VGND sg13g2_and2_1
X_3559_ VGND VPWR s0.shift_out\[14\][0] _1158_ _1161_ _1160_ sg13g2_a21oi_1
X_6278_ net1236 net1144 _0815_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_249 VPWR VGND sg13g2_decap_4
X_5229_ VPWR _0278_ _2664_ VGND sg13g2_inv_1
XFILLER_29_434 VPWR VGND sg13g2_fill_2
XFILLER_45_949 VPWR VGND sg13g2_decap_8
X_6699__134 VPWR VGND net134 sg13g2_tiehi
XFILLER_16_139 VPWR VGND sg13g2_decap_8
XFILLER_13_813 VPWR VGND sg13g2_decap_4
XFILLER_13_835 VPWR VGND sg13g2_decap_4
XFILLER_8_305 VPWR VGND sg13g2_fill_2
XFILLER_13_879 VPWR VGND sg13g2_fill_2
XFILLER_0_761 VPWR VGND sg13g2_decap_8
XFILLER_48_732 VPWR VGND sg13g2_decap_8
XFILLER_47_264 VPWR VGND sg13g2_decap_4
XFILLER_47_286 VPWR VGND sg13g2_fill_2
XFILLER_44_960 VPWR VGND sg13g2_decap_8
XFILLER_43_470 VPWR VGND sg13g2_fill_2
X_4600_ net1074 net571 _2098_ VPWR VGND sg13g2_and2_1
X_5580_ net1011 _2777_ _2985_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1018 VPWR VGND sg13g2_decap_8
X_6615__224 VPWR VGND net224 sg13g2_tiehi
X_4531_ s0.data_out\[6\]\[0\] s0.data_out\[5\]\[0\] net1081 _2030_ VPWR VGND sg13g2_mux2_1
Xhold305 s0.data_out\[1\]\[7\] VPWR VGND net625 sg13g2_dlygate4sd3_1
Xhold316 s0.data_out\[10\]\[6\] VPWR VGND net636 sg13g2_dlygate4sd3_1
X_4462_ _1970_ _1972_ net1431 _1973_ VPWR VGND sg13g2_nand3_1
Xhold349 s0.data_out\[6\]\[4\] VPWR VGND net669 sg13g2_dlygate4sd3_1
Xhold338 _0055_ VPWR VGND net658 sg13g2_dlygate4sd3_1
X_3413_ _1027_ net1219 net602 VPWR VGND sg13g2_nand2_1
Xhold327 s0.data_out\[14\]\[1\] VPWR VGND net647 sg13g2_dlygate4sd3_1
X_6201_ _0692_ _0748_ net1471 _0749_ VPWR VGND sg13g2_nand3_1
X_4393_ net1089 _1901_ _1907_ VPWR VGND sg13g2_nor2_1
X_6132_ s0.data_out\[18\]\[1\] s0.data_out\[17\]\[1\] net1259 _0681_ VPWR VGND sg13g2_mux2_1
XFILLER_30_0 VPWR VGND sg13g2_decap_8
X_6063_ _0624_ net436 net1282 VPWR VGND sg13g2_nand2b_1
X_5014_ net1030 _2463_ _2468_ VPWR VGND sg13g2_nor2_1
X_6622__217 VPWR VGND net217 sg13g2_tiehi
XFILLER_42_908 VPWR VGND sg13g2_decap_8
XFILLER_35_960 VPWR VGND sg13g2_decap_8
X_5916_ _0487_ net1273 _0488_ _0489_ VPWR VGND sg13g2_a21o_1
X_5847_ net1305 VPWR _0428_ VGND _0361_ _0427_ sg13g2_o21ai_1
X_5778_ _0363_ s0.data_out\[20\]\[3\] net1309 VPWR VGND sg13g2_nand2b_1
X_4729_ _2142_ _2214_ net1474 _2215_ VPWR VGND sg13g2_nand3_1
XFILLER_1_547 VPWR VGND sg13g2_decap_8
XFILLER_29_253 VPWR VGND sg13g2_fill_1
XFILLER_29_297 VPWR VGND sg13g2_decap_4
XFILLER_45_779 VPWR VGND sg13g2_decap_8
XFILLER_44_278 VPWR VGND sg13g2_fill_2
XFILLER_26_971 VPWR VGND sg13g2_decap_8
XFILLER_32_407 VPWR VGND sg13g2_fill_2
XFILLER_41_952 VPWR VGND sg13g2_decap_8
XFILLER_16_72 VPWR VGND sg13g2_fill_1
XFILLER_12_153 VPWR VGND sg13g2_fill_2
XFILLER_40_473 VPWR VGND sg13g2_decap_8
XFILLER_13_687 VPWR VGND sg13g2_decap_8
XFILLER_13_698 VPWR VGND sg13g2_fill_2
XFILLER_32_60 VPWR VGND sg13g2_fill_1
XFILLER_5_820 VPWR VGND sg13g2_decap_8
XFILLER_32_93 VPWR VGND sg13g2_fill_2
XFILLER_48_562 VPWR VGND sg13g2_decap_8
XFILLER_36_746 VPWR VGND sg13g2_fill_1
X_6750_ net79 VGND VPWR net357 s0.was_valid_out\[2\][0] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_17_971 VPWR VGND sg13g2_decap_8
X_5701_ VGND VPWR _0298_ net1329 net330 sg13g2_or2_1
X_3962_ VGND VPWR _1528_ net1331 net341 sg13g2_or2_1
X_6681_ net153 VGND VPWR _0191_ s0.shift_out\[8\][0] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_3893_ VGND VPWR _1352_ _1458_ _1459_ net1181 sg13g2_a21oi_1
XFILLER_31_451 VPWR VGND sg13g2_fill_1
XFILLER_32_985 VPWR VGND sg13g2_decap_8
X_5632_ net1303 net1170 _3026_ VPWR VGND sg13g2_nor2b_1
X_5563_ net1323 _2967_ _2968_ _2969_ VPWR VGND sg13g2_nor3_1
X_4514_ net1078 _2012_ _2016_ VPWR VGND sg13g2_nor2_1
Xhold113 _0047_ VPWR VGND net433 sg13g2_dlygate4sd3_1
Xhold135 s0.data_out\[23\]\[6\] VPWR VGND net455 sg13g2_dlygate4sd3_1
X_5494_ _2901_ _2902_ _2903_ VPWR VGND sg13g2_nor2_1
Xhold102 s0.data_out\[11\]\[2\] VPWR VGND net422 sg13g2_dlygate4sd3_1
Xhold124 s0.data_out\[4\]\[3\] VPWR VGND net444 sg13g2_dlygate4sd3_1
Xhold168 s0.data_out\[5\]\[7\] VPWR VGND net488 sg13g2_dlygate4sd3_1
X_4445_ _1956_ _1955_ net1402 _1948_ net1411 VPWR VGND sg13g2_a22oi_1
Xhold157 s0.data_out\[10\]\[3\] VPWR VGND net477 sg13g2_dlygate4sd3_1
Xhold146 _0182_ VPWR VGND net466 sg13g2_dlygate4sd3_1
X_4376_ net1375 _1858_ _1893_ VPWR VGND sg13g2_nor2_1
Xhold179 s0.data_out\[18\]\[7\] VPWR VGND net499 sg13g2_dlygate4sd3_1
X_6115_ VGND VPWR _0667_ _0666_ _0664_ sg13g2_or2_1
X_6046_ VGND VPWR net1274 _0604_ _0607_ _0606_ sg13g2_a21oi_1
XFILLER_26_289 VPWR VGND sg13g2_fill_2
X_6696__137 VPWR VGND net137 sg13g2_tiehi
XFILLER_10_635 VPWR VGND sg13g2_fill_1
XFILLER_2_812 VPWR VGND sg13g2_decap_8
XFILLER_49_315 VPWR VGND sg13g2_decap_8
XFILLER_2_889 VPWR VGND sg13g2_decap_8
XFILLER_49_348 VPWR VGND sg13g2_fill_1
XFILLER_18_713 VPWR VGND sg13g2_decap_4
XFILLER_14_985 VPWR VGND sg13g2_decap_8
XFILLER_13_462 VPWR VGND sg13g2_decap_8
X_6612__227 VPWR VGND net227 sg13g2_tiehi
X_4230_ net1000 _2854_ _1764_ VPWR VGND sg13g2_nor2_1
X_4161_ _1696_ net1118 net673 VPWR VGND sg13g2_nand2_1
X_4092_ _1639_ _1630_ _1638_ VPWR VGND sg13g2_nand2_1
X_4994_ net1360 net388 _2452_ VPWR VGND sg13g2_nor2_1
XFILLER_17_1013 VPWR VGND sg13g2_decap_8
XFILLER_23_18 VPWR VGND sg13g2_decap_8
X_3945_ s0.data_out\[11\]\[4\] s0.data_out\[10\]\[4\] net1176 _1511_ VPWR VGND sg13g2_mux2_1
X_6733_ net97 VGND VPWR net445 s0.data_out\[4\]\[3\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_6664_ net172 VGND VPWR _0174_ s0.data_out\[10\]\[6\] clknet_leaf_20_clk sg13g2_dfrbpq_2
XFILLER_20_922 VPWR VGND sg13g2_decap_4
XFILLER_23_29 VPWR VGND sg13g2_fill_2
X_3876_ _1446_ net1338 net1175 VPWR VGND sg13g2_nand2_1
X_5615_ _3010_ VPWR _3012_ VGND s0.was_valid_out\[21\][0] net1307 sg13g2_o21ai_1
XFILLER_20_955 VPWR VGND sg13g2_decap_8
X_6761__67 VPWR VGND net67 sg13g2_tiehi
X_6595_ net246 VGND VPWR _0105_ s0.data_out\[15\]\[4\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_5546_ s0.data_out\[23\]\[6\] s0.data_out\[22\]\[6\] net1318 _2952_ VPWR VGND sg13g2_mux2_1
XFILLER_2_108 VPWR VGND sg13g2_fill_1
X_5477_ VGND VPWR _2768_ net991 net6 _2890_ sg13g2_a21oi_1
X_4428_ VGND VPWR _1824_ _1938_ _1939_ net1097 sg13g2_a21oi_1
X_4359_ net1110 VPWR _1880_ VGND _1810_ _1879_ sg13g2_o21ai_1
XFILLER_47_808 VPWR VGND sg13g2_decap_8
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
X_6029_ VGND VPWR _0477_ _0589_ _0590_ net1278 sg13g2_a21oi_1
XFILLER_27_510 VPWR VGND sg13g2_fill_1
XFILLER_27_532 VPWR VGND sg13g2_decap_8
X_6563__281 VPWR VGND net281 sg13g2_tiehi
XFILLER_14_204 VPWR VGND sg13g2_fill_2
XFILLER_27_576 VPWR VGND sg13g2_fill_1
XFILLER_30_708 VPWR VGND sg13g2_fill_1
XFILLER_7_904 VPWR VGND sg13g2_decap_8
XFILLER_11_955 VPWR VGND sg13g2_decap_8
XFILLER_6_436 VPWR VGND sg13g2_fill_2
XFILLER_10_487 VPWR VGND sg13g2_decap_4
XFILLER_2_620 VPWR VGND sg13g2_decap_8
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_2_686 VPWR VGND sg13g2_decap_8
XFILLER_49_156 VPWR VGND sg13g2_fill_2
XFILLER_49_134 VPWR VGND sg13g2_fill_1
XFILLER_38_819 VPWR VGND sg13g2_fill_2
XFILLER_1_196 VPWR VGND sg13g2_fill_1
XFILLER_37_329 VPWR VGND sg13g2_fill_2
XFILLER_38_81 VPWR VGND sg13g2_decap_8
XFILLER_46_841 VPWR VGND sg13g2_decap_8
XFILLER_14_760 VPWR VGND sg13g2_fill_1
X_3730_ net1196 net414 _1315_ VPWR VGND sg13g2_and2_1
X_3661_ net1192 net994 _1251_ VPWR VGND sg13g2_nor2_1
X_6380_ _0905_ s0.data_out\[15\]\[1\] net1248 VPWR VGND sg13g2_nand2b_1
X_5400_ VPWR _2818_ net530 VGND sg13g2_inv_1
X_3592_ _1192_ VPWR _1193_ VGND net1477 net591 sg13g2_o21ai_1
XFILLER_6_970 VPWR VGND sg13g2_decap_8
X_5331_ _2749_ net1316 VPWR VGND sg13g2_inv_2
X_5262_ VGND VPWR _2689_ _2688_ net1416 sg13g2_or2_1
X_4213_ net1116 net1159 _1748_ VPWR VGND sg13g2_nor2b_1
X_5193_ _2632_ s0.data_out\[1\]\[4\] net1024 VPWR VGND sg13g2_nand2b_1
X_4144_ VGND VPWR _1682_ _1681_ _1679_ sg13g2_or2_1
X_4075_ _1619_ _1620_ _1622_ VPWR VGND _1621_ sg13g2_nand3b_1
X_6547__298 VPWR VGND net298 sg13g2_tiehi
XFILLER_36_362 VPWR VGND sg13g2_fill_2
XFILLER_36_384 VPWR VGND sg13g2_decap_4
X_6716_ net115 VGND VPWR _0226_ s0.genblk1\[4\].modules.bubble clknet_leaf_13_clk
+ sg13g2_dfrbpq_1
X_4977_ _2383_ _2438_ net1473 _2439_ VPWR VGND sg13g2_nand3_1
X_3928_ s0.data_out\[11\]\[6\] s0.data_out\[10\]\[6\] net1176 _1494_ VPWR VGND sg13g2_mux2_1
Xclkload5 clkload5/Y clknet_leaf_28_clk VPWR VGND sg13g2_inv_2
X_6647_ net190 VGND VPWR net351 s0.was_valid_out\[10\][0] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3859_ _1432_ VPWR _1433_ VGND net1015 _1431_ sg13g2_o21ai_1
XFILLER_30_1010 VPWR VGND sg13g2_decap_8
X_6578_ net264 VGND VPWR _0088_ s0.shift_out\[16\][0] clknet_leaf_32_clk sg13g2_dfrbpq_1
XFILLER_4_929 VPWR VGND sg13g2_decap_8
XFILLER_3_417 VPWR VGND sg13g2_fill_1
X_5529_ net1315 net993 _2935_ VPWR VGND sg13g2_nor2_1
X_6498__55 VPWR VGND net55 sg13g2_tiehi
Xfanout1229 net1230 net1229 VPWR VGND sg13g2_buf_8
Xfanout1218 net365 net1218 VPWR VGND sg13g2_buf_8
Xfanout1207 net1208 net1207 VPWR VGND sg13g2_buf_2
XFILLER_46_104 VPWR VGND sg13g2_fill_1
XFILLER_47_649 VPWR VGND sg13g2_decap_4
XFILLER_28_841 VPWR VGND sg13g2_fill_1
XFILLER_43_811 VPWR VGND sg13g2_decap_4
XFILLER_27_384 VPWR VGND sg13g2_fill_1
XFILLER_27_395 VPWR VGND sg13g2_fill_2
XFILLER_24_94 VPWR VGND sg13g2_decap_8
XFILLER_11_796 VPWR VGND sg13g2_fill_1
XFILLER_40_82 VPWR VGND sg13g2_fill_1
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_19_830 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_14 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_18_340 VPWR VGND sg13g2_fill_2
XFILLER_34_811 VPWR VGND sg13g2_decap_4
X_4900_ net1468 net334 _0250_ VPWR VGND sg13g2_and2_1
X_5880_ net1466 net325 _0039_ VPWR VGND sg13g2_and2_1
XFILLER_46_693 VPWR VGND sg13g2_fill_2
XFILLER_46_682 VPWR VGND sg13g2_decap_8
XFILLER_34_822 VPWR VGND sg13g2_fill_1
X_4831_ _2306_ net1063 _2305_ VPWR VGND sg13g2_nand2b_1
XFILLER_34_877 VPWR VGND sg13g2_decap_8
XFILLER_21_527 VPWR VGND sg13g2_decap_8
XFILLER_34_899 VPWR VGND sg13g2_decap_4
X_4762_ _0235_ _2239_ _2240_ _2867_ net1364 VPWR VGND sg13g2_a22oi_1
X_4693_ _2180_ net492 net1082 VPWR VGND sg13g2_nand2b_1
X_6501_ net52 VGND VPWR net456 s0.data_out\[23\]\[6\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_14_1027 VPWR VGND sg13g2_fill_2
X_3713_ net1191 s0.data_out\[12\]\[0\] _1302_ VPWR VGND sg13g2_and2_1
X_6432_ _0957_ net430 net1248 VPWR VGND sg13g2_nand2b_1
X_3644_ _1234_ net1197 net442 VPWR VGND sg13g2_nand2_1
XFILLER_20_19 VPWR VGND sg13g2_fill_2
X_6363_ _0888_ VPWR _0891_ VGND net1241 _0890_ sg13g2_o21ai_1
X_6553__291 VPWR VGND net291 sg13g2_tiehi
X_3575_ _1177_ net1211 s0.data_out\[13\]\[4\] VPWR VGND sg13g2_nand2_1
X_5314_ VPWR _2732_ net358 VGND sg13g2_inv_1
X_6294_ _0831_ _0827_ _0828_ _0829_ VPWR VGND sg13g2_and3_1
X_5245_ VGND VPWR net1022 net394 _2677_ _2620_ sg13g2_a21oi_1
Xhold17 s0.genblk1\[18\].modules.bubble VPWR VGND net337 sg13g2_dlygate4sd3_1
X_6495__58 VPWR VGND net58 sg13g2_tiehi
Xhold28 s0.was_valid_out\[12\][0] VPWR VGND net348 sg13g2_dlygate4sd3_1
XFILLER_29_39 VPWR VGND sg13g2_fill_1
X_5176_ VGND VPWR s0.shift_out\[0\][0] _2613_ _2615_ _2614_ sg13g2_a21oi_1
Xhold39 _0188_ VPWR VGND net359 sg13g2_dlygate4sd3_1
X_4127_ VGND VPWR net1013 _1636_ _1668_ net1387 sg13g2_a21oi_1
X_4058_ _1605_ net1132 s0.data_out\[9\]\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_37_671 VPWR VGND sg13g2_fill_1
X_6560__284 VPWR VGND net284 sg13g2_tiehi
XFILLER_40_858 VPWR VGND sg13g2_decap_4
XFILLER_4_704 VPWR VGND sg13g2_decap_8
Xfanout1004 net1006 net1004 VPWR VGND sg13g2_buf_8
Xfanout1026 s0.valid_out\[0\][0] net1026 VPWR VGND sg13g2_buf_8
XFILLER_0_943 VPWR VGND sg13g2_decap_8
Xfanout1015 net1016 net1015 VPWR VGND sg13g2_buf_8
Xfanout1037 net1042 net1037 VPWR VGND sg13g2_buf_1
XFILLER_48_914 VPWR VGND sg13g2_decap_8
Xfanout1059 s0.valid_out\[3\][0] net1059 VPWR VGND sg13g2_buf_8
Xfanout1048 net1055 net1048 VPWR VGND sg13g2_buf_1
XFILLER_19_137 VPWR VGND sg13g2_decap_8
XFILLER_28_693 VPWR VGND sg13g2_fill_2
XFILLER_43_663 VPWR VGND sg13g2_decap_8
XFILLER_42_162 VPWR VGND sg13g2_fill_2
XFILLER_15_365 VPWR VGND sg13g2_fill_2
XFILLER_16_888 VPWR VGND sg13g2_decap_4
XFILLER_35_93 VPWR VGND sg13g2_fill_1
XFILLER_30_368 VPWR VGND sg13g2_decap_4
XFILLER_7_564 VPWR VGND sg13g2_fill_2
XFILLER_44_1009 VPWR VGND sg13g2_decap_8
X_5030_ net1027 net1170 _2481_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_947 VPWR VGND sg13g2_decap_8
X_5932_ _0505_ net1283 net486 VPWR VGND sg13g2_nand2_1
X_5863_ _0035_ _0439_ _0440_ _2780_ net1344 VPWR VGND sg13g2_a22oi_1
X_4814_ VGND VPWR net1064 _2286_ _2289_ _2288_ sg13g2_a21oi_1
X_5794_ _0379_ net1296 net432 VPWR VGND sg13g2_nand2_1
X_4745_ net1061 s0.data_out\[4\]\[4\] _2227_ VPWR VGND sg13g2_and2_1
X_4676_ net1439 _2162_ _2163_ VPWR VGND sg13g2_nor2_1
X_6415_ VGND VPWR _0940_ _0931_ net1411 sg13g2_or2_1
X_3627_ _1219_ VPWR _1220_ VGND net1208 _1107_ sg13g2_o21ai_1
X_6346_ _0082_ _0875_ _0876_ _2804_ net1365 VPWR VGND sg13g2_a22oi_1
X_3558_ VGND VPWR _1043_ _1159_ _1160_ net1218 sg13g2_a21oi_1
XFILLER_0_228 VPWR VGND sg13g2_decap_8
X_6277_ s0.data_out\[17\]\[7\] s0.data_out\[16\]\[7\] net1245 _0814_ VPWR VGND sg13g2_mux2_1
X_3489_ net1230 VPWR _1097_ VGND _1057_ _1096_ sg13g2_o21ai_1
Xheichips25_top_sorter_319 VPWR VGND uio_oe[2] sg13g2_tiehi
X_5228_ _2663_ VPWR _2664_ VGND net1464 net683 sg13g2_o21ai_1
XFILLER_5_1025 VPWR VGND sg13g2_decap_4
X_5159_ net1020 net1170 _2598_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_446 VPWR VGND sg13g2_fill_1
XFILLER_45_928 VPWR VGND sg13g2_decap_8
XFILLER_29_468 VPWR VGND sg13g2_decap_8
XFILLER_38_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_36_clk clknet_3_1__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_24_140 VPWR VGND sg13g2_decap_8
XFILLER_25_663 VPWR VGND sg13g2_decap_4
XFILLER_40_666 VPWR VGND sg13g2_decap_8
XFILLER_12_368 VPWR VGND sg13g2_fill_1
XFILLER_40_699 VPWR VGND sg13g2_decap_8
XFILLER_21_95 VPWR VGND sg13g2_fill_2
XFILLER_4_578 VPWR VGND sg13g2_fill_2
XFILLER_0_740 VPWR VGND sg13g2_decap_8
XFILLER_48_711 VPWR VGND sg13g2_decap_8
X_6608__232 VPWR VGND net232 sg13g2_tiehi
XFILLER_48_788 VPWR VGND sg13g2_decap_8
XFILLER_29_980 VPWR VGND sg13g2_decap_8
XFILLER_16_641 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_27_clk clknet_3_5__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_16_696 VPWR VGND sg13g2_decap_8
XFILLER_8_840 VPWR VGND sg13g2_fill_1
X_4530_ net1074 net1172 _2029_ VPWR VGND sg13g2_nor2b_1
Xhold317 s0.data_out\[8\]\[3\] VPWR VGND net637 sg13g2_dlygate4sd3_1
X_4461_ _1972_ _1971_ net1097 VPWR VGND sg13g2_nand2b_1
Xhold306 s0.data_out\[10\]\[0\] VPWR VGND net626 sg13g2_dlygate4sd3_1
Xhold339 s0.data_out\[21\]\[5\] VPWR VGND net659 sg13g2_dlygate4sd3_1
Xhold328 s0.data_out\[21\]\[0\] VPWR VGND net648 sg13g2_dlygate4sd3_1
X_3412_ VPWR VGND _1024_ net1460 _1022_ net1454 _1026_ _1018_ sg13g2_a221oi_1
X_6200_ net1267 VPWR _0748_ VGND _0688_ _0747_ sg13g2_o21ai_1
X_4392_ VGND VPWR _1906_ _1905_ _1903_ sg13g2_or2_1
X_6131_ _0680_ net1260 net529 VPWR VGND sg13g2_nand2_1
X_6062_ _0621_ net1264 _0622_ _0623_ VPWR VGND sg13g2_a21o_1
X_5013_ _2465_ VPWR _2467_ VGND s0.was_valid_out\[1\][0] net1034 sg13g2_o21ai_1
XFILLER_38_221 VPWR VGND sg13g2_fill_2
XFILLER_39_755 VPWR VGND sg13g2_fill_2
Xfanout1390 uio_in[1] net1390 VPWR VGND sg13g2_buf_8
XFILLER_38_298 VPWR VGND sg13g2_decap_8
XFILLER_26_427 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_18_clk clknet_3_6__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
X_5915_ net1273 net1143 _0488_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_460 VPWR VGND sg13g2_fill_2
X_5846_ net1290 s0.data_out\[20\]\[3\] _0427_ VPWR VGND sg13g2_and2_1
XFILLER_21_143 VPWR VGND sg13g2_fill_2
XFILLER_22_677 VPWR VGND sg13g2_decap_8
XFILLER_10_839 VPWR VGND sg13g2_fill_2
X_5777_ _0360_ net1290 _0361_ _0362_ VPWR VGND sg13g2_a21o_1
XFILLER_21_198 VPWR VGND sg13g2_decap_8
X_4728_ net1073 VPWR _2214_ VGND _2143_ _2213_ sg13g2_o21ai_1
X_4659_ _2146_ net1072 _2145_ VPWR VGND sg13g2_nand2b_1
XFILLER_1_526 VPWR VGND sg13g2_decap_8
X_6329_ _0078_ _0862_ _0863_ _2807_ net1366 VPWR VGND sg13g2_a22oi_1
XFILLER_29_243 VPWR VGND sg13g2_fill_2
XFILLER_17_427 VPWR VGND sg13g2_fill_1
XFILLER_45_758 VPWR VGND sg13g2_decap_8
XFILLER_44_235 VPWR VGND sg13g2_fill_2
XFILLER_26_950 VPWR VGND sg13g2_decap_8
XFILLER_40_463 VPWR VGND sg13g2_fill_1
XFILLER_13_666 VPWR VGND sg13g2_decap_8
XFILLER_34_1019 VPWR VGND sg13g2_decap_8
XFILLER_8_169 VPWR VGND sg13g2_decap_8
XFILLER_8_147 VPWR VGND sg13g2_fill_2
XFILLER_36_736 VPWR VGND sg13g2_fill_1
XFILLER_35_213 VPWR VGND sg13g2_fill_2
XFILLER_24_909 VPWR VGND sg13g2_fill_2
X_3961_ _1448_ _1525_ _1526_ _1527_ VPWR VGND sg13g2_nor3_1
X_5700_ _0296_ _3092_ _0297_ VPWR VGND sg13g2_nor2b_1
X_6680_ net154 VGND VPWR _0190_ s0.genblk1\[7\].modules.bubble clknet_leaf_18_clk
+ sg13g2_dfrbpq_1
X_3892_ _1458_ s0.data_out\[10\]\[2\] net1190 VPWR VGND sg13g2_nand2b_1
XFILLER_32_964 VPWR VGND sg13g2_decap_8
X_5631_ _3025_ net1011 _3024_ VPWR VGND sg13g2_nand2_1
X_5562_ net1327 s0.data_out\[22\]\[5\] _2968_ VPWR VGND sg13g2_nor2_1
X_4513_ _2013_ VPWR _2015_ VGND net345 net1083 sg13g2_o21ai_1
XFILLER_7_180 VPWR VGND sg13g2_decap_8
X_5493_ VGND VPWR _2739_ _2750_ _2902_ net1324 sg13g2_a21oi_1
Xhold114 s0.data_out\[3\]\[2\] VPWR VGND net434 sg13g2_dlygate4sd3_1
Xhold103 _0151_ VPWR VGND net423 sg13g2_dlygate4sd3_1
Xhold125 _0243_ VPWR VGND net445 sg13g2_dlygate4sd3_1
X_6689__145 VPWR VGND net145 sg13g2_tiehi
X_4444_ VGND VPWR net1100 _1952_ _1955_ _1954_ sg13g2_a21oi_1
Xhold136 _0011_ VPWR VGND net456 sg13g2_dlygate4sd3_1
Xhold147 s0.data_out\[12\]\[3\] VPWR VGND net467 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_3_2__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold158 _0171_ VPWR VGND net478 sg13g2_dlygate4sd3_1
X_4375_ net1114 VPWR _1892_ VGND _1855_ _1891_ sg13g2_o21ai_1
Xhold169 s0.data_out\[10\]\[1\] VPWR VGND net489 sg13g2_dlygate4sd3_1
X_6114_ net383 net1258 _0666_ VPWR VGND sg13g2_nor2_1
X_6045_ VGND VPWR _0493_ _0605_ _0606_ net1274 sg13g2_a21oi_1
XFILLER_39_552 VPWR VGND sg13g2_fill_1
XFILLER_27_758 VPWR VGND sg13g2_fill_1
XFILLER_42_739 VPWR VGND sg13g2_decap_4
XFILLER_41_238 VPWR VGND sg13g2_fill_1
XFILLER_34_290 VPWR VGND sg13g2_decap_8
X_5829_ _0412_ _0413_ _0414_ VPWR VGND sg13g2_nor2_1
XFILLER_5_128 VPWR VGND sg13g2_fill_1
XFILLER_2_868 VPWR VGND sg13g2_decap_8
XFILLER_40_1023 VPWR VGND sg13g2_decap_4
XFILLER_17_202 VPWR VGND sg13g2_decap_8
XFILLER_45_533 VPWR VGND sg13g2_decap_8
X_6605__235 VPWR VGND net235 sg13g2_tiehi
XFILLER_27_50 VPWR VGND sg13g2_fill_1
XFILLER_27_72 VPWR VGND sg13g2_decap_8
XFILLER_27_83 VPWR VGND sg13g2_fill_1
XFILLER_14_964 VPWR VGND sg13g2_decap_8
XFILLER_9_434 VPWR VGND sg13g2_fill_1
X_4160_ net1111 net1168 _1695_ VPWR VGND sg13g2_nor2b_1
X_4091_ _1635_ _1637_ net1424 _1638_ VPWR VGND sg13g2_nand3_1
XFILLER_48_382 VPWR VGND sg13g2_fill_2
XFILLER_36_588 VPWR VGND sg13g2_fill_1
X_4993_ net1048 VPWR _2451_ VGND _2423_ _2450_ sg13g2_o21ai_1
X_6732_ net98 VGND VPWR _0242_ s0.data_out\[4\]\[2\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3944_ VGND VPWR _1507_ _1509_ _1510_ net1424 sg13g2_a21oi_1
X_6663_ net173 VGND VPWR _0173_ s0.data_out\[10\]\[5\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_32_794 VPWR VGND sg13g2_fill_2
X_3875_ net1185 VPWR _1445_ VGND net1395 net1140 sg13g2_o21ai_1
X_5614_ VGND VPWR net1012 _2895_ _3011_ _3010_ sg13g2_a21oi_1
X_6594_ net247 VGND VPWR net554 s0.data_out\[15\]\[3\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_5545_ _2951_ net1319 net593 VPWR VGND sg13g2_nand2_1
X_5476_ s0.data_out\[23\]\[4\] net991 _2890_ VPWR VGND sg13g2_nor2_1
X_4427_ _1938_ _2760_ net389 VPWR VGND sg13g2_nand2_1
X_4358_ net1098 net408 _1879_ VPWR VGND sg13g2_and2_1
X_4289_ _1812_ net408 net1118 VPWR VGND sg13g2_nand2b_1
X_6028_ _0589_ net410 net1284 VPWR VGND sg13g2_nand2b_1
XFILLER_15_728 VPWR VGND sg13g2_fill_2
XFILLER_42_536 VPWR VGND sg13g2_fill_1
XFILLER_42_569 VPWR VGND sg13g2_decap_8
XFILLER_23_750 VPWR VGND sg13g2_fill_2
XFILLER_13_30 VPWR VGND sg13g2_fill_1
XFILLER_10_466 VPWR VGND sg13g2_fill_2
XFILLER_2_665 VPWR VGND sg13g2_decap_8
XFILLER_1_142 VPWR VGND sg13g2_decap_8
XFILLER_38_809 VPWR VGND sg13g2_fill_1
XFILLER_46_820 VPWR VGND sg13g2_decap_8
Xfanout991 net992 net991 VPWR VGND sg13g2_buf_8
X_6679__155 VPWR VGND net155 sg13g2_tiehi
XFILLER_46_897 VPWR VGND sg13g2_decap_8
XFILLER_20_208 VPWR VGND sg13g2_fill_1
XFILLER_9_231 VPWR VGND sg13g2_fill_2
X_3660_ _1249_ VPWR _1250_ VGND net1197 _2827_ sg13g2_o21ai_1
X_3591_ _1191_ VPWR _1192_ VGND net1018 _1190_ sg13g2_o21ai_1
X_5330_ _2748_ net1058 VPWR VGND sg13g2_inv_2
XFILLER_47_1018 VPWR VGND sg13g2_decap_8
X_5261_ _2687_ VPWR _2688_ VGND net1001 net1151 sg13g2_o21ai_1
X_6686__148 VPWR VGND net148 sg13g2_tiehi
X_4212_ s0.data_out\[9\]\[4\] s0.data_out\[8\]\[4\] net1121 _1747_ VPWR VGND sg13g2_mux2_1
X_5192_ _2631_ net1024 s0.data_out\[0\]\[4\] VPWR VGND sg13g2_nand2_1
X_4143_ net358 net1121 _1681_ VPWR VGND sg13g2_nor2_1
X_4074_ net1405 _1611_ _1621_ VPWR VGND sg13g2_nor2_1
XFILLER_37_820 VPWR VGND sg13g2_fill_2
XFILLER_37_864 VPWR VGND sg13g2_decap_8
XFILLER_37_897 VPWR VGND sg13g2_decap_4
XFILLER_34_18 VPWR VGND sg13g2_decap_4
X_6715_ net116 VGND VPWR _0225_ s0.valid_out\[5\][0] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4976_ net1047 VPWR _2438_ VGND _2379_ _2437_ sg13g2_o21ai_1
X_3927_ _1493_ net1175 net636 VPWR VGND sg13g2_nand2_1
XFILLER_32_591 VPWR VGND sg13g2_fill_1
X_6646_ net191 VGND VPWR net452 s0.data_out\[11\]\[7\] clknet_leaf_22_clk sg13g2_dfrbpq_2
Xclkload6 clknet_leaf_29_clk clkload6/Y VPWR VGND sg13g2_inv_4
X_3858_ VGND VPWR net1015 _1397_ _1432_ net1386 sg13g2_a21oi_1
X_6577_ net265 VGND VPWR _0087_ s0.genblk1\[15\].modules.bubble clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_4_908 VPWR VGND sg13g2_decap_8
X_3789_ VGND VPWR net1193 _1365_ _1368_ _1367_ sg13g2_a21oi_1
X_5528_ _2933_ VPWR _2934_ VGND net1320 _2771_ sg13g2_o21ai_1
X_5459_ VPWR _2877_ net574 VGND sg13g2_inv_1
Xfanout1219 net1220 net1219 VPWR VGND sg13g2_buf_8
Xfanout1208 net1209 net1208 VPWR VGND sg13g2_buf_8
X_6602__238 VPWR VGND net238 sg13g2_tiehi
XFILLER_10_241 VPWR VGND sg13g2_fill_2
XFILLER_11_775 VPWR VGND sg13g2_fill_2
XFILLER_10_263 VPWR VGND sg13g2_fill_2
XFILLER_6_267 VPWR VGND sg13g2_fill_1
XFILLER_3_985 VPWR VGND sg13g2_decap_8
XFILLER_49_70 VPWR VGND sg13g2_decap_4
XFILLER_38_606 VPWR VGND sg13g2_decap_4
XFILLER_18_330 VPWR VGND sg13g2_fill_1
Xheichips25_top_sorter_15 VPWR VGND uio_oe[7] sg13g2_tielo
XFILLER_45_171 VPWR VGND sg13g2_fill_2
XFILLER_33_355 VPWR VGND sg13g2_fill_2
X_4830_ VGND VPWR net1050 _2304_ _2305_ _2302_ sg13g2_a21oi_1
X_6692__141 VPWR VGND net141 sg13g2_tiehi
X_4761_ net1363 _2181_ _2240_ VPWR VGND sg13g2_nor2_1
X_4692_ _2177_ net1066 _2178_ _2179_ VPWR VGND sg13g2_a21o_1
X_6500_ net53 VGND VPWR net460 s0.data_out\[23\]\[5\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_14_1006 VPWR VGND sg13g2_decap_8
X_3712_ VGND VPWR _1296_ _1300_ _0124_ _1301_ sg13g2_a21oi_1
X_6431_ _0954_ net1224 _0955_ _0956_ VPWR VGND sg13g2_a21o_1
X_3643_ VGND VPWR _1233_ _1232_ net1445 sg13g2_or2_1
X_6362_ net362 net1247 _0890_ VPWR VGND sg13g2_nor2_1
X_5313_ VPWR _2731_ net364 VGND sg13g2_inv_1
X_3574_ net1204 net1159 _1176_ VPWR VGND sg13g2_nor2b_1
X_6293_ VPWR _0830_ _0829_ VGND sg13g2_inv_1
X_5244_ VPWR _0281_ _2676_ VGND sg13g2_inv_1
X_5175_ net1022 net1142 _2614_ VPWR VGND sg13g2_nor2b_1
Xhold18 s0.genblk1\[20\].modules.bubble VPWR VGND net338 sg13g2_dlygate4sd3_1
Xhold29 _0133_ VPWR VGND net349 sg13g2_dlygate4sd3_1
X_4126_ VGND VPWR net1128 s0.data_out\[9\]\[5\] _1667_ _1633_ sg13g2_a21oi_1
XFILLER_44_609 VPWR VGND sg13g2_fill_2
X_4057_ _1601_ _1603_ _1604_ VPWR VGND sg13g2_nor2_1
XFILLER_43_108 VPWR VGND sg13g2_decap_8
XFILLER_36_193 VPWR VGND sg13g2_fill_2
XFILLER_24_366 VPWR VGND sg13g2_fill_2
X_4959_ s0.data_out\[3\]\[4\] s0.data_out\[2\]\[4\] net1044 _2422_ VPWR VGND sg13g2_mux2_1
XFILLER_20_572 VPWR VGND sg13g2_fill_1
X_6629_ net209 VGND VPWR _0139_ s0.data_out\[12\]\[3\] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_10_20 VPWR VGND sg13g2_fill_2
XFILLER_3_226 VPWR VGND sg13g2_decap_8
XFILLER_3_248 VPWR VGND sg13g2_fill_1
XFILLER_0_922 VPWR VGND sg13g2_decap_8
Xfanout1016 _2744_ net1016 VPWR VGND sg13g2_buf_8
Xfanout1027 net1029 net1027 VPWR VGND sg13g2_buf_8
Xfanout1038 net1042 net1038 VPWR VGND sg13g2_buf_8
Xfanout1005 net1006 net1005 VPWR VGND sg13g2_buf_2
XFILLER_0_999 VPWR VGND sg13g2_decap_8
Xfanout1049 net1050 net1049 VPWR VGND sg13g2_buf_2
XFILLER_19_84 VPWR VGND sg13g2_fill_1
XFILLER_28_672 VPWR VGND sg13g2_decap_8
XFILLER_35_61 VPWR VGND sg13g2_fill_2
XFILLER_43_686 VPWR VGND sg13g2_fill_1
XFILLER_42_141 VPWR VGND sg13g2_fill_1
XFILLER_43_697 VPWR VGND sg13g2_fill_1
XFILLER_42_174 VPWR VGND sg13g2_decap_4
XFILLER_30_314 VPWR VGND sg13g2_decap_8
XFILLER_30_336 VPWR VGND sg13g2_fill_1
XFILLER_7_532 VPWR VGND sg13g2_fill_1
XFILLER_3_782 VPWR VGND sg13g2_decap_8
XFILLER_2_292 VPWR VGND sg13g2_fill_2
XFILLER_39_926 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_4
XFILLER_19_650 VPWR VGND sg13g2_decap_8
X_5931_ _0501_ _0503_ _0504_ VPWR VGND sg13g2_nor2_1
X_5862_ net1344 _0384_ _0440_ VPWR VGND sg13g2_nor2_1
X_4813_ VGND VPWR _2176_ _2287_ _2288_ net1064 sg13g2_a21oi_1
X_5793_ VGND VPWR net1301 _0375_ _0378_ _0377_ sg13g2_a21oi_1
X_4744_ _0231_ _2225_ _2226_ _2866_ net1363 VPWR VGND sg13g2_a22oi_1
X_4675_ VGND VPWR net1073 _2159_ _2162_ _2161_ sg13g2_a21oi_1
X_6414_ _0939_ _0938_ net1402 _0931_ net1411 VPWR VGND sg13g2_a22oi_1
X_3626_ _1219_ _1218_ _1217_ VPWR VGND sg13g2_nand2b_1
X_6345_ net1365 _0838_ _0876_ VPWR VGND sg13g2_nor2_1
X_3557_ _1159_ s0.data_out\[13\]\[6\] net1222 VPWR VGND sg13g2_nand2b_1
X_6276_ _0813_ net1247 net503 VPWR VGND sg13g2_nand2_1
X_3488_ net1215 s0.data_out\[14\]\[5\] _1096_ VPWR VGND sg13g2_and2_1
X_5227_ _2662_ VPWR _2663_ VGND net1004 _2661_ sg13g2_o21ai_1
XFILLER_5_1004 VPWR VGND sg13g2_decap_8
X_5158_ s0.data_out\[1\]\[0\] s0.data_out\[0\]\[0\] net1026 _2597_ VPWR VGND sg13g2_mux2_1
XFILLER_29_436 VPWR VGND sg13g2_fill_1
XFILLER_45_907 VPWR VGND sg13g2_decap_8
X_5089_ _2505_ _2521_ _2536_ _2539_ _2540_ VPWR VGND sg13g2_or4_1
X_4109_ net1135 VPWR _1654_ VGND _1570_ _1653_ sg13g2_o21ai_1
XFILLER_38_970 VPWR VGND sg13g2_decap_8
XFILLER_25_631 VPWR VGND sg13g2_fill_2
XFILLER_13_859 VPWR VGND sg13g2_decap_8
XFILLER_40_689 VPWR VGND sg13g2_fill_1
XFILLER_21_892 VPWR VGND sg13g2_fill_2
XFILLER_47_222 VPWR VGND sg13g2_decap_4
XFILLER_0_796 VPWR VGND sg13g2_decap_8
XFILLER_48_767 VPWR VGND sg13g2_decap_8
XFILLER_28_480 VPWR VGND sg13g2_fill_2
XFILLER_44_995 VPWR VGND sg13g2_decap_8
XFILLER_30_122 VPWR VGND sg13g2_fill_2
XFILLER_31_667 VPWR VGND sg13g2_fill_2
XFILLER_8_852 VPWR VGND sg13g2_decap_4
XFILLER_7_351 VPWR VGND sg13g2_decap_8
Xhold307 s0.data_out\[7\]\[6\] VPWR VGND net627 sg13g2_dlygate4sd3_1
X_4460_ s0.data_out\[6\]\[4\] s0.data_out\[7\]\[4\] net1105 _1971_ VPWR VGND sg13g2_mux2_1
X_4391_ net364 net1094 _1905_ VPWR VGND sg13g2_nor2_1
Xhold329 s0.was_valid_out\[20\][0] VPWR VGND net649 sg13g2_dlygate4sd3_1
X_3411_ _1011_ VPWR _1025_ VGND net1454 _1018_ sg13g2_o21ai_1
Xhold318 _0195_ VPWR VGND net638 sg13g2_dlygate4sd3_1
X_6130_ net1447 _0678_ _0679_ VPWR VGND sg13g2_nor2_1
X_6550__295 VPWR VGND net295 sg13g2_tiehi
X_6061_ net1264 net1152 _0622_ VPWR VGND sg13g2_nor2b_1
X_5012_ VGND VPWR net1010 _2355_ _2466_ _2465_ sg13g2_a21oi_1
XFILLER_38_233 VPWR VGND sg13g2_fill_2
Xfanout1380 net1383 net1380 VPWR VGND sg13g2_buf_8
XFILLER_16_0 VPWR VGND sg13g2_fill_2
Xfanout1391 uio_in[1] net1391 VPWR VGND sg13g2_buf_1
XFILLER_39_789 VPWR VGND sg13g2_fill_2
X_5914_ s0.data_out\[20\]\[7\] s0.data_out\[19\]\[7\] net1281 _0487_ VPWR VGND sg13g2_mux2_1
XFILLER_35_995 VPWR VGND sg13g2_decap_8
X_5845_ VPWR _0031_ _0426_ VGND sg13g2_inv_1
X_5776_ net1290 net1161 _0361_ VPWR VGND sg13g2_nor2b_1
X_4727_ net1061 s0.data_out\[4\]\[0\] _2213_ VPWR VGND sg13g2_and2_1
X_4658_ VGND VPWR net1061 _2144_ _2145_ _2143_ sg13g2_a21oi_1
X_3609_ _1205_ VPWR _1206_ VGND net1484 net522 sg13g2_o21ai_1
X_4589_ _2088_ _2080_ _2087_ VPWR VGND sg13g2_nand2_1
X_6328_ net1366 _0794_ _0863_ VPWR VGND sg13g2_nor2_1
XFILLER_27_1027 VPWR VGND sg13g2_fill_2
X_6259_ s0.data_out\[17\]\[0\] s0.data_out\[16\]\[0\] net1245 _0796_ VPWR VGND sg13g2_mux2_1
XFILLER_44_214 VPWR VGND sg13g2_fill_2
XFILLER_32_409 VPWR VGND sg13g2_fill_1
XFILLER_41_987 VPWR VGND sg13g2_decap_8
XFILLER_5_899 VPWR VGND sg13g2_decap_8
XFILLER_0_593 VPWR VGND sg13g2_decap_8
XFILLER_48_597 VPWR VGND sg13g2_decap_8
X_3960_ _1500_ _1502_ _1526_ VPWR VGND sg13g2_nor2b_1
XFILLER_44_770 VPWR VGND sg13g2_fill_2
XFILLER_43_291 VPWR VGND sg13g2_fill_2
X_3891_ _1455_ net1136 _1456_ _1457_ VPWR VGND sg13g2_a21o_1
XFILLER_31_442 VPWR VGND sg13g2_decap_8
X_5630_ _2923_ VPWR _3024_ VGND net1321 _2783_ sg13g2_o21ai_1
X_5561_ net459 net1327 _2967_ VPWR VGND sg13g2_nor2b_1
X_4512_ VGND VPWR net998 _1902_ _2014_ _2013_ sg13g2_a21oi_1
X_5492_ net1312 _2894_ _2901_ VPWR VGND sg13g2_nor2_1
Xhold126 s0.shift_out\[6\][0] VPWR VGND net446 sg13g2_dlygate4sd3_1
Xhold104 s0.data_out\[20\]\[2\] VPWR VGND net424 sg13g2_dlygate4sd3_1
Xhold115 _0254_ VPWR VGND net435 sg13g2_dlygate4sd3_1
X_4443_ VGND VPWR _1840_ _1953_ _1954_ net1100 sg13g2_a21oi_1
Xhold148 s0.data_out\[20\]\[5\] VPWR VGND net468 sg13g2_dlygate4sd3_1
Xhold159 s0.data_out\[16\]\[1\] VPWR VGND net479 sg13g2_dlygate4sd3_1
Xhold137 s0.data_out\[13\]\[2\] VPWR VGND net457 sg13g2_dlygate4sd3_1
X_4374_ net1102 net470 _1891_ VPWR VGND sg13g2_and2_1
X_6113_ _0664_ VPWR _0665_ VGND net1262 _0554_ sg13g2_o21ai_1
X_6044_ _0605_ net534 net1281 VPWR VGND sg13g2_nand2b_1
XFILLER_41_217 VPWR VGND sg13g2_fill_2
XFILLER_35_770 VPWR VGND sg13g2_decap_4
X_5828_ _0330_ VPWR _0413_ VGND _0386_ _0388_ sg13g2_o21ai_1
XFILLER_23_987 VPWR VGND sg13g2_decap_8
X_5759_ _0344_ net1007 _0343_ VPWR VGND sg13g2_nand2_1
XFILLER_2_847 VPWR VGND sg13g2_decap_8
XFILLER_40_1002 VPWR VGND sg13g2_decap_8
XFILLER_45_567 VPWR VGND sg13g2_decap_8
XFILLER_14_921 VPWR VGND sg13g2_fill_1
XFILLER_43_83 VPWR VGND sg13g2_fill_2
XFILLER_40_250 VPWR VGND sg13g2_fill_1
XFILLER_9_457 VPWR VGND sg13g2_decap_8
XFILLER_4_140 VPWR VGND sg13g2_fill_2
XFILLER_4_22 VPWR VGND sg13g2_fill_1
X_4090_ _1637_ net1013 _1636_ VPWR VGND sg13g2_nand2_1
XFILLER_1_891 VPWR VGND sg13g2_decap_8
XFILLER_49_884 VPWR VGND sg13g2_decap_8
XFILLER_36_523 VPWR VGND sg13g2_fill_1
XFILLER_36_567 VPWR VGND sg13g2_decap_4
XFILLER_24_729 VPWR VGND sg13g2_fill_2
X_4992_ net1037 net583 _2450_ VPWR VGND sg13g2_and2_1
XFILLER_16_291 VPWR VGND sg13g2_fill_2
X_6731_ net99 VGND VPWR _0241_ s0.data_out\[4\]\[1\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_32_751 VPWR VGND sg13g2_decap_4
X_3943_ _1509_ _1508_ net1184 VPWR VGND sg13g2_nand2b_1
X_6662_ net174 VGND VPWR _0172_ s0.data_out\[10\]\[4\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_3874_ _0143_ _1443_ _1444_ _2830_ net1382 VPWR VGND sg13g2_a22oi_1
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
X_5613_ VGND VPWR net1336 net1307 _3010_ _3009_ sg13g2_a21oi_1
XFILLER_31_272 VPWR VGND sg13g2_decap_4
X_6593_ net248 VGND VPWR net421 s0.data_out\[15\]\[2\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_5544_ net1323 _2948_ _2949_ _2950_ VPWR VGND sg13g2_nor3_1
X_5475_ _2889_ VPWR net5 VGND _2771_ net992 sg13g2_o21ai_1
X_4426_ _1935_ net1087 _1936_ _1937_ VPWR VGND sg13g2_a21o_1
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_4357_ VPWR _0192_ net538 VGND sg13g2_inv_1
XFILLER_24_1019 VPWR VGND sg13g2_decap_8
X_4288_ _1809_ net1098 _1810_ _1811_ VPWR VGND sg13g2_a21o_1
X_6027_ _0586_ net1265 _0587_ _0588_ VPWR VGND sg13g2_a21o_1
XFILLER_42_526 VPWR VGND sg13g2_fill_1
XFILLER_14_228 VPWR VGND sg13g2_decap_4
XFILLER_7_939 VPWR VGND sg13g2_decap_8
XFILLER_6_449 VPWR VGND sg13g2_fill_1
XFILLER_2_644 VPWR VGND sg13g2_decap_8
XFILLER_38_50 VPWR VGND sg13g2_decap_8
Xfanout992 _2885_ net992 VPWR VGND sg13g2_buf_8
XFILLER_46_876 VPWR VGND sg13g2_decap_8
XFILLER_45_364 VPWR VGND sg13g2_fill_2
XFILLER_33_537 VPWR VGND sg13g2_fill_1
XFILLER_9_210 VPWR VGND sg13g2_decap_4
X_3590_ VGND VPWR net1018 _1135_ _1191_ net1378 sg13g2_a21oi_1
X_5260_ net395 net1025 net1023 _2687_ VPWR VGND sg13g2_a21o_1
X_4211_ _1746_ net1120 net670 VPWR VGND sg13g2_nand2_1
X_5191_ _2630_ net1005 _2629_ VPWR VGND sg13g2_nand2_1
X_4142_ _1679_ VPWR _1680_ VGND net1126 _1557_ sg13g2_o21ai_1
X_4073_ VGND VPWR _1620_ _1618_ net1414 sg13g2_or2_1
XFILLER_49_681 VPWR VGND sg13g2_decap_8
XFILLER_48_180 VPWR VGND sg13g2_decap_8
XFILLER_48_191 VPWR VGND sg13g2_fill_1
X_4975_ net1036 s0.data_out\[2\]\[0\] _2437_ VPWR VGND sg13g2_and2_1
X_6714_ net118 VGND VPWR net346 s0.was_valid_out\[5\][0] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3926_ VGND VPWR net1184 _1489_ _1492_ _1491_ sg13g2_a21oi_1
XFILLER_20_743 VPWR VGND sg13g2_fill_1
X_6645_ net192 VGND VPWR _0155_ s0.data_out\[11\]\[6\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_3857_ VGND VPWR net1183 net373 _1431_ _1392_ sg13g2_a21oi_1
Xclkload7 VPWR clkload7/Y clknet_leaf_16_clk VGND sg13g2_inv_1
X_6576_ net266 VGND VPWR _0086_ s0.valid_out\[16\][0] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_3788_ VGND VPWR _1249_ _1366_ _1367_ net1193 sg13g2_a21oi_1
X_5527_ _2933_ net1320 net586 VPWR VGND sg13g2_nand2_1
X_5458_ VPWR _2876_ net387 VGND sg13g2_inv_1
XFILLER_8_1024 VPWR VGND sg13g2_decap_4
Xfanout1209 s0.shift_out\[13\][0] net1209 VPWR VGND sg13g2_buf_8
X_5389_ _2807_ net529 VPWR VGND sg13g2_inv_2
X_4409_ net1085 net1169 _1920_ VPWR VGND sg13g2_nor2b_1
XFILLER_28_832 VPWR VGND sg13g2_decap_8
XFILLER_15_515 VPWR VGND sg13g2_fill_2
XFILLER_30_529 VPWR VGND sg13g2_fill_1
XFILLER_10_286 VPWR VGND sg13g2_fill_1
XFILLER_40_51 VPWR VGND sg13g2_fill_2
XFILLER_3_964 VPWR VGND sg13g2_decap_8
XFILLER_2_441 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_16 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_18_342 VPWR VGND sg13g2_fill_1
XFILLER_45_183 VPWR VGND sg13g2_fill_2
X_4760_ net1076 VPWR _2239_ VGND _2178_ _2238_ sg13g2_o21ai_1
X_4691_ net1065 net1143 _2178_ VPWR VGND sg13g2_nor2b_1
X_3711_ VGND VPWR _1301_ net1332 net343 sg13g2_or2_1
X_6430_ net1224 net1154 _0955_ VPWR VGND sg13g2_nor2b_1
X_3642_ VGND VPWR net1204 _1229_ _1232_ _1231_ sg13g2_a21oi_1
X_6361_ net1223 _0884_ _0889_ VPWR VGND sg13g2_nor2_1
X_5312_ VPWR _2730_ net345 VGND sg13g2_inv_1
X_3573_ VGND VPWR _1170_ _1172_ _1175_ net1423 sg13g2_a21oi_1
XFILLER_46_0 VPWR VGND sg13g2_fill_2
X_6292_ VGND VPWR _0829_ _0819_ net1402 sg13g2_or2_1
X_5243_ _2675_ VPWR _2676_ VGND net1467 net579 sg13g2_o21ai_1
Xhold19 s0.genblk1\[6\].modules.bubble VPWR VGND net339 sg13g2_dlygate4sd3_1
X_5174_ s0.data_out\[1\]\[7\] s0.data_out\[0\]\[7\] net1025 _2613_ VPWR VGND sg13g2_mux2_1
X_4125_ VPWR _0172_ _1666_ VGND sg13g2_inv_1
X_4056_ _1602_ VPWR _1603_ VGND _1590_ _1599_ sg13g2_o21ai_1
X_4958_ net1419 _2418_ _2421_ VPWR VGND sg13g2_nor2_1
X_4889_ _2355_ net1336 net1046 VPWR VGND sg13g2_nand2_1
X_3909_ VPWR VGND _1474_ net1459 _1472_ net1454 _1475_ _1468_ sg13g2_a221oi_1
X_6628_ net210 VGND VPWR _0138_ s0.data_out\[12\]\[2\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_4_739 VPWR VGND sg13g2_decap_8
X_6559_ net285 VGND VPWR net441 s0.data_out\[18\]\[4\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_6669__166 VPWR VGND net166 sg13g2_tiehi
XFILLER_0_901 VPWR VGND sg13g2_decap_8
Xfanout1006 _2754_ net1006 VPWR VGND sg13g2_buf_8
Xfanout1017 _2741_ net1017 VPWR VGND sg13g2_buf_8
Xfanout1028 net1029 net1028 VPWR VGND sg13g2_buf_1
Xfanout1039 net1041 net1039 VPWR VGND sg13g2_buf_8
XFILLER_0_978 VPWR VGND sg13g2_decap_8
XFILLER_48_949 VPWR VGND sg13g2_decap_8
XFILLER_16_868 VPWR VGND sg13g2_fill_2
XFILLER_15_367 VPWR VGND sg13g2_fill_1
XFILLER_35_84 VPWR VGND sg13g2_decap_8
X_6676__159 VPWR VGND net159 sg13g2_tiehi
XFILLER_3_761 VPWR VGND sg13g2_decap_8
XFILLER_19_640 VPWR VGND sg13g2_decap_4
XFILLER_20_1011 VPWR VGND sg13g2_decap_8
X_5930_ _0502_ VPWR _0503_ VGND net1409 _0499_ sg13g2_o21ai_1
X_5861_ net1301 VPWR _0439_ VGND _0381_ _0438_ sg13g2_o21ai_1
X_4812_ _2287_ net484 net1069 VPWR VGND sg13g2_nand2b_1
X_5792_ VGND VPWR _3052_ _0376_ _0377_ net1301 sg13g2_a21oi_1
X_4743_ net1363 _2161_ _2226_ VPWR VGND sg13g2_nor2_1
X_6413_ VGND VPWR net1241 _0935_ _0938_ _0937_ sg13g2_a21oi_1
X_4674_ VGND VPWR _2035_ _2160_ _2161_ net1073 sg13g2_a21oi_1
X_3625_ _1218_ net1337 net1198 VPWR VGND sg13g2_nand2_1
X_6344_ net1251 VPWR _0875_ VGND _0835_ _0874_ sg13g2_o21ai_1
XFILLER_1_709 VPWR VGND sg13g2_decap_8
X_3556_ _1156_ net1206 _1157_ _1158_ VPWR VGND sg13g2_a21o_1
X_6275_ _0811_ VPWR _0812_ VGND _0802_ _0803_ sg13g2_o21ai_1
X_3487_ VPWR _0105_ _1095_ VGND sg13g2_inv_1
X_5226_ VGND VPWR net1004 _2583_ _2662_ net1346 sg13g2_a21oi_1
X_5157_ _2596_ net1004 _2595_ VPWR VGND sg13g2_nand2_1
X_5088_ VGND VPWR _2539_ _2538_ _2537_ sg13g2_or2_1
X_6491__63 VPWR VGND net63 sg13g2_tiehi
X_4108_ net1124 s0.data_out\[9\]\[1\] _1653_ VPWR VGND sg13g2_and2_1
X_4039_ VGND VPWR net1124 _1584_ _1586_ _1585_ sg13g2_a21oi_1
XFILLER_48_746 VPWR VGND sg13g2_decap_8
XFILLER_0_775 VPWR VGND sg13g2_decap_8
X_6682__152 VPWR VGND net152 sg13g2_tiehi
XFILLER_44_974 VPWR VGND sg13g2_decap_8
XFILLER_31_613 VPWR VGND sg13g2_decap_4
XFILLER_8_831 VPWR VGND sg13g2_fill_1
XFILLER_31_679 VPWR VGND sg13g2_decap_4
Xhold308 s0.data_out\[20\]\[3\] VPWR VGND net628 sg13g2_dlygate4sd3_1
X_4390_ _1903_ VPWR _1904_ VGND net1101 _1792_ sg13g2_o21ai_1
Xhold319 s0.data_out\[7\]\[4\] VPWR VGND net639 sg13g2_dlygate4sd3_1
X_3410_ _1024_ _1023_ net1228 VPWR VGND sg13g2_nand2b_1
X_6060_ s0.data_out\[19\]\[5\] s0.data_out\[18\]\[5\] net1269 _0621_ VPWR VGND sg13g2_mux2_1
X_5011_ _2463_ _2464_ _2465_ VPWR VGND sg13g2_nor2_1
XFILLER_39_735 VPWR VGND sg13g2_fill_2
XFILLER_38_201 VPWR VGND sg13g2_fill_2
Xfanout1381 net1383 net1381 VPWR VGND sg13g2_buf_8
Xfanout1392 net1393 net1392 VPWR VGND sg13g2_buf_8
Xfanout1370 net1373 net1370 VPWR VGND sg13g2_buf_8
XFILLER_26_429 VPWR VGND sg13g2_fill_1
XFILLER_35_974 VPWR VGND sg13g2_decap_8
X_5913_ _0486_ net1282 net506 VPWR VGND sg13g2_nand2_1
X_5844_ _0425_ VPWR _0426_ VGND net1462 net624 sg13g2_o21ai_1
XFILLER_21_145 VPWR VGND sg13g2_fill_1
XFILLER_10_819 VPWR VGND sg13g2_decap_4
X_5775_ s0.data_out\[21\]\[3\] s0.data_out\[20\]\[3\] net1297 _0360_ VPWR VGND sg13g2_mux2_1
X_4726_ VGND VPWR _2207_ _2211_ _0227_ _2212_ sg13g2_a21oi_1
X_4657_ s0.data_out\[5\]\[0\] s0.data_out\[4\]\[0\] net1068 _2144_ VPWR VGND sg13g2_mux2_1
X_3608_ _1204_ VPWR _1205_ VGND net1017 _1203_ sg13g2_o21ai_1
X_4588_ _2084_ _2086_ net1422 _2087_ VPWR VGND sg13g2_nand3_1
X_6327_ net1255 VPWR _0862_ VGND _0789_ _0861_ sg13g2_o21ai_1
X_3539_ net1203 net994 _1141_ VPWR VGND sg13g2_nor2_1
XFILLER_27_1006 VPWR VGND sg13g2_decap_8
X_6258_ VGND VPWR net1254 _0792_ _0795_ _0794_ sg13g2_a21oi_1
X_5209_ _2644_ _2647_ _2643_ _2648_ VPWR VGND sg13g2_nand3_1
X_6189_ net1421 _0735_ _0738_ VPWR VGND sg13g2_nor2_1
XFILLER_25_451 VPWR VGND sg13g2_fill_1
XFILLER_26_985 VPWR VGND sg13g2_decap_8
XFILLER_41_966 VPWR VGND sg13g2_decap_8
XFILLER_40_432 VPWR VGND sg13g2_fill_1
XFILLER_8_149 VPWR VGND sg13g2_fill_1
XFILLER_4_300 VPWR VGND sg13g2_fill_2
XFILLER_5_834 VPWR VGND sg13g2_decap_8
XFILLER_4_333 VPWR VGND sg13g2_decap_4
XFILLER_5_878 VPWR VGND sg13g2_decap_8
XFILLER_0_572 VPWR VGND sg13g2_decap_8
XFILLER_48_532 VPWR VGND sg13g2_fill_2
XFILLER_48_576 VPWR VGND sg13g2_decap_8
XFILLER_16_451 VPWR VGND sg13g2_decap_8
XFILLER_32_900 VPWR VGND sg13g2_fill_2
XFILLER_17_985 VPWR VGND sg13g2_decap_8
XFILLER_32_933 VPWR VGND sg13g2_fill_2
X_3890_ net1136 net1164 _1456_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_999 VPWR VGND sg13g2_decap_8
X_5560_ VGND VPWR net1324 _2965_ _2966_ _2962_ sg13g2_a21oi_1
X_4511_ VGND VPWR net1337 net1082 _2013_ _2012_ sg13g2_a21oi_1
X_5491_ VGND VPWR _2900_ _2899_ _2896_ sg13g2_or2_1
X_4442_ _1953_ net404 net1107 VPWR VGND sg13g2_nand2b_1
Xhold116 s0.data_out\[18\]\[5\] VPWR VGND net436 sg13g2_dlygate4sd3_1
Xhold105 _0043_ VPWR VGND net425 sg13g2_dlygate4sd3_1
Xhold149 _0046_ VPWR VGND net469 sg13g2_dlygate4sd3_1
Xhold138 _0127_ VPWR VGND net458 sg13g2_dlygate4sd3_1
Xhold127 _2109_ VPWR VGND net447 sg13g2_dlygate4sd3_1
X_4373_ _0196_ _1889_ _1890_ _2850_ net1375 VPWR VGND sg13g2_a22oi_1
X_6112_ _0664_ _0663_ _0662_ VPWR VGND sg13g2_nand2b_1
X_6043_ _0602_ net1261 _0603_ _0604_ VPWR VGND sg13g2_a21o_1
XFILLER_39_543 VPWR VGND sg13g2_fill_1
XFILLER_2_1008 VPWR VGND sg13g2_decap_8
XFILLER_22_443 VPWR VGND sg13g2_decap_8
XFILLER_23_966 VPWR VGND sg13g2_decap_8
X_5827_ _0389_ _0411_ _0412_ VPWR VGND sg13g2_nor2b_1
X_5758_ s0.data_out\[20\]\[0\] s0.data_out\[21\]\[0\] net1309 _0343_ VPWR VGND sg13g2_mux2_1
XFILLER_33_1021 VPWR VGND sg13g2_decap_8
X_4709_ s0.data_out\[5\]\[5\] s0.data_out\[4\]\[5\] net1070 _2196_ VPWR VGND sg13g2_mux2_1
X_5689_ s0.data_out\[21\]\[5\] s0.data_out\[22\]\[5\] net1319 _3083_ VPWR VGND sg13g2_mux2_1
XFILLER_2_826 VPWR VGND sg13g2_decap_8
XFILLER_1_303 VPWR VGND sg13g2_fill_2
XFILLER_49_329 VPWR VGND sg13g2_decap_8
XFILLER_13_432 VPWR VGND sg13g2_fill_1
XFILLER_25_281 VPWR VGND sg13g2_fill_1
XFILLER_13_476 VPWR VGND sg13g2_decap_8
XFILLER_14_999 VPWR VGND sg13g2_decap_8
XFILLER_41_796 VPWR VGND sg13g2_decap_4
XFILLER_13_487 VPWR VGND sg13g2_fill_1
X_6507__45 VPWR VGND net45 sg13g2_tiehi
XFILLER_5_620 VPWR VGND sg13g2_decap_8
XFILLER_5_675 VPWR VGND sg13g2_fill_1
XFILLER_1_870 VPWR VGND sg13g2_decap_8
XFILLER_0_380 VPWR VGND sg13g2_decap_4
XFILLER_49_863 VPWR VGND sg13g2_decap_8
X_6730_ net100 VGND VPWR _0240_ s0.data_out\[4\]\[0\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_4991_ _0255_ _2448_ _2449_ _2877_ net1348 VPWR VGND sg13g2_a22oi_1
XFILLER_32_741 VPWR VGND sg13g2_decap_4
X_3942_ s0.data_out\[10\]\[5\] s0.data_out\[11\]\[5\] net1189 _1508_ VPWR VGND sg13g2_mux2_1
XFILLER_17_1027 VPWR VGND sg13g2_fill_2
X_3873_ net1382 _1379_ _1444_ VPWR VGND sg13g2_nor2_1
X_6661_ net175 VGND VPWR net478 s0.data_out\[10\]\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_5612_ net1313 VPWR _3009_ VGND net1392 net1300 sg13g2_o21ai_1
X_6592_ net249 VGND VPWR net531 s0.data_out\[15\]\[1\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_32_796 VPWR VGND sg13g2_fill_1
X_5543_ net1327 s0.data_out\[22\]\[6\] _2949_ VPWR VGND sg13g2_nor2_1
XFILLER_20_969 VPWR VGND sg13g2_decap_8
X_5474_ _2889_ net1435 net991 VPWR VGND sg13g2_nand2_1
X_4425_ net1087 net994 _1936_ VPWR VGND sg13g2_nor2_1
X_4356_ _1877_ VPWR _1878_ VGND net1481 net537 sg13g2_o21ai_1
X_4287_ net1098 net1168 _1810_ VPWR VGND sg13g2_nor2b_1
X_6026_ net1265 net993 _0587_ VPWR VGND sg13g2_nor2_1
XFILLER_39_384 VPWR VGND sg13g2_decap_8
XFILLER_27_546 VPWR VGND sg13g2_fill_1
XFILLER_42_516 VPWR VGND sg13g2_fill_1
XFILLER_10_402 VPWR VGND sg13g2_fill_2
XFILLER_11_925 VPWR VGND sg13g2_decap_8
XFILLER_23_752 VPWR VGND sg13g2_fill_1
XFILLER_11_936 VPWR VGND sg13g2_fill_2
XFILLER_7_918 VPWR VGND sg13g2_decap_8
XFILLER_10_468 VPWR VGND sg13g2_fill_1
XFILLER_11_969 VPWR VGND sg13g2_decap_8
X_6504__48 VPWR VGND net48 sg13g2_tiehi
XFILLER_49_148 VPWR VGND sg13g2_fill_2
Xfanout993 _2772_ net993 VPWR VGND sg13g2_buf_8
XFILLER_46_855 VPWR VGND sg13g2_decap_8
XFILLER_45_387 VPWR VGND sg13g2_decap_8
XFILLER_33_549 VPWR VGND sg13g2_fill_2
XFILLER_41_593 VPWR VGND sg13g2_fill_2
XFILLER_9_233 VPWR VGND sg13g2_fill_1
XFILLER_13_262 VPWR VGND sg13g2_fill_2
XFILLER_9_299 VPWR VGND sg13g2_decap_8
XFILLER_10_980 VPWR VGND sg13g2_decap_8
XFILLER_6_984 VPWR VGND sg13g2_decap_8
X_4210_ VGND VPWR _1741_ _1743_ _1745_ net1424 sg13g2_a21oi_1
X_6727__103 VPWR VGND net103 sg13g2_tiehi
X_5190_ s0.data_out\[0\]\[4\] s0.data_out\[1\]\[4\] net1033 _2629_ VPWR VGND sg13g2_mux2_1
X_4141_ _1679_ _1678_ _1677_ VPWR VGND sg13g2_nand2b_1
XFILLER_49_660 VPWR VGND sg13g2_decap_8
X_4072_ _1619_ _1618_ net1414 _1611_ net1405 VPWR VGND sg13g2_a22oi_1
X_4974_ VGND VPWR _2431_ _2435_ _0251_ _2436_ sg13g2_a21oi_1
XFILLER_24_549 VPWR VGND sg13g2_fill_1
X_6713_ net119 VGND VPWR _0223_ s0.data_out\[6\]\[7\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_3925_ VGND VPWR _1374_ _1490_ _1491_ net1185 sg13g2_a21oi_1
X_6644_ net193 VGND VPWR _0154_ s0.data_out\[11\]\[5\] clknet_leaf_22_clk sg13g2_dfrbpq_2
Xclkload8 VPWR clkload8/Y clknet_leaf_26_clk VGND sg13g2_inv_1
X_3856_ _0139_ _1429_ _1430_ _2832_ net1379 VPWR VGND sg13g2_a22oi_1
X_6575_ net268 VGND VPWR _0085_ s0.was_valid_out\[16\][0] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3787_ _1366_ net461 net1197 VPWR VGND sg13g2_nand2b_1
XFILLER_30_1024 VPWR VGND sg13g2_decap_4
X_5526_ VGND VPWR net1328 _2771_ _2932_ _2931_ sg13g2_a21oi_1
X_5457_ VPWR _2875_ net601 VGND sg13g2_inv_1
X_4408_ s0.data_out\[7\]\[1\] s0.data_out\[6\]\[1\] net1092 _1919_ VPWR VGND sg13g2_mux2_1
XFILLER_8_1003 VPWR VGND sg13g2_decap_8
X_5388_ VPWR _2806_ net511 VGND sg13g2_inv_1
X_4339_ net1102 net1158 _1862_ VPWR VGND sg13g2_nor2b_1
X_6009_ _0570_ net1271 net418 VPWR VGND sg13g2_nand2_1
XFILLER_28_877 VPWR VGND sg13g2_decap_8
XFILLER_43_836 VPWR VGND sg13g2_fill_1
XFILLER_15_538 VPWR VGND sg13g2_decap_4
XFILLER_23_571 VPWR VGND sg13g2_fill_1
XFILLER_24_64 VPWR VGND sg13g2_decap_8
XFILLER_10_254 VPWR VGND sg13g2_decap_4
XFILLER_11_777 VPWR VGND sg13g2_fill_1
XFILLER_3_943 VPWR VGND sg13g2_decap_8
XFILLER_49_94 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_17 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_45_140 VPWR VGND sg13g2_fill_2
XFILLER_45_173 VPWR VGND sg13g2_fill_1
XFILLER_34_858 VPWR VGND sg13g2_fill_2
XFILLER_33_357 VPWR VGND sg13g2_fill_1
XFILLER_42_891 VPWR VGND sg13g2_fill_2
X_3710_ _1220_ _1298_ _1299_ _1300_ VPWR VGND sg13g2_nor3_1
X_4690_ s0.data_out\[5\]\[7\] s0.data_out\[4\]\[7\] net1070 _2177_ VPWR VGND sg13g2_mux2_1
X_3641_ VGND VPWR _1116_ _1230_ _1231_ net1204 sg13g2_a21oi_1
X_6360_ _0885_ VPWR _0888_ VGND net362 net1233 sg13g2_o21ai_1
X_3572_ _1173_ VPWR _1174_ VGND net1441 _1145_ sg13g2_o21ai_1
X_5311_ VPWR _2729_ net356 VGND sg13g2_inv_1
XFILLER_5_291 VPWR VGND sg13g2_fill_2
X_6291_ VGND VPWR _0828_ _0826_ net1411 sg13g2_or2_1
X_5242_ _2674_ VPWR _2675_ VGND net1006 _2673_ sg13g2_o21ai_1
X_5173_ s0.data_out\[0\]\[7\] s0.data_out\[1\]\[7\] net1034 _2612_ VPWR VGND sg13g2_mux2_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
X_4124_ _1665_ VPWR _1666_ VGND net1490 net610 sg13g2_o21ai_1
XFILLER_28_107 VPWR VGND sg13g2_decap_8
XFILLER_49_490 VPWR VGND sg13g2_decap_8
X_4055_ _1602_ net1442 _1598_ VPWR VGND sg13g2_nand2_1
XFILLER_40_828 VPWR VGND sg13g2_fill_1
X_4957_ _2419_ VPWR _2420_ VGND net1438 _2393_ sg13g2_o21ai_1
X_4888_ net1052 VPWR _2354_ VGND net1397 net1040 sg13g2_o21ai_1
X_3908_ _1474_ _1473_ net1179 VPWR VGND sg13g2_nand2b_1
XFILLER_20_563 VPWR VGND sg13g2_decap_8
X_6627_ net211 VGND VPWR net443 s0.data_out\[12\]\[1\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3839_ net1178 s0.data_out\[11\]\[0\] _1417_ VPWR VGND sg13g2_and2_1
X_6558_ net286 VGND VPWR net411 s0.data_out\[18\]\[3\] clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_4_718 VPWR VGND sg13g2_decap_8
X_6489_ net1380 _0996_ _0997_ _0098_ VPWR VGND sg13g2_nor3_1
X_5509_ _2915_ net1321 net640 VPWR VGND sg13g2_nand2_1
Xfanout1029 s0.shift_out\[1\][0] net1029 VPWR VGND sg13g2_buf_8
XFILLER_0_957 VPWR VGND sg13g2_decap_8
Xfanout1018 _2741_ net1018 VPWR VGND sg13g2_buf_8
Xfanout1007 net1008 net1007 VPWR VGND sg13g2_buf_8
XFILLER_48_928 VPWR VGND sg13g2_decap_8
XFILLER_19_42 VPWR VGND sg13g2_decap_4
XFILLER_19_53 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_39_clk clknet_3_0__leaf_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_43_611 VPWR VGND sg13g2_fill_1
XFILLER_43_655 VPWR VGND sg13g2_decap_4
XFILLER_37_1008 VPWR VGND sg13g2_decap_8
XFILLER_11_541 VPWR VGND sg13g2_fill_1
XFILLER_7_523 VPWR VGND sg13g2_decap_8
XFILLER_3_740 VPWR VGND sg13g2_decap_8
XFILLER_32_7 VPWR VGND sg13g2_fill_2
XFILLER_47_983 VPWR VGND sg13g2_decap_8
X_5860_ net1286 net432 _0438_ VPWR VGND sg13g2_and2_1
XFILLER_18_162 VPWR VGND sg13g2_decap_4
XFILLER_18_195 VPWR VGND sg13g2_decap_8
X_4811_ _2284_ net1053 _2285_ _2286_ VPWR VGND sg13g2_a21o_1
X_5791_ _0376_ net473 net1308 VPWR VGND sg13g2_nand2b_1
X_4742_ net1073 VPWR _2225_ VGND _2158_ _2224_ sg13g2_o21ai_1
X_4673_ _2160_ net444 net1080 VPWR VGND sg13g2_nand2b_1
X_6412_ VGND VPWR _0813_ _0936_ _0937_ net1241 sg13g2_a21oi_1
X_3624_ net1208 VPWR _1217_ VGND net1395 net1196 sg13g2_o21ai_1
X_6343_ net1236 net475 _0874_ VPWR VGND sg13g2_and2_1
X_3555_ net1206 net1150 _1157_ VPWR VGND sg13g2_nor2b_1
X_3486_ _1094_ VPWR _1095_ VGND net1484 net643 sg13g2_o21ai_1
X_6274_ _0811_ _0810_ net1439 _0787_ net1447 VPWR VGND sg13g2_a22oi_1
X_5225_ VGND VPWR net1019 net386 _2661_ _2585_ sg13g2_a21oi_1
X_5156_ s0.data_out\[0\]\[0\] s0.data_out\[1\]\[0\] net1033 _2595_ VPWR VGND sg13g2_mux2_1
XFILLER_29_405 VPWR VGND sg13g2_decap_4
X_5087_ VGND VPWR _2532_ _2534_ _2538_ net1417 sg13g2_a21oi_1
X_4107_ VPWR _0168_ _1652_ VGND sg13g2_inv_1
X_4038_ net1124 net1164 _1585_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_471 VPWR VGND sg13g2_fill_1
XFILLER_40_603 VPWR VGND sg13g2_decap_8
XFILLER_13_817 VPWR VGND sg13g2_fill_2
X_5989_ net1274 VPWR _0553_ VGND net1393 net1261 sg13g2_o21ai_1
XFILLER_13_839 VPWR VGND sg13g2_fill_1
X_6675__160 VPWR VGND net160 sg13g2_tiehi
XFILLER_20_382 VPWR VGND sg13g2_decap_8
XFILLER_21_894 VPWR VGND sg13g2_fill_1
XFILLER_21_54 VPWR VGND sg13g2_fill_2
XFILLER_43_1012 VPWR VGND sg13g2_decap_8
XFILLER_0_754 VPWR VGND sg13g2_decap_8
XFILLER_48_725 VPWR VGND sg13g2_decap_8
XFILLER_47_257 VPWR VGND sg13g2_decap_8
XFILLER_28_471 VPWR VGND sg13g2_fill_2
XFILLER_29_994 VPWR VGND sg13g2_decap_8
XFILLER_44_953 VPWR VGND sg13g2_decap_8
XFILLER_15_121 VPWR VGND sg13g2_decap_4
XFILLER_15_143 VPWR VGND sg13g2_decap_8
X_6785__65 VPWR VGND net65 sg13g2_tiehi
X_6539__307 VPWR VGND net307 sg13g2_tiehi
XFILLER_30_124 VPWR VGND sg13g2_fill_1
XFILLER_11_393 VPWR VGND sg13g2_fill_2
XFILLER_7_364 VPWR VGND sg13g2_fill_1
XFILLER_7_397 VPWR VGND sg13g2_decap_4
Xhold309 _0044_ VPWR VGND net629 sg13g2_dlygate4sd3_1
X_5010_ net1392 net1034 _2464_ VPWR VGND sg13g2_nor2b_1
Xfanout1393 net1397 net1393 VPWR VGND sg13g2_buf_8
Xfanout1360 net1362 net1360 VPWR VGND sg13g2_buf_8
Xfanout1382 net1383 net1382 VPWR VGND sg13g2_buf_8
Xfanout1371 net1373 net1371 VPWR VGND sg13g2_buf_1
XFILLER_47_780 VPWR VGND sg13g2_decap_8
XFILLER_19_493 VPWR VGND sg13g2_fill_2
XFILLER_35_953 VPWR VGND sg13g2_decap_8
X_5912_ _0484_ VPWR _0485_ VGND _0475_ _0476_ sg13g2_o21ai_1
X_5843_ _0424_ VPWR _0425_ VGND net1007 _0423_ sg13g2_o21ai_1
X_6659__177 VPWR VGND net177 sg13g2_tiehi
X_5774_ _0359_ net1297 net628 VPWR VGND sg13g2_nand2_1
X_4725_ VGND VPWR _2212_ net1329 net331 sg13g2_or2_1
XFILLER_30_691 VPWR VGND sg13g2_fill_2
X_4656_ net1061 net1172 _2143_ VPWR VGND sg13g2_nor2b_1
X_4587_ _2086_ net999 _2085_ VPWR VGND sg13g2_nand2_1
X_3607_ VGND VPWR net1017 _1180_ _1204_ net1380 sg13g2_a21oi_1
XFILLER_1_507 VPWR VGND sg13g2_fill_1
X_3538_ _1139_ VPWR _1140_ VGND net1210 _2822_ sg13g2_o21ai_1
X_6326_ net1238 net479 _0861_ VPWR VGND sg13g2_and2_1
X_6257_ VGND VPWR _0680_ _0793_ _0794_ net1255 sg13g2_a21oi_1
X_3469_ _1081_ VPWR _1082_ VGND net1477 net607 sg13g2_o21ai_1
X_5208_ _2642_ _2638_ net1417 _2647_ VPWR VGND sg13g2_a21o_1
X_6188_ net1430 _0728_ _0737_ VPWR VGND sg13g2_nor2_1
XFILLER_29_202 VPWR VGND sg13g2_decap_4
X_5139_ VGND VPWR _2575_ _2578_ _2581_ _2580_ sg13g2_a21oi_1
XFILLER_29_279 VPWR VGND sg13g2_fill_2
XFILLER_26_964 VPWR VGND sg13g2_decap_8
XFILLER_41_945 VPWR VGND sg13g2_decap_8
X_6519__32 VPWR VGND net32 sg13g2_tiehi
XFILLER_8_128 VPWR VGND sg13g2_fill_2
XFILLER_32_86 VPWR VGND sg13g2_decap_8
XFILLER_10_1022 VPWR VGND sg13g2_decap_8
XFILLER_4_356 VPWR VGND sg13g2_fill_1
XFILLER_4_389 VPWR VGND sg13g2_fill_1
XFILLER_0_551 VPWR VGND sg13g2_decap_8
X_6545__300 VPWR VGND net300 sg13g2_tiehi
XFILLER_17_964 VPWR VGND sg13g2_decap_8
XFILLER_44_783 VPWR VGND sg13g2_decap_4
XFILLER_44_761 VPWR VGND sg13g2_fill_1
XFILLER_16_485 VPWR VGND sg13g2_fill_2
XFILLER_32_912 VPWR VGND sg13g2_fill_2
XFILLER_32_923 VPWR VGND sg13g2_decap_4
XFILLER_43_271 VPWR VGND sg13g2_fill_2
XFILLER_32_978 VPWR VGND sg13g2_decap_8
XFILLER_12_680 VPWR VGND sg13g2_fill_2
X_4510_ net1088 VPWR _2012_ VGND net1396 net1078 sg13g2_o21ai_1
X_5490_ net392 net1318 _2899_ VPWR VGND sg13g2_nor2_1
X_4441_ _1950_ net1089 _1951_ _1952_ VPWR VGND sg13g2_a21o_1
Xhold117 _0653_ VPWR VGND net437 sg13g2_dlygate4sd3_1
Xhold106 s0.data_out\[16\]\[2\] VPWR VGND net426 sg13g2_dlygate4sd3_1
XFILLER_7_194 VPWR VGND sg13g2_decap_4
Xhold139 s0.data_out\[23\]\[5\] VPWR VGND net459 sg13g2_dlygate4sd3_1
Xhold128 _0219_ VPWR VGND net448 sg13g2_dlygate4sd3_1
X_4372_ net1376 _1865_ _1890_ VPWR VGND sg13g2_nor2_1
X_6111_ _0663_ net1337 net1258 VPWR VGND sg13g2_nand2_1
XFILLER_39_500 VPWR VGND sg13g2_fill_2
X_6042_ net1261 net1148 _0603_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_0 VPWR VGND sg13g2_fill_1
XFILLER_27_717 VPWR VGND sg13g2_decap_8
Xfanout1190 s0.valid_out\[11\][0] net1190 VPWR VGND sg13g2_buf_8
XFILLER_26_205 VPWR VGND sg13g2_decap_4
XFILLER_35_750 VPWR VGND sg13g2_fill_1
XFILLER_19_290 VPWR VGND sg13g2_fill_1
XFILLER_34_271 VPWR VGND sg13g2_fill_1
X_5826_ _0405_ VPWR _0411_ VGND _0397_ _0408_ sg13g2_o21ai_1
XFILLER_33_1000 VPWR VGND sg13g2_decap_8
XFILLER_10_628 VPWR VGND sg13g2_fill_2
X_5757_ VGND VPWR net1305 _0339_ _0342_ _0341_ sg13g2_a21oi_1
XFILLER_22_488 VPWR VGND sg13g2_fill_1
X_4708_ _2195_ net1069 s0.data_out\[4\]\[5\] VPWR VGND sg13g2_nand2_1
X_6516__35 VPWR VGND net35 sg13g2_tiehi
X_6672__163 VPWR VGND net163 sg13g2_tiehi
X_5688_ _3082_ net1313 _3081_ VPWR VGND sg13g2_nand2b_1
X_4639_ _2126_ VPWR _2129_ VGND s0.was_valid_out\[4\][0] net1070 sg13g2_o21ai_1
XFILLER_2_805 VPWR VGND sg13g2_decap_8
X_6309_ _0722_ VPWR _0846_ VGND net1257 _2810_ sg13g2_o21ai_1
X_6529__317 VPWR VGND net317 sg13g2_tiehi
XFILLER_18_717 VPWR VGND sg13g2_fill_2
XFILLER_45_547 VPWR VGND sg13g2_fill_2
XFILLER_17_249 VPWR VGND sg13g2_fill_2
XFILLER_14_912 VPWR VGND sg13g2_fill_2
XFILLER_32_219 VPWR VGND sg13g2_fill_2
XFILLER_40_241 VPWR VGND sg13g2_fill_2
XFILLER_13_455 VPWR VGND sg13g2_decap_8
XFILLER_14_978 VPWR VGND sg13g2_decap_8
XFILLER_43_85 VPWR VGND sg13g2_fill_1
XFILLER_5_665 VPWR VGND sg13g2_fill_1
XFILLER_4_142 VPWR VGND sg13g2_fill_1
XFILLER_49_842 VPWR VGND sg13g2_decap_8
X_6649__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_48_330 VPWR VGND sg13g2_decap_8
XFILLER_36_536 VPWR VGND sg13g2_fill_1
X_4990_ net1348 _2392_ _2449_ VPWR VGND sg13g2_nor2_1
XFILLER_44_580 VPWR VGND sg13g2_fill_2
XFILLER_16_293 VPWR VGND sg13g2_fill_1
XFILLER_17_1006 VPWR VGND sg13g2_decap_8
X_3941_ _1507_ net1184 _1506_ VPWR VGND sg13g2_nand2b_1
X_6660_ net176 VGND VPWR _0170_ s0.data_out\[10\]\[2\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3872_ net1195 VPWR _1443_ VGND _1376_ _1442_ sg13g2_o21ai_1
X_5611_ _0012_ _3007_ _3008_ _2764_ net1339 VPWR VGND sg13g2_a22oi_1
XFILLER_20_948 VPWR VGND sg13g2_decap_8
X_6591_ net250 VGND VPWR _0101_ s0.data_out\[15\]\[0\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_5542_ net455 net1327 _2948_ VPWR VGND sg13g2_nor2b_1
XFILLER_9_982 VPWR VGND sg13g2_decap_8
X_5473_ VGND VPWR net1334 net992 net4 _2888_ sg13g2_a21oi_1
X_4424_ _1934_ VPWR _1935_ VGND net1093 _2857_ sg13g2_o21ai_1
X_4355_ _1821_ _1876_ net1481 _1877_ VPWR VGND sg13g2_nand3_1
X_4286_ _1808_ VPWR _1809_ VGND net1105 _2853_ sg13g2_o21ai_1
XFILLER_39_341 VPWR VGND sg13g2_fill_1
X_6025_ _0585_ VPWR _0586_ VGND net1270 _2794_ sg13g2_o21ai_1
XFILLER_27_525 VPWR VGND sg13g2_decap_8
XFILLER_23_720 VPWR VGND sg13g2_fill_2
X_5809_ _0394_ net1305 _0393_ VPWR VGND sg13g2_nand2b_1
XFILLER_11_948 VPWR VGND sg13g2_decap_8
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_2_679 VPWR VGND sg13g2_decap_8
XFILLER_38_30 VPWR VGND sg13g2_fill_2
Xfanout994 _2772_ net994 VPWR VGND sg13g2_buf_8
XFILLER_46_834 VPWR VGND sg13g2_decap_8
XFILLER_18_525 VPWR VGND sg13g2_fill_2
X_6542__303 VPWR VGND net303 sg13g2_tiehi
XFILLER_6_963 VPWR VGND sg13g2_decap_8
X_4140_ _1678_ net1338 net1121 VPWR VGND sg13g2_nand2_1
X_4071_ VGND VPWR net1139 _1615_ _1618_ _1617_ sg13g2_a21oi_1
XFILLER_36_333 VPWR VGND sg13g2_fill_2
XFILLER_36_355 VPWR VGND sg13g2_decap_8
XFILLER_24_528 VPWR VGND sg13g2_decap_4
X_4973_ VGND VPWR _2436_ net1330 net340 sg13g2_or2_1
XFILLER_36_388 VPWR VGND sg13g2_fill_2
X_6712_ net120 VGND VPWR _0222_ s0.data_out\[6\]\[6\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_3924_ _1490_ s0.data_out\[10\]\[7\] net1189 VPWR VGND sg13g2_nand2b_1
X_6643_ net194 VGND VPWR _0153_ s0.data_out\[11\]\[4\] clknet_leaf_23_clk sg13g2_dfrbpq_2
Xclkload9 clknet_leaf_20_clk clkload9/Y VPWR VGND sg13g2_inv_4
X_3855_ net1379 _1367_ _1430_ VPWR VGND sg13g2_nor2_1
X_6574_ net269 VGND VPWR _0084_ s0.data_out\[17\]\[7\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3786_ _1363_ net1180 _1364_ _1365_ VPWR VGND sg13g2_a21o_1
XFILLER_30_1003 VPWR VGND sg13g2_decap_8
X_5525_ _2770_ _2750_ net1326 _2931_ VPWR VGND sg13g2_a21o_1
X_5456_ VPWR _2874_ net484 VGND sg13g2_inv_1
X_4407_ _1918_ net1092 net501 VPWR VGND sg13g2_nand2_1
X_5387_ VPWR _2805_ net689 VGND sg13g2_inv_1
X_4338_ s0.data_out\[8\]\[4\] s0.data_out\[7\]\[4\] net1108 _1861_ VPWR VGND sg13g2_mux2_1
X_4269_ _1793_ VPWR _1795_ VGND s0.was_valid_out\[7\][0] net1107 sg13g2_o21ai_1
X_6008_ VGND VPWR _0569_ _0568_ net1443 sg13g2_or2_1
XFILLER_39_182 VPWR VGND sg13g2_fill_2
XFILLER_43_804 VPWR VGND sg13g2_decap_8
XFILLER_15_506 VPWR VGND sg13g2_decap_4
XFILLER_43_848 VPWR VGND sg13g2_decap_4
XFILLER_11_789 VPWR VGND sg13g2_decap_8
XFILLER_40_31 VPWR VGND sg13g2_fill_1
XFILLER_3_922 VPWR VGND sg13g2_decap_8
XFILLER_2_421 VPWR VGND sg13g2_fill_1
XFILLER_3_999 VPWR VGND sg13g2_decap_8
XFILLER_49_51 VPWR VGND sg13g2_fill_1
XFILLER_37_108 VPWR VGND sg13g2_decap_4
XFILLER_19_801 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_18 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_18_311 VPWR VGND sg13g2_fill_2
XFILLER_46_675 VPWR VGND sg13g2_decap_8
XFILLER_19_889 VPWR VGND sg13g2_fill_2
XFILLER_34_804 VPWR VGND sg13g2_decap_8
XFILLER_45_185 VPWR VGND sg13g2_fill_1
XFILLER_33_314 VPWR VGND sg13g2_decap_4
XFILLER_42_881 VPWR VGND sg13g2_fill_1
XFILLER_41_380 VPWR VGND sg13g2_fill_2
X_3640_ _1230_ s0.data_out\[12\]\[2\] net1212 VPWR VGND sg13g2_nand2b_1
X_3571_ _1170_ _1172_ net1423 _1173_ VPWR VGND sg13g2_nand3_1
X_5310_ VGND VPWR net1467 _2716_ _0295_ _2728_ sg13g2_a21oi_1
X_6290_ _0827_ _0826_ net1411 _0819_ net1402 VPWR VGND sg13g2_a22oi_1
X_5241_ VGND VPWR net1006 _2637_ _2674_ net1347 sg13g2_a21oi_1
X_5172_ _2610_ VPWR _2611_ VGND _2602_ _2603_ sg13g2_o21ai_1
X_4123_ _1664_ VPWR _1665_ VGND net1013 _1663_ sg13g2_o21ai_1
X_4054_ _1582_ _1591_ _1599_ _1600_ _1601_ VPWR VGND sg13g2_nor4_1
XFILLER_37_686 VPWR VGND sg13g2_fill_2
XFILLER_36_130 VPWR VGND sg13g2_fill_1
X_4956_ _2419_ net1419 _2418_ VPWR VGND sg13g2_nand2_1
X_4887_ _0247_ _2352_ _2353_ _2869_ net1361 VPWR VGND sg13g2_a22oi_1
X_3907_ s0.data_out\[10\]\[0\] s0.data_out\[11\]\[0\] net1187 _1473_ VPWR VGND sg13g2_mux2_1
X_6626_ net212 VGND VPWR _0136_ s0.data_out\[12\]\[0\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3838_ VGND VPWR _1411_ _1415_ _0135_ _1416_ sg13g2_a21oi_1
X_6557_ net287 VGND VPWR net429 s0.data_out\[18\]\[2\] clknet_leaf_35_clk sg13g2_dfrbpq_2
XFILLER_3_218 VPWR VGND sg13g2_decap_4
X_5508_ VGND VPWR net1328 _2776_ _2914_ _2913_ sg13g2_a21oi_1
X_3769_ s0.data_out\[12\]\[0\] s0.data_out\[11\]\[0\] net1187 _1348_ VPWR VGND sg13g2_mux2_1
X_6488_ VGND VPWR _2735_ _0998_ _0097_ _1003_ sg13g2_a21oi_1
X_5439_ VPWR _2857_ net632 VGND sg13g2_inv_1
XFILLER_0_936 VPWR VGND sg13g2_decap_8
Xfanout1008 _2752_ net1008 VPWR VGND sg13g2_buf_8
Xfanout1019 net1021 net1019 VPWR VGND sg13g2_buf_8
XFILLER_48_907 VPWR VGND sg13g2_decap_8
XFILLER_47_406 VPWR VGND sg13g2_fill_1
XFILLER_15_303 VPWR VGND sg13g2_fill_1
XFILLER_28_686 VPWR VGND sg13g2_decap_8
XFILLER_27_196 VPWR VGND sg13g2_decap_8
XFILLER_24_870 VPWR VGND sg13g2_decap_4
X_6717__114 VPWR VGND net114 sg13g2_tiehi
XFILLER_11_597 VPWR VGND sg13g2_decap_8
XFILLER_3_796 VPWR VGND sg13g2_decap_8
XFILLER_2_262 VPWR VGND sg13g2_decap_8
X_6724__107 VPWR VGND net107 sg13g2_tiehi
XFILLER_47_962 VPWR VGND sg13g2_decap_8
XFILLER_19_664 VPWR VGND sg13g2_fill_1
XFILLER_19_675 VPWR VGND sg13g2_fill_2
X_4810_ net1053 net1143 _2285_ VPWR VGND sg13g2_nor2b_1
X_5790_ _0373_ net1286 _0374_ _0375_ VPWR VGND sg13g2_a21o_1
X_4741_ net995 _2871_ _2224_ VPWR VGND sg13g2_nor2_1
X_4672_ _2157_ net1062 _2158_ _2159_ VPWR VGND sg13g2_a21o_1
X_6411_ _0936_ s0.data_out\[15\]\[7\] net1247 VPWR VGND sg13g2_nand2b_1
X_3623_ _0120_ _1215_ _1216_ _2819_ net1381 VPWR VGND sg13g2_a22oi_1
XFILLER_6_590 VPWR VGND sg13g2_decap_4
X_6342_ VPWR _0081_ _0873_ VGND sg13g2_inv_1
X_3554_ _1155_ VPWR _1156_ VGND net1211 _2820_ sg13g2_o21ai_1
X_3485_ _1069_ _1093_ net1484 _1094_ VPWR VGND sg13g2_nand3_1
X_6273_ VGND VPWR net1254 _0807_ _0810_ _0809_ sg13g2_a21oi_1
X_5224_ _0277_ _2659_ _2660_ _2884_ net1346 VPWR VGND sg13g2_a22oi_1
XFILLER_5_1018 VPWR VGND sg13g2_decap_8
X_5155_ VGND VPWR net1029 _2593_ _2594_ _2590_ sg13g2_a21oi_1
X_5086_ VGND VPWR _2525_ _2527_ _2537_ net1429 sg13g2_a21oi_1
X_4106_ _1651_ VPWR _1652_ VGND net1488 net626 sg13g2_o21ai_1
XFILLER_38_984 VPWR VGND sg13g2_decap_8
X_4037_ s0.data_out\[10\]\[2\] s0.data_out\[9\]\[2\] net1133 _1584_ VPWR VGND sg13g2_mux2_1
X_5988_ _0048_ _0551_ _0552_ _2784_ net1353 VPWR VGND sg13g2_a22oi_1
XFILLER_13_829 VPWR VGND sg13g2_fill_2
XFILLER_24_155 VPWR VGND sg13g2_fill_2
XFILLER_25_678 VPWR VGND sg13g2_decap_4
X_4939_ _2402_ net1045 net580 VPWR VGND sg13g2_nand2_1
XFILLER_21_873 VPWR VGND sg13g2_fill_1
X_6609_ net231 VGND VPWR net546 s0.data_out\[14\]\[6\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_0_733 VPWR VGND sg13g2_decap_8
XFILLER_48_704 VPWR VGND sg13g2_decap_8
XFILLER_29_973 VPWR VGND sg13g2_decap_8
XFILLER_46_63 VPWR VGND sg13g2_fill_1
XFILLER_44_932 VPWR VGND sg13g2_decap_8
XFILLER_15_100 VPWR VGND sg13g2_fill_1
XFILLER_15_111 VPWR VGND sg13g2_fill_2
XFILLER_43_464 VPWR VGND sg13g2_fill_1
XFILLER_31_637 VPWR VGND sg13g2_fill_2
XFILLER_8_822 VPWR VGND sg13g2_decap_4
X_6730__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_38_203 VPWR VGND sg13g2_fill_1
XFILLER_23_4 VPWR VGND sg13g2_decap_8
Xfanout1350 net1351 net1350 VPWR VGND sg13g2_buf_8
Xfanout1372 net1373 net1372 VPWR VGND sg13g2_buf_8
XFILLER_39_737 VPWR VGND sg13g2_fill_1
Xfanout1361 net1362 net1361 VPWR VGND sg13g2_buf_1
Xfanout1383 net1389 net1383 VPWR VGND sg13g2_buf_8
Xfanout1394 net1396 net1394 VPWR VGND sg13g2_buf_8
XFILLER_35_910 VPWR VGND sg13g2_fill_1
X_5911_ _0484_ _0483_ net1437 _0460_ net1444 VPWR VGND sg13g2_a22oi_1
X_5842_ VGND VPWR net1007 _0354_ _0424_ net1345 sg13g2_a21oi_1
XFILLER_34_453 VPWR VGND sg13g2_fill_2
X_5773_ _0358_ net1334 _0356_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_136 VPWR VGND sg13g2_decap_8
X_4724_ _2209_ _2210_ _2211_ VPWR VGND sg13g2_nor2_1
X_4655_ _2142_ _2141_ net1072 VPWR VGND sg13g2_nand2b_1
X_4586_ s0.data_out\[5\]\[5\] s0.data_out\[6\]\[5\] net1095 _2085_ VPWR VGND sg13g2_mux2_1
X_3606_ VGND VPWR net1204 net491 _1203_ _1176_ sg13g2_a21oi_1
X_3537_ _1139_ net1210 net532 VPWR VGND sg13g2_nand2_1
X_6325_ VPWR _0077_ _0860_ VGND sg13g2_inv_1
XFILLER_1_519 VPWR VGND sg13g2_decap_8
X_6256_ _0793_ net479 net1260 VPWR VGND sg13g2_nand2b_1
X_3468_ _1024_ _1080_ net1477 _1081_ VPWR VGND sg13g2_nand3_1
X_5207_ VGND VPWR _2638_ _2642_ _2646_ net1417 sg13g2_a21oi_1
X_6187_ _0736_ _0735_ net1421 _0728_ net1430 VPWR VGND sg13g2_a22oi_1
X_3399_ _1013_ net1219 net647 VPWR VGND sg13g2_nand2_1
X_5138_ _2579_ VPWR _2580_ VGND net1022 _2574_ sg13g2_o21ai_1
XFILLER_29_236 VPWR VGND sg13g2_decap_8
XFILLER_45_707 VPWR VGND sg13g2_decap_4
X_5069_ net1399 _2511_ _2520_ VPWR VGND sg13g2_nor2_1
XFILLER_26_943 VPWR VGND sg13g2_decap_8
XFILLER_13_615 VPWR VGND sg13g2_fill_1
XFILLER_13_648 VPWR VGND sg13g2_fill_1
XFILLER_32_21 VPWR VGND sg13g2_fill_1
XFILLER_4_302 VPWR VGND sg13g2_fill_1
XFILLER_10_1001 VPWR VGND sg13g2_decap_8
XFILLER_0_530 VPWR VGND sg13g2_decap_8
XFILLER_17_910 VPWR VGND sg13g2_fill_1
XFILLER_17_921 VPWR VGND sg13g2_decap_8
XFILLER_43_250 VPWR VGND sg13g2_fill_1
XFILLER_32_957 VPWR VGND sg13g2_decap_8
X_4440_ net1089 net1144 _1951_ VPWR VGND sg13g2_nor2b_1
Xhold107 s0.was_valid_out\[0\][0] VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold129 s0.data_out\[5\]\[6\] VPWR VGND net449 sg13g2_dlygate4sd3_1
Xhold118 s0.data_out\[23\]\[7\] VPWR VGND net438 sg13g2_dlygate4sd3_1
X_4371_ net1114 VPWR _1889_ VGND _1862_ _1888_ sg13g2_o21ai_1
XFILLER_4_880 VPWR VGND sg13g2_decap_8
X_6110_ net1262 VPWR _0662_ VGND net1394 net1249 sg13g2_o21ai_1
X_6041_ s0.data_out\[19\]\[6\] s0.data_out\[18\]\[6\] net1269 _0602_ VPWR VGND sg13g2_mux2_1
X_6665__171 VPWR VGND net171 sg13g2_tiehi
Xfanout1191 net1192 net1191 VPWR VGND sg13g2_buf_8
XFILLER_27_707 VPWR VGND sg13g2_fill_2
Xfanout1180 net1181 net1180 VPWR VGND sg13g2_buf_8
X_5825_ _0371_ _0389_ _0406_ _0409_ _0410_ VPWR VGND sg13g2_or4_1
X_5756_ VGND VPWR _3017_ _0340_ _0341_ net1306 sg13g2_a21oi_1
X_4707_ _2191_ _2193_ net1427 _2194_ VPWR VGND sg13g2_nand3_1
X_5687_ VGND VPWR net1300 _3079_ _3081_ _3080_ sg13g2_a21oi_1
X_4638_ _2126_ _2127_ _2128_ VPWR VGND sg13g2_nor2_1
X_4569_ VGND VPWR _1942_ _2067_ _2068_ net1088 sg13g2_a21oi_1
XFILLER_1_305 VPWR VGND sg13g2_fill_1
X_6308_ _0845_ net1250 _0844_ VPWR VGND sg13g2_nand2b_1
X_6239_ _0779_ _0776_ _0778_ VPWR VGND sg13g2_nand2_1
XFILLER_40_1027 VPWR VGND sg13g2_fill_2
XFILLER_40_1016 VPWR VGND sg13g2_decap_8
XFILLER_26_784 VPWR VGND sg13g2_fill_2
XFILLER_14_935 VPWR VGND sg13g2_fill_2
XFILLER_14_957 VPWR VGND sg13g2_decap_8
XFILLER_25_272 VPWR VGND sg13g2_decap_8
XFILLER_9_427 VPWR VGND sg13g2_fill_2
XFILLER_40_297 VPWR VGND sg13g2_decap_4
XFILLER_49_821 VPWR VGND sg13g2_decap_8
XFILLER_0_393 VPWR VGND sg13g2_decap_8
XFILLER_49_898 VPWR VGND sg13g2_decap_8
XFILLER_1_1010 VPWR VGND sg13g2_decap_8
X_3940_ VGND VPWR net1140 _1504_ _1506_ _1505_ sg13g2_a21oi_1
XFILLER_17_795 VPWR VGND sg13g2_fill_2
X_3871_ net1182 net451 _1442_ VPWR VGND sg13g2_and2_1
X_6590_ net251 VGND VPWR _0100_ s0.shift_out\[15\][0] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_5610_ net1339 _2942_ _3008_ VPWR VGND sg13g2_nor2_1
X_5541_ VGND VPWR net1323 _2946_ _2947_ _2942_ sg13g2_a21oi_1
XFILLER_9_961 VPWR VGND sg13g2_decap_8
XFILLER_8_460 VPWR VGND sg13g2_decap_8
X_5472_ s0.data_out\[23\]\[2\] net992 _2888_ VPWR VGND sg13g2_nor2_1
X_6513__39 VPWR VGND net39 sg13g2_tiehi
X_4423_ _1934_ net1093 net389 VPWR VGND sg13g2_nand2_1
X_4354_ net1110 VPWR _1876_ VGND _1817_ _1875_ sg13g2_o21ai_1
X_6024_ _0585_ net1270 net410 VPWR VGND sg13g2_nand2_1
X_4285_ _1808_ net1105 net408 VPWR VGND sg13g2_nand2_1
XFILLER_35_570 VPWR VGND sg13g2_fill_2
XFILLER_11_938 VPWR VGND sg13g2_fill_1
X_5808_ VGND VPWR net1292 _0392_ _0393_ _0390_ sg13g2_a21oi_1
XFILLER_22_253 VPWR VGND sg13g2_decap_4
X_5739_ net1393 _2753_ _0327_ VPWR VGND sg13g2_nor2_1
XFILLER_10_459 VPWR VGND sg13g2_decap_8
X_6535__311 VPWR VGND net311 sg13g2_tiehi
XFILLER_2_658 VPWR VGND sg13g2_decap_8
Xfanout995 _2762_ net995 VPWR VGND sg13g2_buf_8
XFILLER_46_813 VPWR VGND sg13g2_decap_8
XFILLER_14_732 VPWR VGND sg13g2_fill_2
XFILLER_14_776 VPWR VGND sg13g2_fill_2
XFILLER_41_595 VPWR VGND sg13g2_fill_1
X_6655__181 VPWR VGND net181 sg13g2_tiehi
XFILLER_6_942 VPWR VGND sg13g2_decap_8
X_6503__50 VPWR VGND net50 sg13g2_tiehi
XFILLER_5_485 VPWR VGND sg13g2_decap_4
X_4070_ VGND VPWR _1493_ _1616_ _1617_ net1138 sg13g2_a21oi_1
XFILLER_23_1022 VPWR VGND sg13g2_decap_8
XFILLER_49_695 VPWR VGND sg13g2_decap_8
X_6662__174 VPWR VGND net174 sg13g2_tiehi
X_4972_ _2357_ _2433_ _2434_ _2435_ VPWR VGND sg13g2_nor3_1
XFILLER_17_570 VPWR VGND sg13g2_fill_1
X_6711_ net121 VGND VPWR _0221_ s0.data_out\[6\]\[5\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_3923_ _1487_ net1138 _1488_ _1489_ VPWR VGND sg13g2_a21o_1
X_3854_ net1193 VPWR _1429_ VGND _1364_ _1428_ sg13g2_o21ai_1
X_6642_ net195 VGND VPWR net462 s0.data_out\[11\]\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_6573_ net270 VGND VPWR _0083_ s0.data_out\[17\]\[6\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3785_ net1180 net1161 _1364_ VPWR VGND sg13g2_nor2b_1
X_5524_ VGND VPWR _2920_ _2928_ _2930_ _2929_ sg13g2_a21oi_1
X_5455_ VPWR _2873_ net642 VGND sg13g2_inv_1
X_4406_ net1447 _1916_ _1917_ VPWR VGND sg13g2_nor2_1
X_5386_ VPWR _2804_ net368 VGND sg13g2_inv_1
X_4337_ _1860_ net1422 _1859_ VPWR VGND sg13g2_nand2_1
X_4268_ VGND VPWR _2759_ _1678_ _1794_ _1793_ sg13g2_a21oi_1
X_6007_ VGND VPWR net1278 _0565_ _0568_ _0567_ sg13g2_a21oi_1
X_4199_ net1414 _1725_ _1734_ VPWR VGND sg13g2_nor2_1
XFILLER_24_11 VPWR VGND sg13g2_decap_4
XFILLER_24_33 VPWR VGND sg13g2_decap_4
XFILLER_10_234 VPWR VGND sg13g2_decap_8
XFILLER_11_768 VPWR VGND sg13g2_decap_8
X_6639__198 VPWR VGND net198 sg13g2_tiehi
XFILLER_3_901 VPWR VGND sg13g2_decap_8
XFILLER_3_978 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
Xhold290 s0.data_out\[10\]\[4\] VPWR VGND net610 sg13g2_dlygate4sd3_1
X_6500__53 VPWR VGND net53 sg13g2_tiehi
XFILLER_19_824 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_19 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_19_857 VPWR VGND sg13g2_fill_1
XFILLER_45_131 VPWR VGND sg13g2_decap_4
XFILLER_18_356 VPWR VGND sg13g2_fill_2
XFILLER_34_827 VPWR VGND sg13g2_fill_2
XFILLER_18_378 VPWR VGND sg13g2_fill_1
XFILLER_34_838 VPWR VGND sg13g2_fill_2
XFILLER_41_392 VPWR VGND sg13g2_fill_1
X_3570_ _1172_ _2741_ _1171_ VPWR VGND sg13g2_nand2_1
X_5240_ VGND VPWR net1023 net395 _2673_ _2640_ sg13g2_a21oi_1
XFILLER_5_271 VPWR VGND sg13g2_fill_1
XFILLER_5_293 VPWR VGND sg13g2_fill_1
X_5171_ _2610_ _2609_ net1436 _2588_ net1443 VPWR VGND sg13g2_a22oi_1
X_4122_ VGND VPWR net1013 _1628_ _1664_ net1387 sg13g2_a21oi_1
X_4053_ net1455 _1574_ _1600_ VPWR VGND sg13g2_nor2_1
XFILLER_24_315 VPWR VGND sg13g2_fill_2
X_4955_ VGND VPWR net1051 _2415_ _2418_ _2417_ sg13g2_a21oi_1
X_3906_ _1472_ net1179 _1471_ VPWR VGND sg13g2_nand2b_1
X_4886_ net1360 _2288_ _2353_ VPWR VGND sg13g2_nor2_1
X_6625_ net213 VGND VPWR _0135_ s0.shift_out\[12\][0] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_3837_ VGND VPWR _1416_ net1331 net342 sg13g2_or2_1
X_6556_ net288 VGND VPWR net419 s0.data_out\[18\]\[1\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3768_ net1178 net1171 _1347_ VPWR VGND sg13g2_nor2b_1
X_5507_ _2775_ _2750_ net1325 _2913_ VPWR VGND sg13g2_a21o_1
X_6532__314 VPWR VGND net314 sg13g2_tiehi
X_6487_ net1484 VPWR _1003_ VGND _1000_ _1002_ sg13g2_o21ai_1
X_3699_ VGND VPWR net1205 _1286_ _1289_ _1288_ sg13g2_a21oi_1
X_5438_ VPWR _2856_ net470 VGND sg13g2_inv_1
XFILLER_0_915 VPWR VGND sg13g2_decap_8
X_5369_ _2787_ net496 VPWR VGND sg13g2_inv_2
Xfanout1009 net1010 net1009 VPWR VGND sg13g2_buf_8
XFILLER_19_11 VPWR VGND sg13g2_fill_1
XFILLER_19_22 VPWR VGND sg13g2_fill_2
XFILLER_19_77 VPWR VGND sg13g2_decap_8
XFILLER_42_178 VPWR VGND sg13g2_fill_2
XFILLER_23_392 VPWR VGND sg13g2_decap_8
X_6652__184 VPWR VGND net184 sg13g2_tiehi
XFILLER_3_775 VPWR VGND sg13g2_decap_8
XFILLER_32_9 VPWR VGND sg13g2_fill_1
XFILLER_25_8 VPWR VGND sg13g2_fill_2
XFILLER_47_941 VPWR VGND sg13g2_decap_8
XFILLER_18_120 VPWR VGND sg13g2_decap_8
XFILLER_20_1025 VPWR VGND sg13g2_decap_4
XFILLER_19_687 VPWR VGND sg13g2_fill_2
XFILLER_15_860 VPWR VGND sg13g2_fill_1
XFILLER_15_871 VPWR VGND sg13g2_fill_2
XFILLER_14_381 VPWR VGND sg13g2_decap_4
X_4740_ VPWR _0230_ _2223_ VGND sg13g2_inv_1
XFILLER_30_841 VPWR VGND sg13g2_fill_2
X_4671_ net1062 net993 _2158_ VPWR VGND sg13g2_nor2_1
X_6410_ _0933_ net1224 _0934_ _0935_ VPWR VGND sg13g2_a21o_1
X_3622_ net1381 _1153_ _1216_ VPWR VGND sg13g2_nor2_1
X_6341_ _0872_ VPWR _0873_ VGND net1478 net668 sg13g2_o21ai_1
X_3553_ _1155_ net1211 s0.data_out\[13\]\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_44_0 VPWR VGND sg13g2_decap_4
X_3484_ net1230 VPWR _1093_ VGND _1065_ _1092_ sg13g2_o21ai_1
X_6272_ VGND VPWR _0696_ _0808_ _0809_ net1254 sg13g2_a21oi_1
X_5223_ net1346 _2590_ _2660_ VPWR VGND sg13g2_nor2_1
X_5154_ _2591_ net1020 _2592_ _2593_ VPWR VGND sg13g2_a21o_1
X_4105_ _1576_ _1650_ net1488 _1651_ VPWR VGND sg13g2_nand3_1
X_5085_ _2536_ _2528_ _2535_ VPWR VGND sg13g2_nand2_1
XFILLER_38_963 VPWR VGND sg13g2_decap_8
X_4036_ _1583_ net1131 net465 VPWR VGND sg13g2_nand2_1
XFILLER_37_462 VPWR VGND sg13g2_decap_8
XFILLER_24_101 VPWR VGND sg13g2_decap_8
XFILLER_13_808 VPWR VGND sg13g2_fill_1
XFILLER_36_1021 VPWR VGND sg13g2_decap_8
X_5987_ net1353 _0491_ _0552_ VPWR VGND sg13g2_nor2_1
X_4938_ VGND VPWR net1051 _2398_ _2401_ _2400_ sg13g2_a21oi_1
X_4869_ _0243_ _2338_ _2339_ _2871_ net1358 VPWR VGND sg13g2_a22oi_1
X_6608_ net232 VGND VPWR _0118_ s0.data_out\[14\]\[5\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_6539_ net307 VGND VPWR net367 s0.was_valid_out\[19\][0] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_0_712 VPWR VGND sg13g2_decap_8
XFILLER_0_789 VPWR VGND sg13g2_decap_8
XFILLER_29_952 VPWR VGND sg13g2_decap_8
XFILLER_44_911 VPWR VGND sg13g2_decap_8
XFILLER_16_613 VPWR VGND sg13g2_fill_1
XFILLER_16_635 VPWR VGND sg13g2_fill_1
XFILLER_44_988 VPWR VGND sg13g2_decap_8
XFILLER_8_845 VPWR VGND sg13g2_decap_8
XFILLER_11_351 VPWR VGND sg13g2_fill_1
XFILLER_3_561 VPWR VGND sg13g2_fill_1
Xfanout1340 net1343 net1340 VPWR VGND sg13g2_buf_8
Xfanout1362 net1364 net1362 VPWR VGND sg13g2_buf_1
Xfanout1384 net1388 net1384 VPWR VGND sg13g2_buf_8
Xfanout1351 net1389 net1351 VPWR VGND sg13g2_buf_8
Xfanout1373 net1377 net1373 VPWR VGND sg13g2_buf_8
Xfanout1395 net1396 net1395 VPWR VGND sg13g2_buf_8
X_5910_ VGND VPWR net1294 _0480_ _0483_ _0482_ sg13g2_a21oi_1
XFILLER_19_473 VPWR VGND sg13g2_fill_1
XFILLER_35_988 VPWR VGND sg13g2_decap_8
X_5841_ VGND VPWR net1291 net424 _0423_ _0350_ sg13g2_a21oi_1
X_5772_ VGND VPWR _0357_ _0356_ net1334 sg13g2_or2_1
X_4723_ _2128_ VPWR _2210_ VGND _2183_ _2185_ sg13g2_o21ai_1
X_4654_ s0.data_out\[4\]\[0\] s0.data_out\[5\]\[0\] net1080 _2141_ VPWR VGND sg13g2_mux2_1
X_4585_ _2084_ net1090 _2083_ VPWR VGND sg13g2_nand2b_1
X_3605_ _0116_ _1201_ _1202_ _2822_ net1378 VPWR VGND sg13g2_a22oi_1
X_3536_ _1123_ VPWR _1138_ VGND net1454 _1130_ sg13g2_o21ai_1
X_6324_ _0859_ VPWR _0860_ VGND net1478 net653 sg13g2_o21ai_1
X_6255_ _0791_ net1239 _0789_ _0792_ VPWR VGND sg13g2_a21o_1
X_3467_ net1228 VPWR _1080_ VGND _1020_ _1079_ sg13g2_o21ai_1
X_5206_ net1436 _2609_ _2645_ VPWR VGND sg13g2_nor2_1
X_6186_ VGND VPWR net1263 _0732_ _0735_ _0734_ sg13g2_a21oi_1
X_3398_ net1213 net1168 _1012_ VPWR VGND sg13g2_nor2b_1
X_5137_ net1006 VPWR _2579_ VGND net427 net1034 sg13g2_o21ai_1
X_6707__125 VPWR VGND net125 sg13g2_tiehi
X_5068_ VGND VPWR _2519_ _2517_ net1408 sg13g2_or2_1
XFILLER_44_229 VPWR VGND sg13g2_fill_1
X_4019_ net1147 net1407 net1390 _0165_ VPWR VGND sg13g2_mux2_1
XFILLER_37_270 VPWR VGND sg13g2_fill_2
X_6767__23 VPWR VGND net23 sg13g2_tiehi
XFILLER_26_999 VPWR VGND sg13g2_decap_8
XFILLER_40_413 VPWR VGND sg13g2_decap_4
XFILLER_25_498 VPWR VGND sg13g2_decap_4
XFILLER_32_44 VPWR VGND sg13g2_fill_1
X_6714__118 VPWR VGND net118 sg13g2_tiehi
XFILLER_5_848 VPWR VGND sg13g2_fill_2
XFILLER_48_524 VPWR VGND sg13g2_decap_4
XFILLER_0_586 VPWR VGND sg13g2_decap_8
XFILLER_35_207 VPWR VGND sg13g2_fill_2
XFILLER_16_465 VPWR VGND sg13g2_decap_4
XFILLER_17_999 VPWR VGND sg13g2_decap_8
XFILLER_31_402 VPWR VGND sg13g2_fill_2
XFILLER_16_487 VPWR VGND sg13g2_fill_1
XFILLER_16_498 VPWR VGND sg13g2_fill_1
X_6771__267 VPWR VGND net267 sg13g2_tiehi
X_6525__26 VPWR VGND net26 sg13g2_tiehi
Xhold108 s0.data_out\[18\]\[2\] VPWR VGND net428 sg13g2_dlygate4sd3_1
X_4370_ net1102 net639 _1888_ VPWR VGND sg13g2_and2_1
Xhold119 _0012_ VPWR VGND net439 sg13g2_dlygate4sd3_1
X_6040_ _0601_ net1272 net534 VPWR VGND sg13g2_nand2_1
XFILLER_26_1020 VPWR VGND sg13g2_decap_8
Xfanout1192 net1193 net1192 VPWR VGND sg13g2_buf_1
Xfanout1170 net1173 net1170 VPWR VGND sg13g2_buf_8
Xfanout1181 net1186 net1181 VPWR VGND sg13g2_buf_8
X_5824_ VGND VPWR _0409_ _0408_ _0407_ sg13g2_or2_1
XFILLER_23_947 VPWR VGND sg13g2_decap_4
X_6776__189 VPWR VGND net189 sg13g2_tiehi
X_5755_ _0340_ s0.data_out\[20\]\[1\] net1309 VPWR VGND sg13g2_nand2b_1
X_4706_ _2193_ _2192_ net1073 VPWR VGND sg13g2_nand2b_1
X_5686_ net1300 net1151 _3080_ VPWR VGND sg13g2_nor2b_1
X_4637_ VGND VPWR net1336 net1082 _2127_ net1076 sg13g2_a21oi_1
X_4568_ _2067_ net449 net1094 VPWR VGND sg13g2_nand2b_1
X_4499_ net1372 _1964_ _2004_ VPWR VGND sg13g2_nor2_1
X_6307_ VGND VPWR net1237 _0843_ _0844_ _0841_ sg13g2_a21oi_1
X_3519_ VGND VPWR _1004_ _1120_ _1121_ net1216 sg13g2_a21oi_1
X_6238_ net1002 VPWR _0778_ VGND net370 net1257 sg13g2_o21ai_1
X_6169_ _0718_ _0717_ net1411 _0710_ net1402 VPWR VGND sg13g2_a22oi_1
XFILLER_17_218 VPWR VGND sg13g2_fill_2
X_6720__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_41_700 VPWR VGND sg13g2_fill_1
XFILLER_14_914 VPWR VGND sg13g2_fill_1
XFILLER_41_722 VPWR VGND sg13g2_fill_2
XFILLER_41_766 VPWR VGND sg13g2_fill_2
XFILLER_40_243 VPWR VGND sg13g2_fill_1
XFILLER_25_295 VPWR VGND sg13g2_fill_1
XFILLER_43_76 VPWR VGND sg13g2_fill_2
XFILLER_22_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_20_clk clknet_3_7__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
X_6522__29 VPWR VGND net29 sg13g2_tiehi
XFILLER_49_800 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_4
XFILLER_1_884 VPWR VGND sg13g2_decap_8
XFILLER_49_877 VPWR VGND sg13g2_decap_8
XFILLER_32_700 VPWR VGND sg13g2_decap_4
X_3870_ _0142_ _1440_ _1441_ _2831_ net1382 VPWR VGND sg13g2_a22oi_1
XFILLER_31_243 VPWR VGND sg13g2_fill_1
XFILLER_32_755 VPWR VGND sg13g2_fill_2
XFILLER_13_980 VPWR VGND sg13g2_decap_8
XFILLER_32_777 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_11_clk clknet_3_2__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_5540_ _2944_ net1311 _2945_ _2946_ VPWR VGND sg13g2_a21o_1
XFILLER_9_940 VPWR VGND sg13g2_decap_8
X_5471_ _2887_ VPWR net3 VGND _2776_ net992 sg13g2_o21ai_1
X_4422_ _1917_ _1931_ _1932_ _1933_ VPWR VGND sg13g2_nor3_1
X_4353_ net1098 s0.data_out\[7\]\[0\] _1875_ VPWR VGND sg13g2_and2_1
X_4284_ VGND VPWR _1807_ _1806_ net1446 sg13g2_or2_1
X_6023_ _0569_ VPWR _0584_ VGND net1452 _0576_ sg13g2_o21ai_1
X_6704__128 VPWR VGND net128 sg13g2_tiehi
XFILLER_23_722 VPWR VGND sg13g2_fill_1
X_3999_ net1137 VPWR _1556_ VGND net1396 net1129 sg13g2_o21ai_1
X_5807_ s0.data_out\[21\]\[4\] s0.data_out\[20\]\[4\] net1297 _0392_ VPWR VGND sg13g2_mux2_1
X_5738_ net1301 VPWR _0326_ VGND net1393 net1286 sg13g2_o21ai_1
XFILLER_6_409 VPWR VGND sg13g2_fill_2
X_5669_ _3063_ s0.data_out\[21\]\[6\] net1319 VPWR VGND sg13g2_nand2b_1
X_6512__40 VPWR VGND net40 sg13g2_tiehi
Xfanout996 _2762_ net996 VPWR VGND sg13g2_buf_8
XFILLER_46_869 VPWR VGND sg13g2_decap_8
XFILLER_18_527 VPWR VGND sg13g2_fill_1
XFILLER_18_549 VPWR VGND sg13g2_decap_4
XFILLER_26_571 VPWR VGND sg13g2_decap_4
XFILLER_13_243 VPWR VGND sg13g2_fill_2
XFILLER_14_766 VPWR VGND sg13g2_decap_4
XFILLER_9_203 VPWR VGND sg13g2_decap_8
XFILLER_6_921 VPWR VGND sg13g2_decap_8
XFILLER_10_994 VPWR VGND sg13g2_decap_8
XFILLER_6_998 VPWR VGND sg13g2_decap_8
XFILLER_5_464 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_1_681 VPWR VGND sg13g2_decap_8
XFILLER_23_1001 VPWR VGND sg13g2_decap_8
XFILLER_49_674 VPWR VGND sg13g2_decap_8
XFILLER_48_151 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
X_4971_ _2409_ _2411_ _2434_ VPWR VGND sg13g2_nor2b_1
X_3922_ net1138 net1144 _1488_ VPWR VGND sg13g2_nor2b_1
X_6710_ net122 VGND VPWR _0220_ s0.data_out\[6\]\[4\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_3853_ net1180 net461 _1428_ VPWR VGND sg13g2_and2_1
X_6641_ net196 VGND VPWR net423 s0.data_out\[11\]\[2\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_6572_ net271 VGND VPWR _0082_ s0.data_out\[17\]\[5\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3784_ s0.data_out\[12\]\[3\] s0.data_out\[11\]\[3\] net1187 _1363_ VPWR VGND sg13g2_mux2_1
X_5523_ _2912_ VPWR _2929_ VGND net1449 _2919_ sg13g2_o21ai_1
X_5454_ VPWR _2872_ net676 VGND sg13g2_inv_1
X_5385_ VPWR _2803_ net560 VGND sg13g2_inv_1
X_4405_ VGND VPWR net1097 _1913_ _1916_ _1915_ sg13g2_a21oi_1
X_4336_ VGND VPWR net1114 _1856_ _1859_ _1858_ sg13g2_a21oi_1
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_1017 VPWR VGND sg13g2_decap_8
X_4267_ _1791_ _1792_ _1793_ VPWR VGND sg13g2_nor2_1
X_4198_ _1733_ _1732_ net1405 _1725_ net1414 VPWR VGND sg13g2_a22oi_1
X_6006_ VGND VPWR _0454_ _0566_ _0567_ net1278 sg13g2_a21oi_1
XFILLER_27_302 VPWR VGND sg13g2_fill_1
XFILLER_27_346 VPWR VGND sg13g2_decap_4
XFILLER_27_368 VPWR VGND sg13g2_decap_4
XFILLER_40_44 VPWR VGND sg13g2_decap_8
XFILLER_46_1023 VPWR VGND sg13g2_decap_4
XFILLER_3_957 VPWR VGND sg13g2_decap_8
Xhold280 s0.data_out\[4\]\[0\] VPWR VGND net600 sg13g2_dlygate4sd3_1
XFILLER_49_42 VPWR VGND sg13g2_decap_8
Xhold291 _1543_ VPWR VGND net611 sg13g2_dlygate4sd3_1
XFILLER_18_313 VPWR VGND sg13g2_fill_1
XFILLER_19_869 VPWR VGND sg13g2_decap_8
XFILLER_45_165 VPWR VGND sg13g2_fill_2
X_5170_ VGND VPWR net1005 _2604_ _2609_ _2608_ sg13g2_a21oi_1
X_4121_ VGND VPWR net1130 net675 _1663_ _1623_ sg13g2_a21oi_1
X_4052_ net1441 _1598_ _1599_ VPWR VGND sg13g2_nor2_1
XFILLER_49_471 VPWR VGND sg13g2_fill_1
X_4954_ VGND VPWR _2311_ _2416_ _2417_ net1051 sg13g2_a21oi_1
XFILLER_33_850 VPWR VGND sg13g2_fill_2
XFILLER_20_500 VPWR VGND sg13g2_fill_2
X_3905_ VGND VPWR net1135 _1469_ _1471_ _1470_ sg13g2_a21oi_1
X_4885_ net1066 VPWR _2352_ VGND _2285_ _2351_ sg13g2_o21ai_1
XFILLER_32_382 VPWR VGND sg13g2_decap_4
XFILLER_33_894 VPWR VGND sg13g2_fill_1
X_3836_ _1413_ _1414_ _1415_ VPWR VGND sg13g2_nor2_1
X_6624_ net214 VGND VPWR _0134_ s0.valid_out\[12\][0] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_6555_ net289 VGND VPWR _0065_ s0.data_out\[18\]\[0\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_3767_ _1346_ net1016 _1345_ VPWR VGND sg13g2_nand2_1
X_5506_ VGND VPWR _2912_ _2911_ net1443 sg13g2_or2_1
X_6486_ _0999_ VPWR _1002_ VGND net1229 _1001_ sg13g2_o21ai_1
X_3698_ VGND VPWR _1177_ _1287_ _1288_ net1205 sg13g2_a21oi_1
X_5437_ VPWR _2855_ net555 VGND sg13g2_inv_1
XFILLER_10_58 VPWR VGND sg13g2_fill_2
X_5368_ _2786_ net468 VPWR VGND sg13g2_inv_2
X_4319_ net1102 net1144 _1842_ VPWR VGND sg13g2_nor2b_1
X_5299_ net1465 net386 _2723_ VPWR VGND sg13g2_nor2_1
XFILLER_19_67 VPWR VGND sg13g2_fill_1
XFILLER_28_633 VPWR VGND sg13g2_fill_2
X_6645__192 VPWR VGND net192 sg13g2_tiehi
XFILLER_15_327 VPWR VGND sg13g2_decap_4
XFILLER_30_308 VPWR VGND sg13g2_fill_2
XFILLER_35_77 VPWR VGND sg13g2_decap_8
XFILLER_7_548 VPWR VGND sg13g2_fill_2
XFILLER_13_1022 VPWR VGND sg13g2_decap_8
XFILLER_3_754 VPWR VGND sg13g2_decap_8
XFILLER_47_920 VPWR VGND sg13g2_decap_8
XFILLER_20_1004 VPWR VGND sg13g2_decap_8
XFILLER_19_644 VPWR VGND sg13g2_fill_2
XFILLER_47_997 VPWR VGND sg13g2_decap_8
XFILLER_46_463 VPWR VGND sg13g2_fill_1
XFILLER_19_677 VPWR VGND sg13g2_fill_1
X_4670_ _2156_ VPWR _2157_ VGND net1068 _2866_ sg13g2_o21ai_1
X_3621_ net1218 VPWR _1215_ VGND _1150_ _1214_ sg13g2_o21ai_1
X_6340_ _0871_ VPWR _0872_ VGND net1002 _0870_ sg13g2_o21ai_1
X_3552_ VGND VPWR net1218 _1151_ _1154_ _1153_ sg13g2_a21oi_1
X_3483_ net1018 _2821_ _1092_ VPWR VGND sg13g2_nor2_1
X_6271_ _0808_ net482 net1259 VPWR VGND sg13g2_nand2b_1
X_5222_ net1029 VPWR _2659_ VGND _2592_ _2658_ sg13g2_o21ai_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_5153_ net1020 net1166 _2592_ VPWR VGND sg13g2_nor2b_1
X_4104_ net1135 VPWR _1650_ VGND _1577_ _1649_ sg13g2_o21ai_1
XFILLER_38_942 VPWR VGND sg13g2_decap_8
X_5084_ _2532_ _2534_ net1417 _2535_ VPWR VGND sg13g2_nand3_1
X_4035_ VPWR VGND _1581_ net1459 _1576_ net1455 _1582_ _1574_ sg13g2_a221oi_1
X_6779__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_37_496 VPWR VGND sg13g2_fill_2
X_6599__242 VPWR VGND net242 sg13g2_tiehi
XFILLER_36_1000 VPWR VGND sg13g2_decap_8
X_5986_ net1287 VPWR _0551_ VGND _0488_ _0550_ sg13g2_o21ai_1
X_4937_ VGND VPWR _2283_ _2399_ _2400_ net1051 sg13g2_a21oi_1
X_4868_ net1358 _2279_ _2339_ VPWR VGND sg13g2_nor2_1
X_6607_ net233 VGND VPWR _0117_ s0.data_out\[14\]\[4\] clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_20_374 VPWR VGND sg13g2_fill_2
X_3819_ _1398_ net1015 _1397_ VPWR VGND sg13g2_nand2_1
XFILLER_20_396 VPWR VGND sg13g2_fill_2
X_4799_ _2274_ net1056 net574 VPWR VGND sg13g2_nand2_1
X_6538_ net308 VGND VPWR net474 s0.data_out\[20\]\[7\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_21_79 VPWR VGND sg13g2_fill_2
X_6469_ net1223 s0.data_out\[15\]\[6\] _0987_ VPWR VGND sg13g2_and2_1
XFILLER_43_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_768 VPWR VGND sg13g2_decap_8
XFILLER_48_739 VPWR VGND sg13g2_decap_8
XFILLER_28_463 VPWR VGND sg13g2_fill_2
XFILLER_44_967 VPWR VGND sg13g2_decap_8
XFILLER_15_113 VPWR VGND sg13g2_fill_1
XFILLER_15_135 VPWR VGND sg13g2_fill_2
XFILLER_16_658 VPWR VGND sg13g2_fill_2
XFILLER_11_363 VPWR VGND sg13g2_decap_4
XFILLER_30_7 VPWR VGND sg13g2_fill_1
Xfanout1341 net1343 net1341 VPWR VGND sg13g2_buf_8
Xfanout1330 net1333 net1330 VPWR VGND sg13g2_buf_8
Xfanout1363 net1364 net1363 VPWR VGND sg13g2_buf_8
Xfanout1352 net1354 net1352 VPWR VGND sg13g2_buf_8
Xfanout1374 net1376 net1374 VPWR VGND sg13g2_buf_8
Xfanout1396 net1397 net1396 VPWR VGND sg13g2_buf_8
XFILLER_4_1020 VPWR VGND sg13g2_decap_8
Xfanout1385 net1388 net1385 VPWR VGND sg13g2_buf_8
XFILLER_47_794 VPWR VGND sg13g2_decap_8
XFILLER_35_967 VPWR VGND sg13g2_decap_8
X_5840_ _0030_ _0421_ _0422_ _2782_ net1345 VPWR VGND sg13g2_a22oi_1
X_5771_ _0355_ VPWR _0356_ VGND net1007 _0353_ sg13g2_o21ai_1
X_4722_ _2186_ _2208_ _2209_ VPWR VGND sg13g2_nor2b_1
X_4653_ VGND VPWR net1072 _2137_ _2140_ _2139_ sg13g2_a21oi_1
X_4584_ VGND VPWR net1078 _2081_ _2083_ _2082_ sg13g2_a21oi_1
X_3604_ net1378 _1144_ _1202_ VPWR VGND sg13g2_nor2_1
X_3535_ VPWR VGND _1136_ net1459 _1134_ net1454 _1137_ _1130_ sg13g2_a221oi_1
X_6323_ _0801_ _0858_ net1478 _0859_ VPWR VGND sg13g2_nand3_1
X_6254_ _0790_ VPWR _0791_ VGND net1246 _2807_ sg13g2_o21ai_1
X_3466_ net1213 s0.data_out\[14\]\[0\] _1079_ VPWR VGND sg13g2_and2_1
X_5205_ _2630_ _2635_ net1426 _2644_ VPWR VGND sg13g2_nand3_1
X_6185_ VGND VPWR _0620_ _0733_ _0734_ net1263 sg13g2_a21oi_1
X_3397_ VGND VPWR _1011_ _1010_ net1445 sg13g2_or2_1
X_5136_ VGND VPWR _2578_ net1026 net427 sg13g2_or2_1
X_5067_ _2518_ _2517_ net1408 _2511_ net1399 VPWR VGND sg13g2_a22oi_1
XFILLER_29_249 VPWR VGND sg13g2_decap_4
X_4018_ net1151 net1416 net1390 _0164_ VPWR VGND sg13g2_mux2_1
XFILLER_26_923 VPWR VGND sg13g2_fill_2
XFILLER_25_422 VPWR VGND sg13g2_decap_8
XFILLER_26_978 VPWR VGND sg13g2_decap_8
X_6642__195 VPWR VGND net195 sg13g2_tiehi
XFILLER_41_959 VPWR VGND sg13g2_decap_8
XFILLER_12_116 VPWR VGND sg13g2_fill_2
XFILLER_13_628 VPWR VGND sg13g2_fill_1
X_5969_ _2755_ _2794_ _0538_ VPWR VGND sg13g2_nor2_1
XFILLER_21_650 VPWR VGND sg13g2_decap_8
XFILLER_21_683 VPWR VGND sg13g2_fill_1
XFILLER_20_171 VPWR VGND sg13g2_fill_2
XFILLER_5_827 VPWR VGND sg13g2_decap_8
XFILLER_0_565 VPWR VGND sg13g2_decap_8
XFILLER_48_569 VPWR VGND sg13g2_fill_2
XFILLER_16_444 VPWR VGND sg13g2_fill_2
XFILLER_17_978 VPWR VGND sg13g2_decap_8
XFILLER_31_469 VPWR VGND sg13g2_fill_1
XFILLER_40_981 VPWR VGND sg13g2_decap_8
XFILLER_8_632 VPWR VGND sg13g2_decap_4
XFILLER_8_698 VPWR VGND sg13g2_fill_1
XFILLER_7_142 VPWR VGND sg13g2_decap_8
Xhold109 _0067_ VPWR VGND net429 sg13g2_dlygate4sd3_1
X_6589__252 VPWR VGND net252 sg13g2_tiehi
Xfanout1160 net704 net1160 VPWR VGND sg13g2_buf_8
Xfanout1171 net1172 net1171 VPWR VGND sg13g2_buf_8
Xfanout1182 net1183 net1182 VPWR VGND sg13g2_buf_8
Xfanout1193 net391 net1193 VPWR VGND sg13g2_buf_8
XFILLER_26_219 VPWR VGND sg13g2_fill_2
XFILLER_34_241 VPWR VGND sg13g2_fill_2
X_5823_ VGND VPWR _0402_ _0404_ _0408_ net1418 sg13g2_a21oi_1
X_6596__245 VPWR VGND net245 sg13g2_tiehi
X_5754_ _0337_ net1290 _0338_ _0339_ VPWR VGND sg13g2_a21o_1
XFILLER_33_1014 VPWR VGND sg13g2_decap_8
X_5685_ s0.data_out\[22\]\[5\] s0.data_out\[21\]\[5\] net1307 _3079_ VPWR VGND sg13g2_mux2_1
XFILLER_31_992 VPWR VGND sg13g2_decap_8
X_4705_ s0.data_out\[4\]\[4\] s0.data_out\[5\]\[4\] net1080 _2192_ VPWR VGND sg13g2_mux2_1
X_4636_ VGND VPWR net1336 net1070 _2126_ _2125_ sg13g2_a21oi_1
X_4567_ _2064_ net1079 _2065_ _2066_ VPWR VGND sg13g2_a21o_1
X_6306_ s0.data_out\[17\]\[4\] s0.data_out\[16\]\[4\] net1245 _0843_ VPWR VGND sg13g2_mux2_1
XFILLER_2_819 VPWR VGND sg13g2_decap_8
X_4498_ net1101 VPWR _2003_ VGND _1961_ _2002_ sg13g2_o21ai_1
X_3518_ _1120_ net457 net1220 VPWR VGND sg13g2_nand2b_1
X_6237_ net1236 _0773_ _0777_ VPWR VGND sg13g2_nor2_1
X_3449_ _1063_ net1221 s0.data_out\[14\]\[4\] VPWR VGND sg13g2_nand2_1
X_6168_ VGND VPWR net1262 _0714_ _0717_ _0716_ sg13g2_a21oi_1
X_5119_ VGND VPWR net1030 s0.data_out\[1\]\[5\] _2564_ _2530_ sg13g2_a21oi_1
X_6099_ net1353 _0625_ _0654_ VPWR VGND sg13g2_nor2_1
XFILLER_26_720 VPWR VGND sg13g2_fill_2
XFILLER_26_775 VPWR VGND sg13g2_decap_4
XFILLER_40_211 VPWR VGND sg13g2_fill_2
XFILLER_13_403 VPWR VGND sg13g2_fill_1
XFILLER_25_263 VPWR VGND sg13g2_decap_4
XFILLER_40_277 VPWR VGND sg13g2_fill_2
XFILLER_13_469 VPWR VGND sg13g2_decap_8
XFILLER_49_1010 VPWR VGND sg13g2_decap_8
XFILLER_1_863 VPWR VGND sg13g2_decap_8
XFILLER_0_362 VPWR VGND sg13g2_fill_1
XFILLER_49_856 VPWR VGND sg13g2_decap_8
XFILLER_32_745 VPWR VGND sg13g2_fill_2
X_6739__90 VPWR VGND net90 sg13g2_tiehi
XFILLER_31_299 VPWR VGND sg13g2_fill_1
XFILLER_8_451 VPWR VGND sg13g2_decap_4
XFILLER_9_996 VPWR VGND sg13g2_decap_8
X_5470_ _2887_ net1449 _2885_ VPWR VGND sg13g2_nand2_1
X_4421_ VPWR VGND _1930_ net1460 _1928_ net1453 _1932_ _1924_ sg13g2_a221oi_1
X_4352_ net324 net1331 _1874_ _0191_ VPWR VGND sg13g2_nor3_1
X_6521__30 VPWR VGND net30 sg13g2_tiehi
XFILLER_4_690 VPWR VGND sg13g2_decap_8
X_4283_ VGND VPWR net1110 _1803_ _1806_ _1805_ sg13g2_a21oi_1
X_6022_ VPWR VGND _0582_ net1460 _0580_ net1452 _0583_ _0576_ sg13g2_a221oi_1
XFILLER_39_399 VPWR VGND sg13g2_decap_8
XFILLER_27_539 VPWR VGND sg13g2_decap_8
X_3998_ _0156_ _1554_ _1555_ _2834_ net1387 VPWR VGND sg13g2_a22oi_1
X_5806_ _0391_ net1298 net496 VPWR VGND sg13g2_nand2_1
XFILLER_11_918 VPWR VGND sg13g2_decap_8
X_5737_ _0024_ net528 _0325_ _2763_ net1340 VPWR VGND sg13g2_a22oi_1
XFILLER_10_428 VPWR VGND sg13g2_fill_1
X_5668_ _3060_ net1300 _3061_ _3062_ VPWR VGND sg13g2_a21o_1
X_4619_ _2112_ VPWR _2113_ VGND net998 _2111_ sg13g2_o21ai_1
X_5599_ _0009_ _2998_ _2999_ _2769_ net1339 VPWR VGND sg13g2_a22oi_1
XFILLER_2_627 VPWR VGND sg13g2_decap_4
XFILLER_49_119 VPWR VGND sg13g2_fill_1
XFILLER_38_88 VPWR VGND sg13g2_decap_4
Xfanout997 net998 net997 VPWR VGND sg13g2_buf_8
XFILLER_46_848 VPWR VGND sg13g2_decap_8
XFILLER_14_734 VPWR VGND sg13g2_fill_1
XFILLER_14_778 VPWR VGND sg13g2_fill_1
XFILLER_13_288 VPWR VGND sg13g2_fill_2
XFILLER_13_299 VPWR VGND sg13g2_decap_4
XFILLER_6_900 VPWR VGND sg13g2_decap_8
XFILLER_10_973 VPWR VGND sg13g2_decap_8
XFILLER_6_977 VPWR VGND sg13g2_decap_8
XFILLER_1_660 VPWR VGND sg13g2_decap_8
XFILLER_0_181 VPWR VGND sg13g2_fill_2
XFILLER_0_170 VPWR VGND sg13g2_decap_8
XFILLER_49_653 VPWR VGND sg13g2_decap_8
X_4970_ _2412_ _2432_ _2433_ VPWR VGND sg13g2_nor2b_1
X_3921_ s0.data_out\[11\]\[7\] s0.data_out\[10\]\[7\] net1175 _1487_ VPWR VGND sg13g2_mux2_1
X_6640_ net197 VGND VPWR _0150_ s0.data_out\[11\]\[1\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_3852_ VPWR _0138_ _1427_ VGND sg13g2_inv_1
X_6593__248 VPWR VGND net248 sg13g2_tiehi
X_6571_ net272 VGND VPWR _0081_ s0.data_out\[17\]\[4\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_20_748 VPWR VGND sg13g2_decap_8
X_5522_ net1458 _2927_ _2928_ VPWR VGND sg13g2_nor2_1
XFILLER_30_1017 VPWR VGND sg13g2_decap_8
X_3783_ _1362_ net1187 net461 VPWR VGND sg13g2_nand2_1
XFILLER_9_793 VPWR VGND sg13g2_decap_4
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
X_5453_ VPWR _2871_ net444 VGND sg13g2_inv_1
X_5384_ VPWR _2802_ net418 VGND sg13g2_inv_1
X_4404_ VGND VPWR _1800_ _1914_ _1915_ net1096 sg13g2_a21oi_1
X_6710__122 VPWR VGND net122 sg13g2_tiehi
X_4335_ VGND VPWR _1737_ _1857_ _1858_ net1114 sg13g2_a21oi_1
X_4266_ net1394 _2760_ _1792_ VPWR VGND sg13g2_nor2_1
X_4197_ VGND VPWR net1126 _1729_ _1732_ _1731_ sg13g2_a21oi_1
X_6005_ _0566_ net428 net1283 VPWR VGND sg13g2_nand2b_1
XFILLER_42_306 VPWR VGND sg13g2_fill_1
XFILLER_11_704 VPWR VGND sg13g2_fill_2
XFILLER_24_57 VPWR VGND sg13g2_decap_8
XFILLER_11_737 VPWR VGND sg13g2_fill_1
XFILLER_11_748 VPWR VGND sg13g2_fill_1
XFILLER_10_247 VPWR VGND sg13g2_decap_8
X_6769_ net293 VGND VPWR _0279_ s0.data_out\[1\]\[3\] clknet_leaf_9_clk sg13g2_dfrbpq_2
XFILLER_40_78 VPWR VGND sg13g2_decap_4
XFILLER_3_936 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_46_1002 VPWR VGND sg13g2_decap_8
Xhold270 _0183_ VPWR VGND net590 sg13g2_dlygate4sd3_1
Xhold281 s0.data_out\[3\]\[5\] VPWR VGND net601 sg13g2_dlygate4sd3_1
Xhold292 s0.data_out\[14\]\[7\] VPWR VGND net612 sg13g2_dlygate4sd3_1
XFILLER_49_87 VPWR VGND sg13g2_decap_8
XFILLER_19_837 VPWR VGND sg13g2_fill_1
XFILLER_18_358 VPWR VGND sg13g2_fill_1
XFILLER_46_689 VPWR VGND sg13g2_decap_4
XFILLER_14_531 VPWR VGND sg13g2_decap_8
XFILLER_26_391 VPWR VGND sg13g2_decap_4
XFILLER_6_763 VPWR VGND sg13g2_fill_2
XFILLER_2_980 VPWR VGND sg13g2_decap_8
X_4120_ _0171_ _1661_ _1662_ _2840_ net1388 VPWR VGND sg13g2_a22oi_1
X_4051_ VGND VPWR net1137 _1595_ _1598_ _1597_ sg13g2_a21oi_1
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_49_483 VPWR VGND sg13g2_decap_8
XFILLER_24_317 VPWR VGND sg13g2_fill_1
X_4953_ _2416_ net576 net1058 VPWR VGND sg13g2_nand2b_1
XFILLER_36_199 VPWR VGND sg13g2_decap_8
X_3904_ net1135 net1171 _1470_ VPWR VGND sg13g2_nor2b_1
X_4884_ net1053 net484 _2351_ VPWR VGND sg13g2_and2_1
X_6623_ net216 VGND VPWR net349 s0.was_valid_out\[12\][0] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_3835_ _1332_ VPWR _1414_ VGND _1388_ _1390_ sg13g2_o21ai_1
X_6554_ net290 VGND VPWR _0064_ s0.shift_out\[18\][0] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3766_ s0.data_out\[11\]\[0\] s0.data_out\[12\]\[0\] net1197 _1345_ VPWR VGND sg13g2_mux2_1
X_6485_ s0.was_valid_out\[14\][0] net1234 _1001_ VPWR VGND sg13g2_nor2_1
X_5505_ VGND VPWR net1325 _2910_ _2911_ _2907_ sg13g2_a21oi_1
X_3697_ _1287_ net414 net1211 VPWR VGND sg13g2_nand2b_1
X_5436_ _2854_ net537 VPWR VGND sg13g2_inv_2
X_5367_ VPWR _2785_ net432 VGND sg13g2_inv_1
X_4318_ s0.data_out\[8\]\[7\] s0.data_out\[7\]\[7\] net1108 _1841_ VPWR VGND sg13g2_mux2_1
X_5298_ VGND VPWR net1464 _2691_ _0289_ _2722_ sg13g2_a21oi_1
X_4249_ _1752_ _1778_ net1488 _1779_ VPWR VGND sg13g2_nand3_1
XFILLER_16_807 VPWR VGND sg13g2_fill_1
XFILLER_27_144 VPWR VGND sg13g2_fill_1
XFILLER_43_604 VPWR VGND sg13g2_decap_8
XFILLER_15_317 VPWR VGND sg13g2_fill_2
XFILLER_43_659 VPWR VGND sg13g2_fill_1
XFILLER_13_1001 VPWR VGND sg13g2_decap_8
XFILLER_3_733 VPWR VGND sg13g2_decap_8
XFILLER_2_232 VPWR VGND sg13g2_fill_2
XFILLER_47_976 VPWR VGND sg13g2_decap_8
XFILLER_46_442 VPWR VGND sg13g2_fill_1
XFILLER_18_144 VPWR VGND sg13g2_decap_4
XFILLER_18_166 VPWR VGND sg13g2_fill_2
XFILLER_15_873 VPWR VGND sg13g2_fill_1
XFILLER_30_843 VPWR VGND sg13g2_fill_1
X_3620_ net1206 net406 _1214_ VPWR VGND sg13g2_and2_1
X_3551_ VGND VPWR _1036_ _1152_ _1153_ net1218 sg13g2_a21oi_1
X_3482_ _0104_ _1090_ _1091_ _2816_ net1367 VPWR VGND sg13g2_a22oi_1
X_6270_ _0805_ net1239 _0806_ _0807_ VPWR VGND sg13g2_a21o_1
X_5221_ net1020 net375 _2658_ VPWR VGND sg13g2_and2_1
X_5152_ s0.data_out\[1\]\[1\] s0.data_out\[0\]\[1\] net1026 _2591_ VPWR VGND sg13g2_mux2_1
XFILLER_29_409 VPWR VGND sg13g2_fill_1
X_4103_ net1123 s0.data_out\[9\]\[0\] _1649_ VPWR VGND sg13g2_and2_1
X_5083_ _2534_ _2751_ _2533_ VPWR VGND sg13g2_nand2_1
XFILLER_49_291 VPWR VGND sg13g2_fill_2
X_4034_ _1581_ net1135 _1580_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_998 VPWR VGND sg13g2_decap_8
X_5985_ net1003 _2791_ _0550_ VPWR VGND sg13g2_nor2_1
XFILLER_24_147 VPWR VGND sg13g2_decap_4
X_4936_ _2399_ s0.data_out\[2\]\[7\] net1058 VPWR VGND sg13g2_nand2b_1
XFILLER_32_180 VPWR VGND sg13g2_decap_8
X_4867_ net1063 VPWR _2338_ VGND _2276_ _2337_ sg13g2_o21ai_1
X_6606_ net234 VGND VPWR _0116_ s0.data_out\[14\]\[3\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_20_353 VPWR VGND sg13g2_fill_2
X_3818_ _1283_ VPWR _1397_ VGND net1198 _2835_ sg13g2_o21ai_1
X_6537_ net309 VGND VPWR net433 s0.data_out\[20\]\[6\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_4798_ _2258_ VPWR _2273_ VGND net1451 _2265_ sg13g2_o21ai_1
X_3749_ net1395 _2745_ _1330_ VPWR VGND sg13g2_nor2_1
X_6468_ _0094_ _0985_ _0986_ _2809_ net1368 VPWR VGND sg13g2_a22oi_1
X_6399_ _0923_ VPWR _0924_ VGND _0914_ _0915_ sg13g2_o21ai_1
X_5419_ VPWR _2837_ net422 VGND sg13g2_inv_1
XFILLER_43_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_747 VPWR VGND sg13g2_decap_8
XFILLER_48_718 VPWR VGND sg13g2_decap_8
XFILLER_29_987 VPWR VGND sg13g2_decap_8
XFILLER_44_946 VPWR VGND sg13g2_decap_8
XFILLER_43_445 VPWR VGND sg13g2_fill_2
XFILLER_12_865 VPWR VGND sg13g2_fill_1
XFILLER_8_836 VPWR VGND sg13g2_decap_4
XFILLER_7_16 VPWR VGND sg13g2_decap_4
XFILLER_7_335 VPWR VGND sg13g2_fill_1
XFILLER_7_38 VPWR VGND sg13g2_fill_1
XFILLER_11_91 VPWR VGND sg13g2_decap_8
XFILLER_39_707 VPWR VGND sg13g2_fill_2
Xfanout1320 net1322 net1320 VPWR VGND sg13g2_buf_8
Xfanout1331 net1333 net1331 VPWR VGND sg13g2_buf_8
Xfanout1375 net1376 net1375 VPWR VGND sg13g2_buf_8
Xfanout1353 net1354 net1353 VPWR VGND sg13g2_buf_1
Xfanout1342 net1343 net1342 VPWR VGND sg13g2_buf_1
Xfanout1364 net1389 net1364 VPWR VGND sg13g2_buf_8
Xfanout1397 uio_in[0] net1397 VPWR VGND sg13g2_buf_8
Xfanout1386 net1388 net1386 VPWR VGND sg13g2_buf_8
XFILLER_47_773 VPWR VGND sg13g2_decap_8
XFILLER_34_467 VPWR VGND sg13g2_fill_2
X_5770_ _0355_ net1007 _0354_ VPWR VGND sg13g2_nand2_1
XFILLER_22_629 VPWR VGND sg13g2_fill_1
X_4721_ _2202_ VPWR _2208_ VGND _2194_ _2205_ sg13g2_o21ai_1
X_4652_ VGND VPWR _2020_ _2138_ _2139_ net1072 sg13g2_a21oi_1
X_3603_ net1216 VPWR _1201_ VGND _1141_ _1200_ sg13g2_o21ai_1
X_4583_ net1078 net1153 _2082_ VPWR VGND sg13g2_nor2b_1
X_6322_ net1255 VPWR _0858_ VGND _0797_ _0857_ sg13g2_o21ai_1
X_3534_ _1136_ net1018 _1135_ VPWR VGND sg13g2_nand2_1
X_3465_ net323 net1332 _1078_ _0100_ VPWR VGND sg13g2_nor3_1
X_6253_ _0790_ net1245 net479 VPWR VGND sg13g2_nand2_1
X_5204_ _2638_ _2642_ net1417 _2643_ VPWR VGND sg13g2_nand3_1
X_6184_ _0733_ net368 net1269 VPWR VGND sg13g2_nand2b_1
X_3396_ VGND VPWR net1227 _1007_ _1010_ _1009_ sg13g2_a21oi_1
X_5135_ _2576_ VPWR _2577_ VGND net1031 _2464_ sg13g2_o21ai_1
XFILLER_29_206 VPWR VGND sg13g2_fill_2
X_5066_ VGND VPWR net1039 _2514_ _2517_ _2516_ sg13g2_a21oi_1
XFILLER_38_773 VPWR VGND sg13g2_fill_2
XFILLER_38_762 VPWR VGND sg13g2_decap_8
X_4017_ VGND VPWR net1390 _2768_ _0163_ _1567_ sg13g2_a21oi_1
XFILLER_37_272 VPWR VGND sg13g2_fill_1
XFILLER_26_957 VPWR VGND sg13g2_decap_8
XFILLER_13_607 VPWR VGND sg13g2_decap_4
XFILLER_41_938 VPWR VGND sg13g2_decap_8
X_5968_ _0043_ _0536_ _0537_ _2789_ net1354 VPWR VGND sg13g2_a22oi_1
X_4919_ s0.data_out\[2\]\[0\] s0.data_out\[3\]\[0\] net1056 _2382_ VPWR VGND sg13g2_mux2_1
X_5899_ _0472_ net1293 _0471_ VPWR VGND sg13g2_nand2b_1
XFILLER_20_183 VPWR VGND sg13g2_fill_1
XFILLER_4_316 VPWR VGND sg13g2_fill_2
XFILLER_10_1015 VPWR VGND sg13g2_decap_8
XFILLER_20_194 VPWR VGND sg13g2_decap_8
XFILLER_0_544 VPWR VGND sg13g2_decap_8
XFILLER_29_762 VPWR VGND sg13g2_fill_1
XFILLER_44_721 VPWR VGND sg13g2_fill_2
XFILLER_28_272 VPWR VGND sg13g2_fill_1
XFILLER_44_776 VPWR VGND sg13g2_decap_8
XFILLER_44_787 VPWR VGND sg13g2_fill_1
XFILLER_43_264 VPWR VGND sg13g2_fill_2
XFILLER_31_404 VPWR VGND sg13g2_fill_1
XFILLER_32_927 VPWR VGND sg13g2_fill_2
XFILLER_40_960 VPWR VGND sg13g2_decap_8
XFILLER_12_673 VPWR VGND sg13g2_decap_8
XFILLER_11_172 VPWR VGND sg13g2_fill_1
XFILLER_11_183 VPWR VGND sg13g2_fill_2
XFILLER_7_198 VPWR VGND sg13g2_fill_1
XFILLER_7_187 VPWR VGND sg13g2_fill_2
XFILLER_4_894 VPWR VGND sg13g2_decap_8
Xfanout1150 net709 net1150 VPWR VGND sg13g2_buf_8
XFILLER_39_548 VPWR VGND sg13g2_decap_4
Xfanout1172 net1173 net1172 VPWR VGND sg13g2_buf_8
Xfanout1183 net1186 net1183 VPWR VGND sg13g2_buf_8
Xfanout1161 s0.data_new_delayed\[3\] net1161 VPWR VGND sg13g2_buf_8
Xfanout1194 net391 net1194 VPWR VGND sg13g2_buf_2
XFILLER_35_743 VPWR VGND sg13g2_decap_8
X_5822_ VGND VPWR _0394_ _0396_ _0407_ net1427 sg13g2_a21oi_1
X_5753_ net1290 net1166 _0338_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_297 VPWR VGND sg13g2_fill_2
X_4704_ _2191_ net1073 _2190_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_971 VPWR VGND sg13g2_decap_8
X_5684_ _3078_ net1308 s0.data_out\[21\]\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_30_492 VPWR VGND sg13g2_decap_4
X_4635_ net1076 VPWR _2125_ VGND net1393 net1065 sg13g2_o21ai_1
X_4566_ net1078 net1148 _2065_ VPWR VGND sg13g2_nor2b_1
X_6305_ _0842_ net1247 net525 VPWR VGND sg13g2_nand2_1
X_3517_ _1117_ net1203 _1118_ _1119_ VPWR VGND sg13g2_a21o_1
X_4497_ net1090 s0.data_out\[6\]\[5\] _2002_ VPWR VGND sg13g2_and2_1
X_6236_ _0774_ VPWR _0776_ VGND net370 net1245 sg13g2_o21ai_1
X_3448_ net1423 _1061_ _1062_ VPWR VGND sg13g2_nor2_1
X_6167_ VGND VPWR _0601_ _0715_ _0716_ net1262 sg13g2_a21oi_1
X_5118_ VPWR _0268_ net584 VGND sg13g2_inv_1
X_6098_ net1275 VPWR _0653_ VGND _0622_ _0652_ sg13g2_o21ai_1
XFILLER_17_209 VPWR VGND sg13g2_decap_4
X_5049_ net1435 _2499_ _2500_ VPWR VGND sg13g2_nor2_1
XFILLER_27_79 VPWR VGND sg13g2_decap_4
XFILLER_13_448 VPWR VGND sg13g2_decap_8
XFILLER_40_289 VPWR VGND sg13g2_fill_2
XFILLER_5_603 VPWR VGND sg13g2_fill_1
X_6770__280 VPWR VGND net280 sg13g2_tiehi
XFILLER_0_330 VPWR VGND sg13g2_decap_8
XFILLER_1_842 VPWR VGND sg13g2_decap_8
XFILLER_49_835 VPWR VGND sg13g2_decap_8
XFILLER_36_529 VPWR VGND sg13g2_decap_8
XFILLER_1_1024 VPWR VGND sg13g2_decap_4
XFILLER_17_721 VPWR VGND sg13g2_decap_8
XFILLER_17_743 VPWR VGND sg13g2_fill_2
XFILLER_17_754 VPWR VGND sg13g2_fill_2
XFILLER_32_724 VPWR VGND sg13g2_fill_2
XFILLER_40_790 VPWR VGND sg13g2_decap_4
XFILLER_9_975 VPWR VGND sg13g2_decap_8
XFILLER_8_496 VPWR VGND sg13g2_fill_1
X_4420_ net1453 _1924_ _1931_ VPWR VGND sg13g2_nor2_1
X_4351_ VPWR VGND _1851_ _1873_ _1872_ _1832_ _1874_ _1871_ sg13g2_a221oi_1
X_4282_ VGND VPWR _1687_ _1804_ _1805_ net1110 sg13g2_a21oi_1
X_6021_ _0582_ net1003 _0581_ VPWR VGND sg13g2_nand2_1
X_6785_ net65 VGND VPWR _0295_ s0.data_out\[0\]\[7\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_3997_ net1387 _1491_ _1555_ VPWR VGND sg13g2_nor2_1
X_5805_ net1292 net1157 _0390_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_779 VPWR VGND sg13g2_fill_2
X_5736_ net1343 net378 _0325_ VPWR VGND sg13g2_nor2_1
XFILLER_10_418 VPWR VGND sg13g2_fill_2
X_5667_ net1300 net1147 _3061_ VPWR VGND sg13g2_nor2b_1
X_4618_ VGND VPWR net998 _2078_ _2112_ net1370 sg13g2_a21oi_1
X_5598_ net1339 _2962_ _2999_ VPWR VGND sg13g2_nor2_1
X_4549_ _2048_ net997 _2047_ VPWR VGND sg13g2_nand2_1
X_6219_ _0069_ _0761_ _0762_ _2799_ net1356 VPWR VGND sg13g2_a22oi_1
Xfanout998 _2761_ net998 VPWR VGND sg13g2_buf_8
XFILLER_18_507 VPWR VGND sg13g2_fill_1
XFILLER_46_827 VPWR VGND sg13g2_decap_8
XFILLER_18_518 VPWR VGND sg13g2_decap_8
X_6579__263 VPWR VGND net263 sg13g2_tiehi
X_6736__94 VPWR VGND net94 sg13g2_tiehi
XFILLER_10_952 VPWR VGND sg13g2_decap_8
XFILLER_6_956 VPWR VGND sg13g2_decap_8
XFILLER_49_632 VPWR VGND sg13g2_decap_8
X_6586__256 VPWR VGND net256 sg13g2_tiehi
XFILLER_36_348 VPWR VGND sg13g2_fill_2
X_3920_ _1486_ net1175 net536 VPWR VGND sg13g2_nand2_1
XFILLER_45_893 VPWR VGND sg13g2_decap_8
X_3851_ _1426_ VPWR _1427_ VGND net1488 net651 sg13g2_o21ai_1
XFILLER_32_543 VPWR VGND sg13g2_decap_4
X_6570_ net273 VGND VPWR _0080_ s0.data_out\[17\]\[3\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3782_ net1455 _1344_ _1361_ VPWR VGND sg13g2_nor2_1
XFILLER_32_598 VPWR VGND sg13g2_fill_2
X_5521_ VGND VPWR net1325 _2926_ _2927_ _2922_ sg13g2_a21oi_1
X_5452_ VPWR _2870_ net507 VGND sg13g2_inv_1
X_5383_ VPWR _2801_ net428 VGND sg13g2_inv_1
X_4403_ _1914_ s0.data_out\[6\]\[2\] net1105 VPWR VGND sg13g2_nand2b_1
X_4334_ _1857_ net470 net1120 VPWR VGND sg13g2_nand2b_1
XFILLER_5_71 VPWR VGND sg13g2_fill_1
X_4265_ net1114 VPWR _1791_ VGND net1394 net1103 sg13g2_o21ai_1
X_6004_ _0563_ net1265 _0564_ _0565_ VPWR VGND sg13g2_a21o_1
X_4196_ VGND VPWR _1605_ _1730_ _1731_ net1126 sg13g2_a21oi_1
XFILLER_39_1010 VPWR VGND sg13g2_decap_8
XFILLER_24_47 VPWR VGND sg13g2_fill_1
XFILLER_10_204 VPWR VGND sg13g2_fill_2
X_6768_ net306 VGND VPWR _0278_ s0.data_out\[1\]\[2\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_6699_ net134 VGND VPWR net471 s0.data_out\[7\]\[5\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_5719_ _0020_ _0310_ _0311_ _2770_ net1342 VPWR VGND sg13g2_a22oi_1
XFILLER_3_915 VPWR VGND sg13g2_decap_8
X_6733__97 VPWR VGND net97 sg13g2_tiehi
Xhold260 s0.data_out\[2\]\[6\] VPWR VGND net580 sg13g2_dlygate4sd3_1
Xhold271 s0.data_out\[14\]\[0\] VPWR VGND net591 sg13g2_dlygate4sd3_1
Xhold293 s0.data_out\[10\]\[5\] VPWR VGND net613 sg13g2_dlygate4sd3_1
XFILLER_2_458 VPWR VGND sg13g2_fill_2
XFILLER_2_469 VPWR VGND sg13g2_fill_2
Xhold282 s0.data_out\[14\]\[3\] VPWR VGND net602 sg13g2_dlygate4sd3_1
XFILLER_18_304 VPWR VGND sg13g2_decap_8
XFILLER_46_646 VPWR VGND sg13g2_fill_1
XFILLER_42_830 VPWR VGND sg13g2_fill_2
X_4050_ VGND VPWR _1477_ _1596_ _1597_ net1137 sg13g2_a21oi_1
XFILLER_37_657 VPWR VGND sg13g2_fill_2
X_4952_ _2413_ net1040 _2414_ _2415_ VPWR VGND sg13g2_a21o_1
X_4883_ _0246_ _2349_ _2350_ _2870_ net1360 VPWR VGND sg13g2_a22oi_1
X_3903_ s0.data_out\[11\]\[0\] s0.data_out\[10\]\[0\] net1174 _1469_ VPWR VGND sg13g2_mux2_1
XFILLER_33_852 VPWR VGND sg13g2_fill_1
X_6622_ net217 VGND VPWR net407 s0.data_out\[13\]\[7\] clknet_leaf_28_clk sg13g2_dfrbpq_2
XFILLER_20_502 VPWR VGND sg13g2_fill_1
XFILLER_20_513 VPWR VGND sg13g2_fill_2
X_3834_ _1391_ _1412_ _1413_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_535 VPWR VGND sg13g2_decap_4
XFILLER_32_395 VPWR VGND sg13g2_fill_1
X_6553_ net291 VGND VPWR _0063_ s0.genblk1\[17\].modules.bubble clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_3765_ VGND VPWR net1192 _1341_ _1344_ _1343_ sg13g2_a21oi_1
X_6484_ net1217 _0994_ _1000_ VPWR VGND sg13g2_nor2_1
X_3696_ _1284_ net1196 _1285_ _1286_ VPWR VGND sg13g2_a21o_1
X_5504_ _2908_ net1315 _2909_ _2910_ VPWR VGND sg13g2_a21o_1
XFILLER_10_16 VPWR VGND sg13g2_decap_4
X_5435_ VPWR _2853_ net673 VGND sg13g2_inv_1
X_5366_ VPWR _2784_ net473 VGND sg13g2_inv_1
XFILLER_0_929 VPWR VGND sg13g2_decap_8
X_4317_ _1840_ net1107 net555 VPWR VGND sg13g2_nand2_1
X_5297_ net1464 net375 _2722_ VPWR VGND sg13g2_nor2_1
X_4248_ net1125 VPWR _1778_ VGND _1748_ _1777_ sg13g2_o21ai_1
XFILLER_28_602 VPWR VGND sg13g2_fill_2
X_4179_ _1714_ _2747_ s0.data_out\[8\]\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_28_657 VPWR VGND sg13g2_fill_2
XFILLER_28_679 VPWR VGND sg13g2_decap_8
XFILLER_27_178 VPWR VGND sg13g2_fill_1
XFILLER_24_863 VPWR VGND sg13g2_decap_8
XFILLER_24_874 VPWR VGND sg13g2_fill_2
XFILLER_24_896 VPWR VGND sg13g2_decap_4
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
X_6576__266 VPWR VGND net266 sg13g2_tiehi
XFILLER_11_579 VPWR VGND sg13g2_decap_8
XFILLER_3_712 VPWR VGND sg13g2_decap_8
XFILLER_3_789 VPWR VGND sg13g2_decap_8
X_6583__259 VPWR VGND net259 sg13g2_tiehi
XFILLER_47_955 VPWR VGND sg13g2_decap_8
XFILLER_19_657 VPWR VGND sg13g2_decap_8
XFILLER_34_605 VPWR VGND sg13g2_fill_2
X_6700__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_15_885 VPWR VGND sg13g2_decap_4
XFILLER_15_896 VPWR VGND sg13g2_fill_1
XFILLER_30_822 VPWR VGND sg13g2_decap_4
X_3550_ _1152_ net406 net1222 VPWR VGND sg13g2_nand2b_1
XFILLER_6_594 VPWR VGND sg13g2_fill_1
XFILLER_6_583 VPWR VGND sg13g2_decap_8
X_3481_ net1367 _1032_ _1091_ VPWR VGND sg13g2_nor2_1
X_5220_ VPWR _0276_ _2657_ VGND sg13g2_inv_1
X_5151_ VGND VPWR _2472_ _2589_ _2590_ net1029 sg13g2_a21oi_1
X_4102_ VGND VPWR _1643_ _1647_ _0167_ _1648_ sg13g2_a21oi_1
X_5082_ s0.data_out\[1\]\[5\] s0.data_out\[2\]\[5\] net1045 _2533_ VPWR VGND sg13g2_mux2_1
XFILLER_38_922 VPWR VGND sg13g2_decap_8
X_4033_ VGND VPWR net1124 _1579_ _1580_ _1577_ sg13g2_a21oi_1
XFILLER_38_977 VPWR VGND sg13g2_decap_8
XFILLER_37_476 VPWR VGND sg13g2_decap_8
XFILLER_25_627 VPWR VGND sg13g2_decap_4
X_5984_ _0047_ _0548_ _0549_ _2785_ net1352 VPWR VGND sg13g2_a22oi_1
X_4935_ _2396_ net1040 _2397_ _2398_ VPWR VGND sg13g2_a21o_1
XFILLER_21_866 VPWR VGND sg13g2_decap_8
X_4866_ net1050 s0.data_out\[3\]\[3\] _2337_ VPWR VGND sg13g2_and2_1
X_6605_ net235 VGND VPWR _0115_ s0.data_out\[14\]\[2\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_3817_ _1396_ net1196 _1395_ VPWR VGND sg13g2_nand2b_1
X_4797_ VPWR VGND _2271_ net1458 _2269_ net1451 _2272_ _2265_ sg13g2_a221oi_1
X_6536_ net310 VGND VPWR net469 s0.data_out\[20\]\[5\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_20_376 VPWR VGND sg13g2_fill_1
XFILLER_20_398 VPWR VGND sg13g2_fill_1
X_3748_ net1196 VPWR _1329_ VGND net1395 net1183 sg13g2_o21ai_1
X_6467_ net1368 _0958_ _0986_ VPWR VGND sg13g2_nor2_1
X_3679_ _1269_ s0.data_out\[12\]\[6\] net1212 VPWR VGND sg13g2_nand2b_1
X_6398_ _0923_ _0922_ net1440 _0899_ net1446 VPWR VGND sg13g2_a22oi_1
X_5418_ VPWR _2836_ net461 VGND sg13g2_inv_1
X_5349_ VPWR _2767_ net459 VGND sg13g2_inv_1
XFILLER_0_726 VPWR VGND sg13g2_decap_8
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_922 VPWR VGND sg13g2_fill_1
XFILLER_29_911 VPWR VGND sg13g2_fill_2
XFILLER_29_966 VPWR VGND sg13g2_decap_8
XFILLER_44_925 VPWR VGND sg13g2_decap_8
XFILLER_28_465 VPWR VGND sg13g2_fill_1
XFILLER_15_137 VPWR VGND sg13g2_fill_1
XFILLER_7_358 VPWR VGND sg13g2_fill_1
XFILLER_11_70 VPWR VGND sg13g2_fill_1
Xfanout1310 net539 net1310 VPWR VGND sg13g2_buf_8
Xfanout1321 net1322 net1321 VPWR VGND sg13g2_buf_1
Xfanout1332 net1333 net1332 VPWR VGND sg13g2_buf_8
Xfanout1343 net1351 net1343 VPWR VGND sg13g2_buf_8
Xfanout1354 net1357 net1354 VPWR VGND sg13g2_buf_8
Xfanout1365 net1377 net1365 VPWR VGND sg13g2_buf_8
Xfanout1398 net1401 net1398 VPWR VGND sg13g2_buf_8
Xfanout1376 net1377 net1376 VPWR VGND sg13g2_buf_8
Xfanout1387 net1388 net1387 VPWR VGND sg13g2_buf_1
XFILLER_47_752 VPWR VGND sg13g2_decap_8
XFILLER_43_991 VPWR VGND sg13g2_decap_8
XFILLER_15_660 VPWR VGND sg13g2_decap_8
X_4720_ _2206_ VPWR _2207_ VGND _2166_ _2168_ sg13g2_o21ai_1
XFILLER_30_630 VPWR VGND sg13g2_decap_8
X_4651_ _2138_ net642 net1080 VPWR VGND sg13g2_nand2b_1
XFILLER_30_652 VPWR VGND sg13g2_decap_8
X_3602_ net1203 net532 _1200_ VPWR VGND sg13g2_and2_1
X_4582_ s0.data_out\[6\]\[5\] s0.data_out\[5\]\[5\] net1083 _2081_ VPWR VGND sg13g2_mux2_1
X_3533_ s0.data_out\[13\]\[0\] s0.data_out\[14\]\[0\] net1219 _1135_ VPWR VGND sg13g2_mux2_1
X_6321_ net1238 s0.data_out\[16\]\[0\] _0857_ VPWR VGND sg13g2_and2_1
XFILLER_42_0 VPWR VGND sg13g2_decap_4
X_3464_ VPWR VGND _1054_ _1077_ _1076_ _1035_ _1078_ _1075_ sg13g2_a221oi_1
X_6252_ net1239 net1169 _0789_ VPWR VGND sg13g2_nor2b_1
X_5203_ _2642_ net1031 _2641_ VPWR VGND sg13g2_nand2b_1
X_6183_ _0730_ net1251 _0731_ _0732_ VPWR VGND sg13g2_a21o_1
X_5134_ VPWR _2576_ _2575_ VGND sg13g2_inv_1
X_3395_ VGND VPWR _0893_ _1008_ _1009_ net1227 sg13g2_a21oi_1
X_5065_ VGND VPWR _2402_ _2515_ _2516_ net1039 sg13g2_a21oi_1
XFILLER_38_741 VPWR VGND sg13g2_fill_2
XFILLER_38_730 VPWR VGND sg13g2_decap_8
XFILLER_37_240 VPWR VGND sg13g2_decap_4
X_4016_ net1390 net1156 _1567_ VPWR VGND sg13g2_nor2_1
XFILLER_25_402 VPWR VGND sg13g2_fill_2
XFILLER_26_936 VPWR VGND sg13g2_decap_8
XFILLER_40_405 VPWR VGND sg13g2_fill_2
XFILLER_12_118 VPWR VGND sg13g2_fill_1
X_5967_ net1354 _0459_ _0537_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_32_clk clknet_3_4__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
XFILLER_12_129 VPWR VGND sg13g2_fill_1
X_4918_ _2381_ net1047 _2380_ VPWR VGND sg13g2_nand2b_1
XFILLER_34_991 VPWR VGND sg13g2_decap_8
X_5898_ VGND VPWR net1276 _0469_ _0471_ _0470_ sg13g2_a21oi_1
XFILLER_32_14 VPWR VGND sg13g2_decap_8
X_4849_ _2319_ VPWR _2324_ VGND _2309_ _2318_ sg13g2_o21ai_1
XFILLER_20_173 VPWR VGND sg13g2_fill_1
XFILLER_32_58 VPWR VGND sg13g2_fill_2
X_6519_ net32 VGND VPWR _0029_ s0.data_out\[21\]\[0\] clknet_leaf_4_clk sg13g2_dfrbpq_2
XFILLER_0_523 VPWR VGND sg13g2_decap_8
XFILLER_29_730 VPWR VGND sg13g2_fill_2
XFILLER_29_774 VPWR VGND sg13g2_fill_2
XFILLER_44_711 VPWR VGND sg13g2_fill_1
XFILLER_43_210 VPWR VGND sg13g2_fill_1
XFILLER_44_766 VPWR VGND sg13g2_decap_4
XFILLER_25_980 VPWR VGND sg13g2_decap_8
XFILLER_32_939 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_23_clk clknet_3_7__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_31_449 VPWR VGND sg13g2_fill_2
XFILLER_7_111 VPWR VGND sg13g2_fill_1
XFILLER_4_873 VPWR VGND sg13g2_decap_8
Xfanout1140 net1141 net1140 VPWR VGND sg13g2_buf_8
Xfanout1173 net705 net1173 VPWR VGND sg13g2_buf_8
Xfanout1151 net1155 net1151 VPWR VGND sg13g2_buf_8
Xfanout1162 net700 net1162 VPWR VGND sg13g2_buf_8
Xfanout1195 net1196 net1195 VPWR VGND sg13g2_buf_8
Xfanout1184 net1185 net1184 VPWR VGND sg13g2_buf_8
XFILLER_47_560 VPWR VGND sg13g2_decap_8
XFILLER_19_251 VPWR VGND sg13g2_fill_1
X_5821_ _0406_ _0397_ _0405_ VPWR VGND sg13g2_nand2_1
XFILLER_16_980 VPWR VGND sg13g2_decap_8
X_5752_ s0.data_out\[21\]\[1\] s0.data_out\[20\]\[1\] net1297 _0337_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_14_clk clknet_3_3__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_6637__200 VPWR VGND net200 sg13g2_tiehi
X_4703_ VGND VPWR net1062 _2189_ _2190_ _2187_ sg13g2_a21oi_1
X_5683_ _3074_ _3076_ net1426 _3077_ VPWR VGND sg13g2_nand3_1
X_4634_ _0223_ _2123_ _2124_ _2860_ net1372 VPWR VGND sg13g2_a22oi_1
XFILLER_8_71 VPWR VGND sg13g2_fill_1
X_4565_ s0.data_out\[6\]\[6\] s0.data_out\[5\]\[6\] net1083 _2064_ VPWR VGND sg13g2_mux2_1
X_6304_ net1237 net1158 _0841_ VPWR VGND sg13g2_nor2b_1
X_3516_ net1203 net1164 _1118_ VPWR VGND sg13g2_nor2b_1
X_4496_ VPWR _0208_ _2001_ VGND sg13g2_inv_1
X_6235_ VGND VPWR net1002 _0663_ _0775_ _0774_ sg13g2_a21oi_1
X_3447_ VGND VPWR net1230 _1058_ _1061_ _1060_ sg13g2_a21oi_1
X_6166_ _0715_ s0.data_out\[17\]\[6\] net1269 VPWR VGND sg13g2_nand2b_1
XFILLER_40_1009 VPWR VGND sg13g2_decap_8
X_6097_ net1264 net436 _0652_ VPWR VGND sg13g2_and2_1
X_5117_ _2562_ VPWR _2563_ VGND net1468 net583 sg13g2_o21ai_1
X_5048_ VGND VPWR net1038 _2496_ _2499_ _2498_ sg13g2_a21oi_1
XFILLER_25_232 VPWR VGND sg13g2_decap_8
XFILLER_26_755 VPWR VGND sg13g2_decap_8
X_6748__81 VPWR VGND net81 sg13g2_tiehi
XFILLER_40_268 VPWR VGND sg13g2_decap_4
XFILLER_22_994 VPWR VGND sg13g2_decap_8
XFILLER_4_103 VPWR VGND sg13g2_fill_2
XFILLER_4_125 VPWR VGND sg13g2_fill_1
XFILLER_1_821 VPWR VGND sg13g2_decap_8
XFILLER_49_814 VPWR VGND sg13g2_decap_8
XFILLER_1_898 VPWR VGND sg13g2_decap_8
XFILLER_1_1003 VPWR VGND sg13g2_decap_8
XFILLER_29_582 VPWR VGND sg13g2_fill_2
XFILLER_16_210 VPWR VGND sg13g2_fill_1
XFILLER_9_954 VPWR VGND sg13g2_decap_8
XFILLER_13_994 VPWR VGND sg13g2_decap_8
X_4350_ _1794_ VPWR _1873_ VGND _1847_ _1850_ sg13g2_o21ai_1
X_4281_ _1804_ net453 net1118 VPWR VGND sg13g2_nand2b_1
X_6020_ s0.data_out\[18\]\[0\] s0.data_out\[19\]\[0\] net1284 _0581_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_3_clk clknet_3_0__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
XFILLER_39_302 VPWR VGND sg13g2_decap_4
X_5804_ _0386_ _0387_ _0389_ VPWR VGND _0388_ sg13g2_nand3b_1
X_6784_ net78 VGND VPWR _0294_ s0.data_out\[0\]\[6\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_3996_ net1184 VPWR _1554_ VGND _1488_ _1553_ sg13g2_o21ai_1
XFILLER_22_235 VPWR VGND sg13g2_fill_1
XFILLER_22_257 VPWR VGND sg13g2_fill_1
X_5735_ net1313 VPWR _0324_ VGND _3054_ _0323_ sg13g2_o21ai_1
X_5666_ s0.data_out\[22\]\[6\] s0.data_out\[21\]\[6\] net1307 _3060_ VPWR VGND sg13g2_mux2_1
X_6745__84 VPWR VGND net84 sg13g2_tiehi
X_4617_ VGND VPWR net1075 net570 _2111_ _2074_ sg13g2_a21oi_1
X_5597_ net1324 VPWR _2998_ VGND _2964_ _2997_ sg13g2_o21ai_1
X_4548_ s0.data_out\[5\]\[2\] s0.data_out\[6\]\[2\] net1092 _2047_ VPWR VGND sg13g2_mux2_1
X_4479_ VPWR _0204_ _1988_ VGND sg13g2_inv_1
X_6218_ net1356 _0727_ _0762_ VPWR VGND sg13g2_nor2_1
XFILLER_46_806 VPWR VGND sg13g2_decap_8
Xfanout999 _2761_ net999 VPWR VGND sg13g2_buf_1
XFILLER_38_57 VPWR VGND sg13g2_fill_2
X_6149_ net1253 s0.data_new_delayed\[3\] _0698_ VPWR VGND sg13g2_nor2b_1
XFILLER_41_511 VPWR VGND sg13g2_fill_1
XFILLER_14_747 VPWR VGND sg13g2_fill_1
XFILLER_14_758 VPWR VGND sg13g2_fill_2
XFILLER_41_577 VPWR VGND sg13g2_fill_2
XFILLER_16_1022 VPWR VGND sg13g2_decap_8
XFILLER_10_931 VPWR VGND sg13g2_decap_8
XFILLER_6_935 VPWR VGND sg13g2_decap_8
XFILLER_5_412 VPWR VGND sg13g2_fill_2
XFILLER_5_445 VPWR VGND sg13g2_decap_4
XFILLER_5_489 VPWR VGND sg13g2_fill_1
XFILLER_49_611 VPWR VGND sg13g2_decap_8
XFILLER_1_695 VPWR VGND sg13g2_decap_8
XFILLER_23_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_688 VPWR VGND sg13g2_decap_8
XFILLER_48_187 VPWR VGND sg13g2_decap_4
XFILLER_45_872 VPWR VGND sg13g2_fill_2
XFILLER_45_861 VPWR VGND sg13g2_fill_2
XFILLER_45_850 VPWR VGND sg13g2_decap_8
X_3850_ _1425_ VPWR _1426_ VGND net1016 _1424_ sg13g2_o21ai_1
XFILLER_20_717 VPWR VGND sg13g2_decap_4
X_3781_ _1360_ net1335 _1358_ VPWR VGND sg13g2_xnor2_1
X_5520_ _2924_ net1315 _2925_ _2926_ VPWR VGND sg13g2_a21o_1
X_5451_ VPWR _2869_ net492 VGND sg13g2_inv_1
X_6742__87 VPWR VGND net87 sg13g2_tiehi
X_5382_ VPWR _2800_ net410 VGND sg13g2_inv_1
X_4402_ _1911_ net1086 _1912_ _1913_ VPWR VGND sg13g2_a21o_1
X_4333_ _1854_ net1102 _1855_ _1856_ VPWR VGND sg13g2_a21o_1
XFILLER_5_990 VPWR VGND sg13g2_decap_8
X_4264_ _0187_ _1789_ _1790_ _2846_ net1384 VPWR VGND sg13g2_a22oi_1
X_6003_ net1266 net1162 _0564_ VPWR VGND sg13g2_nor2b_1
X_4195_ _1730_ net371 net1132 VPWR VGND sg13g2_nand2b_1
XFILLER_28_839 VPWR VGND sg13g2_fill_2
XFILLER_36_894 VPWR VGND sg13g2_fill_2
XFILLER_35_382 VPWR VGND sg13g2_fill_1
XFILLER_11_706 VPWR VGND sg13g2_fill_1
XFILLER_24_26 VPWR VGND sg13g2_decap_8
XFILLER_24_37 VPWR VGND sg13g2_fill_1
XFILLER_10_216 VPWR VGND sg13g2_fill_1
X_6767_ net23 VGND VPWR net495 s0.data_out\[1\]\[1\] clknet_leaf_8_clk sg13g2_dfrbpq_2
XFILLER_10_227 VPWR VGND sg13g2_decap_8
X_5718_ net1341 _3037_ _0311_ VPWR VGND sg13g2_nor2_1
X_3979_ net1384 _1482_ _1541_ VPWR VGND sg13g2_nor2_1
X_6698_ net135 VGND VPWR _0208_ s0.data_out\[7\]\[4\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_5649_ s0.data_out\[21\]\[2\] s0.data_out\[22\]\[2\] net1320 _3043_ VPWR VGND sg13g2_mux2_1
Xhold261 _0270_ VPWR VGND net581 sg13g2_dlygate4sd3_1
Xhold250 s0.data_out\[5\]\[4\] VPWR VGND net570 sg13g2_dlygate4sd3_1
XFILLER_2_448 VPWR VGND sg13g2_fill_1
Xhold294 _1670_ VPWR VGND net614 sg13g2_dlygate4sd3_1
Xhold283 s0.data_out\[22\]\[0\] VPWR VGND net603 sg13g2_dlygate4sd3_1
Xhold272 _1193_ VPWR VGND net592 sg13g2_dlygate4sd3_1
XFILLER_49_56 VPWR VGND sg13g2_decap_8
XFILLER_42_853 VPWR VGND sg13g2_fill_2
XFILLER_14_70 VPWR VGND sg13g2_decap_4
XFILLER_49_430 VPWR VGND sg13g2_fill_1
XFILLER_49_463 VPWR VGND sg13g2_fill_1
X_4951_ net1040 net1152 _2414_ VPWR VGND sg13g2_nor2b_1
X_4882_ net1361 _2295_ _2350_ VPWR VGND sg13g2_nor2_1
X_3902_ VGND VPWR net1179 _1465_ _1468_ _1467_ sg13g2_a21oi_1
X_6621_ net218 VGND VPWR _0131_ s0.data_out\[13\]\[6\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_3833_ _1406_ VPWR _1412_ VGND _1399_ _1409_ sg13g2_o21ai_1
XFILLER_32_363 VPWR VGND sg13g2_fill_2
XFILLER_32_374 VPWR VGND sg13g2_fill_2
X_6552_ net292 VGND VPWR _0062_ s0.valid_out\[18\][0] clknet_leaf_36_clk sg13g2_dfrbpq_1
XFILLER_9_570 VPWR VGND sg13g2_decap_4
X_3764_ VGND VPWR _1234_ _1342_ _1343_ net1191 sg13g2_a21oi_1
X_6483_ _0996_ VPWR _0999_ VGND s0.was_valid_out\[14\][0] net1221 sg13g2_o21ai_1
X_3695_ net1196 net1159 _1285_ VPWR VGND sg13g2_nor2b_1
X_5503_ net1315 net1162 _2909_ VPWR VGND sg13g2_nor2b_1
X_5434_ VPWR _2852_ net518 VGND sg13g2_inv_1
XFILLER_0_908 VPWR VGND sg13g2_decap_8
X_5365_ VPWR _2783_ s0.data_out\[21\]\[0\] VGND sg13g2_inv_1
X_4316_ VGND VPWR net1114 _1836_ _1839_ _1838_ sg13g2_a21oi_1
X_5296_ net547 net1346 _2721_ _0288_ VPWR VGND sg13g2_a21o_1
X_4247_ net1000 _2850_ _1777_ VPWR VGND sg13g2_nor2_1
X_6569__274 VPWR VGND net274 sg13g2_tiehi
X_4178_ _1711_ net1113 _1712_ _1713_ VPWR VGND sg13g2_a21o_1
XFILLER_35_36 VPWR VGND sg13g2_fill_2
XFILLER_35_47 VPWR VGND sg13g2_fill_1
XFILLER_3_768 VPWR VGND sg13g2_decap_8
XFILLER_2_234 VPWR VGND sg13g2_fill_1
XFILLER_47_934 VPWR VGND sg13g2_decap_8
XFILLER_18_113 VPWR VGND sg13g2_decap_8
XFILLER_19_625 VPWR VGND sg13g2_fill_2
XFILLER_20_1018 VPWR VGND sg13g2_decap_8
XFILLER_14_374 VPWR VGND sg13g2_decap_8
XFILLER_41_171 VPWR VGND sg13g2_decap_8
X_3480_ net1227 VPWR _1090_ VGND _1029_ _1089_ sg13g2_o21ai_1
XFILLER_44_4 VPWR VGND sg13g2_fill_2
X_5150_ _2589_ net375 net1033 VPWR VGND sg13g2_nand2b_1
X_4101_ VGND VPWR _1648_ net1331 net329 sg13g2_or2_1
X_5081_ _2532_ net1039 _2531_ VPWR VGND sg13g2_nand2b_1
X_4032_ s0.data_out\[10\]\[0\] s0.data_out\[9\]\[0\] net1131 _1579_ VPWR VGND sg13g2_mux2_1
XFILLER_38_956 VPWR VGND sg13g2_decap_8
X_5983_ net1352 _0498_ _0549_ VPWR VGND sg13g2_nor2_1
X_4934_ net1040 net1142 _2397_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_1014 VPWR VGND sg13g2_decap_8
XFILLER_21_801 VPWR VGND sg13g2_fill_2
XFILLER_21_834 VPWR VGND sg13g2_fill_1
X_4865_ _0242_ _2335_ _2336_ _2872_ net1359 VPWR VGND sg13g2_a22oi_1
X_6604_ net236 VGND VPWR _0114_ s0.data_out\[14\]\[1\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3816_ VGND VPWR net1183 _1394_ _1395_ _1392_ sg13g2_a21oi_1
X_4796_ _2271_ net995 _2270_ VPWR VGND sg13g2_nand2_1
X_6535_ net311 VGND VPWR net497 s0.data_out\[20\]\[4\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_3747_ _0132_ _1327_ _1328_ _2825_ net1382 VPWR VGND sg13g2_a22oi_1
X_6466_ net1241 VPWR _0985_ VGND _0955_ _0984_ sg13g2_o21ai_1
X_3678_ _1266_ net1194 _1267_ _1268_ VPWR VGND sg13g2_a21o_1
XFILLER_0_705 VPWR VGND sg13g2_decap_8
X_6397_ VGND VPWR net1242 _0919_ _0922_ _0921_ sg13g2_a21oi_1
X_5417_ VPWR _2835_ net373 VGND sg13g2_inv_1
X_5348_ VPWR _2766_ net455 VGND sg13g2_inv_1
X_5279_ _2706_ _2768_ _2705_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_422 VPWR VGND sg13g2_fill_2
XFILLER_29_945 VPWR VGND sg13g2_decap_8
XFILLER_44_904 VPWR VGND sg13g2_decap_8
X_6582__260 VPWR VGND net260 sg13g2_tiehi
XFILLER_16_606 VPWR VGND sg13g2_fill_2
XFILLER_11_300 VPWR VGND sg13g2_fill_1
XFILLER_11_60 VPWR VGND sg13g2_fill_1
XFILLER_3_532 VPWR VGND sg13g2_fill_1
XFILLER_2_0 VPWR VGND sg13g2_fill_2
XFILLER_11_82 VPWR VGND sg13g2_decap_4
XFILLER_39_709 VPWR VGND sg13g2_fill_1
Xfanout1311 net1314 net1311 VPWR VGND sg13g2_buf_8
Xfanout1322 s0.valid_out\[22\][0] net1322 VPWR VGND sg13g2_buf_2
Xfanout1300 net1302 net1300 VPWR VGND sg13g2_buf_8
Xfanout1344 net1351 net1344 VPWR VGND sg13g2_buf_8
Xfanout1355 net1356 net1355 VPWR VGND sg13g2_buf_8
Xfanout1366 net1377 net1366 VPWR VGND sg13g2_buf_2
Xfanout1333 _2983_ net1333 VPWR VGND sg13g2_buf_8
XFILLER_47_731 VPWR VGND sg13g2_decap_8
Xfanout1399 net1401 net1399 VPWR VGND sg13g2_buf_2
Xfanout1377 net1389 net1377 VPWR VGND sg13g2_buf_8
Xfanout1388 net1389 net1388 VPWR VGND sg13g2_buf_8
XFILLER_19_466 VPWR VGND sg13g2_decap_8
XFILLER_43_970 VPWR VGND sg13g2_decap_8
XFILLER_15_694 VPWR VGND sg13g2_fill_2
X_4650_ _2135_ net1061 _2136_ _2137_ VPWR VGND sg13g2_a21o_1
X_3601_ _0115_ _1198_ _1199_ _2823_ net1380 VPWR VGND sg13g2_a22oi_1
X_4581_ _2077_ _2079_ net1430 _2080_ VPWR VGND sg13g2_nand3_1
X_6320_ net322 net1331 _0856_ _0076_ VPWR VGND sg13g2_nor3_1
X_3532_ _1134_ net1214 _1133_ VPWR VGND sg13g2_nand2b_1
X_3463_ _0998_ VPWR _1077_ VGND _1050_ _1053_ sg13g2_o21ai_1
X_6251_ VGND VPWR _0788_ _0787_ net1447 sg13g2_or2_1
X_5202_ VGND VPWR net1022 _2639_ _2641_ _2640_ sg13g2_a21oi_1
X_6182_ net1249 net1153 _0731_ VPWR VGND sg13g2_nor2b_1
X_5133_ VGND VPWR net1336 net1025 _2575_ _2574_ sg13g2_a21oi_1
X_3394_ _1008_ s0.data_out\[14\]\[2\] net1232 VPWR VGND sg13g2_nand2b_1
XFILLER_35_0 VPWR VGND sg13g2_decap_4
X_5064_ _2515_ s0.data_out\[1\]\[6\] net1045 VPWR VGND sg13g2_nand2b_1
X_6566__277 VPWR VGND net277 sg13g2_tiehi
X_4015_ _1566_ VPWR _0162_ VGND net1391 net993 sg13g2_o21ai_1
XFILLER_41_907 VPWR VGND sg13g2_fill_2
XFILLER_40_417 VPWR VGND sg13g2_fill_2
X_5966_ net1293 VPWR _0536_ VGND _0456_ _0535_ sg13g2_o21ai_1
XFILLER_34_970 VPWR VGND sg13g2_decap_8
X_5897_ net1276 net1173 _0470_ VPWR VGND sg13g2_nor2b_1
X_4917_ VGND VPWR net1036 _2378_ _2380_ _2379_ sg13g2_a21oi_1
X_4848_ _2301_ _2309_ _2320_ _2322_ _2323_ VPWR VGND sg13g2_and4_1
XFILLER_21_664 VPWR VGND sg13g2_fill_2
X_4779_ _2252_ net1049 _2253_ _2254_ VPWR VGND sg13g2_a21o_1
X_6518_ net33 VGND VPWR _0028_ s0.shift_out\[21\][0] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_4_318 VPWR VGND sg13g2_fill_1
X_6449_ net1225 s0.data_out\[15\]\[1\] _0972_ VPWR VGND sg13g2_and2_1
XFILLER_0_502 VPWR VGND sg13g2_decap_8
XFILLER_0_579 VPWR VGND sg13g2_decap_8
XFILLER_48_528 VPWR VGND sg13g2_fill_1
XFILLER_16_458 VPWR VGND sg13g2_decap_8
XFILLER_40_995 VPWR VGND sg13g2_decap_8
XFILLER_8_646 VPWR VGND sg13g2_fill_1
XFILLER_7_189 VPWR VGND sg13g2_fill_1
XFILLER_4_852 VPWR VGND sg13g2_decap_8
XFILLER_26_1013 VPWR VGND sg13g2_decap_8
Xfanout1141 net360 net1141 VPWR VGND sg13g2_buf_8
Xfanout1130 s0.shift_out\[9\][0] net1130 VPWR VGND sg13g2_buf_1
Xfanout1174 net1177 net1174 VPWR VGND sg13g2_buf_8
Xfanout1152 net1155 net1152 VPWR VGND sg13g2_buf_2
Xfanout1163 s0.data_new_delayed\[2\] net1163 VPWR VGND sg13g2_buf_1
Xfanout1196 net391 net1196 VPWR VGND sg13g2_buf_8
Xfanout1185 net1186 net1185 VPWR VGND sg13g2_buf_8
XFILLER_35_778 VPWR VGND sg13g2_fill_2
X_5820_ _0402_ _0404_ net1418 _0405_ VPWR VGND sg13g2_nand3_1
XFILLER_15_480 VPWR VGND sg13g2_fill_1
X_5751_ _0336_ net1297 net633 VPWR VGND sg13g2_nand2_1
XFILLER_22_428 VPWR VGND sg13g2_fill_2
XFILLER_34_299 VPWR VGND sg13g2_fill_1
X_6757__71 VPWR VGND net71 sg13g2_tiehi
X_4702_ s0.data_out\[5\]\[4\] s0.data_out\[4\]\[4\] net1068 _2189_ VPWR VGND sg13g2_mux2_1
X_5682_ _3076_ net1012 _3075_ VPWR VGND sg13g2_nand2_1
XFILLER_30_472 VPWR VGND sg13g2_decap_8
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
X_4633_ net1372 net405 _2124_ VPWR VGND sg13g2_nor2_1
XFILLER_8_61 VPWR VGND sg13g2_fill_2
X_4564_ _2063_ net1082 net449 VPWR VGND sg13g2_nand2_1
X_6303_ _0840_ net1421 _0839_ VPWR VGND sg13g2_nand2_1
X_3515_ s0.data_out\[14\]\[2\] s0.data_out\[13\]\[2\] net1210 _1117_ VPWR VGND sg13g2_mux2_1
X_4495_ _2000_ VPWR _2001_ VGND net1479 net639 sg13g2_o21ai_1
X_6234_ VGND VPWR net1337 net1245 _0774_ _0773_ sg13g2_a21oi_1
X_3446_ VGND VPWR _0953_ _1059_ _1060_ net1230 sg13g2_a21oi_1
X_6165_ _0712_ net1249 _0713_ _0714_ VPWR VGND sg13g2_a21o_1
X_6096_ _0057_ _0650_ _0651_ _2793_ net1353 VPWR VGND sg13g2_a22oi_1
X_5116_ _2561_ VPWR _2562_ VGND net1010 _2560_ sg13g2_o21ai_1
XFILLER_45_509 VPWR VGND sg13g2_fill_2
X_5047_ VGND VPWR _2387_ _2497_ _2498_ net1038 sg13g2_a21oi_1
XFILLER_27_48 VPWR VGND sg13g2_fill_2
X_5949_ net1427 _0511_ _0522_ VPWR VGND sg13g2_nor2_1
XFILLER_22_973 VPWR VGND sg13g2_decap_8
XFILLER_5_627 VPWR VGND sg13g2_fill_1
XFILLER_49_1024 VPWR VGND sg13g2_decap_4
XFILLER_1_800 VPWR VGND sg13g2_decap_8
XFILLER_0_310 VPWR VGND sg13g2_fill_2
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_1_877 VPWR VGND sg13g2_decap_8
XFILLER_44_542 VPWR VGND sg13g2_fill_2
XFILLER_32_726 VPWR VGND sg13g2_fill_1
XFILLER_9_933 VPWR VGND sg13g2_decap_8
XFILLER_13_973 VPWR VGND sg13g2_decap_8
X_6754__74 VPWR VGND net74 sg13g2_tiehi
X_4280_ _1801_ net1099 _1802_ _1803_ VPWR VGND sg13g2_a21o_1
XFILLER_35_531 VPWR VGND sg13g2_fill_2
XFILLER_35_597 VPWR VGND sg13g2_fill_2
X_5803_ net1398 _0378_ _0388_ VPWR VGND sg13g2_nor2_1
XFILLER_22_203 VPWR VGND sg13g2_fill_1
X_6783_ net91 VGND VPWR _0293_ s0.data_out\[0\]\[5\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_3995_ _2746_ _2841_ _1553_ VPWR VGND sg13g2_nor2_1
X_5734_ net1008 _2779_ _0323_ VPWR VGND sg13g2_nor2_1
X_5665_ _3059_ net1308 net650 VPWR VGND sg13g2_nand2_1
XFILLER_31_792 VPWR VGND sg13g2_fill_2
X_4616_ _0219_ net447 _2110_ _2862_ net1370 VPWR VGND sg13g2_a22oi_1
X_5596_ net1312 s0.data_out\[22\]\[4\] _2997_ VPWR VGND sg13g2_and2_1
X_4547_ VGND VPWR net1074 _2044_ _2046_ _2045_ sg13g2_a21oi_1
X_4478_ _1987_ VPWR _1988_ VGND net1479 net521 sg13g2_o21ai_1
X_3429_ _1043_ net1221 net545 VPWR VGND sg13g2_nand2_1
X_6217_ net1268 VPWR _0761_ VGND _0724_ _0760_ sg13g2_o21ai_1
X_6148_ s0.data_out\[18\]\[3\] s0.data_out\[17\]\[3\] net1259 _0697_ VPWR VGND sg13g2_mux2_1
XFILLER_45_306 VPWR VGND sg13g2_fill_2
X_6079_ _0638_ VPWR _0639_ VGND net1471 net597 sg13g2_o21ai_1
XFILLER_14_704 VPWR VGND sg13g2_fill_1
XFILLER_13_203 VPWR VGND sg13g2_fill_2
XFILLER_26_575 VPWR VGND sg13g2_fill_1
XFILLER_41_545 VPWR VGND sg13g2_decap_4
XFILLER_13_236 VPWR VGND sg13g2_decap_8
XFILLER_16_1001 VPWR VGND sg13g2_decap_8
XFILLER_6_914 VPWR VGND sg13g2_decap_8
XFILLER_10_987 VPWR VGND sg13g2_decap_8
X_6751__77 VPWR VGND net77 sg13g2_tiehi
XFILLER_1_674 VPWR VGND sg13g2_decap_8
X_6627__211 VPWR VGND net211 sg13g2_tiehi
XFILLER_49_667 VPWR VGND sg13g2_decap_8
XFILLER_0_195 VPWR VGND sg13g2_fill_2
XFILLER_17_531 VPWR VGND sg13g2_decap_4
XFILLER_29_391 VPWR VGND sg13g2_decap_8
XFILLER_32_556 VPWR VGND sg13g2_decap_8
X_3780_ VGND VPWR _1359_ _1358_ net1335 sg13g2_or2_1
XFILLER_32_589 VPWR VGND sg13g2_fill_2
XFILLER_9_752 VPWR VGND sg13g2_decap_4
X_6634__204 VPWR VGND net204 sg13g2_tiehi
X_5450_ VPWR _2868_ net449 VGND sg13g2_inv_1
X_4401_ net1085 net1165 _1912_ VPWR VGND sg13g2_nor2b_1
X_5381_ VPWR _2799_ net440 VGND sg13g2_inv_1
X_4332_ net1102 net1153 _1855_ VPWR VGND sg13g2_nor2b_1
X_4263_ net1384 net372 _1790_ VPWR VGND sg13g2_nor2_1
XFILLER_4_490 VPWR VGND sg13g2_fill_1
X_6002_ s0.data_out\[19\]\[2\] s0.data_out\[18\]\[2\] net1270 _0563_ VPWR VGND sg13g2_mux2_1
X_4194_ _1727_ net1117 _1728_ _1729_ VPWR VGND sg13g2_a21o_1
XFILLER_39_111 VPWR VGND sg13g2_fill_2
XFILLER_39_188 VPWR VGND sg13g2_decap_4
XFILLER_23_512 VPWR VGND sg13g2_decap_4
XFILLER_10_206 VPWR VGND sg13g2_fill_1
X_6766_ net36 VGND VPWR _0276_ s0.data_out\[1\]\[0\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_3978_ net1181 VPWR _1540_ VGND _1479_ _1539_ sg13g2_o21ai_1
X_5717_ net1316 VPWR _0310_ VGND _3034_ _0309_ sg13g2_o21ai_1
X_6697_ net136 VGND VPWR _0207_ s0.data_out\[7\]\[3\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5648_ VGND VPWR net1304 _3040_ _3042_ _3041_ sg13g2_a21oi_1
X_5579_ VGND VPWR _2979_ _2982_ _0004_ _2984_ sg13g2_a21oi_1
Xhold240 s0.data_out\[17\]\[7\] VPWR VGND net560 sg13g2_dlygate4sd3_1
Xhold262 s0.data_out\[2\]\[2\] VPWR VGND net582 sg13g2_dlygate4sd3_1
Xhold251 s0.data_out\[5\]\[0\] VPWR VGND net571 sg13g2_dlygate4sd3_1
XFILLER_49_35 VPWR VGND sg13g2_decap_8
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_1016 VPWR VGND sg13g2_decap_8
Xhold295 s0.was_valid_out\[14\][0] VPWR VGND net615 sg13g2_dlygate4sd3_1
Xhold273 s0.data_out\[22\]\[6\] VPWR VGND net593 sg13g2_dlygate4sd3_1
Xhold284 _0017_ VPWR VGND net604 sg13g2_dlygate4sd3_1
XFILLER_49_79 VPWR VGND sg13g2_decap_4
XFILLER_45_147 VPWR VGND sg13g2_fill_2
XFILLER_27_873 VPWR VGND sg13g2_fill_2
XFILLER_14_545 VPWR VGND sg13g2_decap_8
XFILLER_10_784 VPWR VGND sg13g2_fill_1
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_2_994 VPWR VGND sg13g2_decap_8
XFILLER_49_442 VPWR VGND sg13g2_decap_8
XFILLER_37_615 VPWR VGND sg13g2_decap_4
XFILLER_49_497 VPWR VGND sg13g2_decap_4
X_4950_ s0.data_out\[3\]\[5\] s0.data_out\[2\]\[5\] net1045 _2413_ VPWR VGND sg13g2_mux2_1
XFILLER_33_832 VPWR VGND sg13g2_fill_1
X_4881_ net1064 VPWR _2349_ VGND _2292_ _2348_ sg13g2_o21ai_1
X_3901_ VGND VPWR _1338_ _1466_ _1467_ net1178 sg13g2_a21oi_1
XFILLER_33_843 VPWR VGND sg13g2_decap_8
X_6620_ net219 VGND VPWR _0130_ s0.data_out\[13\]\[5\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_3832_ _1373_ _1391_ _1407_ _1410_ _1411_ VPWR VGND sg13g2_or4_1
X_6551_ net294 VGND VPWR net544 s0.was_valid_out\[18\][0] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_32_386 VPWR VGND sg13g2_fill_1
X_5502_ s0.data_out\[23\]\[2\] s0.data_out\[22\]\[2\] net1320 _2908_ VPWR VGND sg13g2_mux2_1
X_3763_ _1342_ s0.data_out\[11\]\[1\] net1197 VPWR VGND sg13g2_nand2b_1
X_6482_ _0996_ _0997_ _0998_ VPWR VGND sg13g2_nor2_1
X_3694_ s0.data_out\[13\]\[4\] s0.data_out\[12\]\[4\] net1198 _1284_ VPWR VGND sg13g2_mux2_1
X_5433_ VPWR _2851_ net637 VGND sg13g2_inv_1
X_5364_ VPWR _2782_ net557 VGND sg13g2_inv_1
X_4315_ VGND VPWR _1719_ _1837_ _1838_ net1115 sg13g2_a21oi_1
X_5295_ VGND VPWR _2692_ _2693_ _2721_ net1346 sg13g2_a21oi_1
X_4246_ _0183_ _1775_ _1776_ _2844_ net1375 VPWR VGND sg13g2_a22oi_1
X_4177_ net1112 net994 _1712_ VPWR VGND sg13g2_nor2_1
XFILLER_43_629 VPWR VGND sg13g2_fill_2
XFILLER_42_139 VPWR VGND sg13g2_fill_2
XFILLER_11_526 VPWR VGND sg13g2_decap_4
XFILLER_11_537 VPWR VGND sg13g2_decap_4
X_6749_ net80 VGND VPWR net485 s0.data_out\[3\]\[7\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_13_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_747 VPWR VGND sg13g2_decap_8
XFILLER_47_913 VPWR VGND sg13g2_decap_8
XFILLER_19_604 VPWR VGND sg13g2_decap_4
X_6624__214 VPWR VGND net214 sg13g2_tiehi
XFILLER_46_489 VPWR VGND sg13g2_fill_2
XFILLER_27_681 VPWR VGND sg13g2_decap_4
XFILLER_33_139 VPWR VGND sg13g2_fill_1
X_6631__207 VPWR VGND net207 sg13g2_tiehi
XFILLER_29_1022 VPWR VGND sg13g2_decap_8
X_4100_ _1645_ _1646_ _1647_ VPWR VGND sg13g2_nor2_1
X_5080_ VGND VPWR net1030 _2529_ _2531_ _2530_ sg13g2_a21oi_1
XFILLER_2_791 VPWR VGND sg13g2_decap_8
X_4031_ _1578_ net1131 net596 VPWR VGND sg13g2_nand2_1
XFILLER_49_272 VPWR VGND sg13g2_decap_8
XFILLER_38_935 VPWR VGND sg13g2_decap_8
XFILLER_37_412 VPWR VGND sg13g2_fill_2
X_5982_ net1287 VPWR _0548_ VGND _0495_ _0547_ sg13g2_o21ai_1
X_4933_ s0.data_out\[3\]\[7\] s0.data_out\[2\]\[7\] net1046 _2396_ VPWR VGND sg13g2_mux2_1
X_4864_ net1359 _2256_ _2336_ VPWR VGND sg13g2_nor2_1
X_6603_ net237 VGND VPWR _0113_ s0.data_out\[14\]\[0\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3815_ s0.data_out\[12\]\[4\] s0.data_out\[11\]\[4\] net1188 _1394_ VPWR VGND sg13g2_mux2_1
X_4795_ s0.data_out\[3\]\[0\] s0.data_out\[4\]\[0\] net1067 _2270_ VPWR VGND sg13g2_mux2_1
X_3746_ net1382 _1263_ _1328_ VPWR VGND sg13g2_nor2_1
X_6534_ net312 VGND VPWR net629 s0.data_out\[20\]\[3\] clknet_leaf_4_clk sg13g2_dfrbpq_2
XFILLER_20_389 VPWR VGND sg13g2_decap_8
X_6465_ net1224 net430 _0984_ VPWR VGND sg13g2_and2_1
X_5416_ VPWR _2834_ net451 VGND sg13g2_inv_1
X_3677_ net1194 net1150 _1267_ VPWR VGND sg13g2_nor2b_1
X_6396_ VGND VPWR _0804_ _0920_ _0921_ net1242 sg13g2_a21oi_1
X_5347_ VPWR _2765_ net593 VGND sg13g2_inv_1
XFILLER_43_1019 VPWR VGND sg13g2_decap_8
X_5278_ _2704_ VPWR _2705_ VGND net1001 net1156 sg13g2_o21ai_1
X_4229_ VGND VPWR _1758_ _1762_ _0179_ _1763_ sg13g2_a21oi_1
XFILLER_29_913 VPWR VGND sg13g2_fill_1
XFILLER_43_404 VPWR VGND sg13g2_fill_2
XFILLER_16_629 VPWR VGND sg13g2_fill_2
XFILLER_7_305 VPWR VGND sg13g2_fill_1
XFILLER_11_356 VPWR VGND sg13g2_decap_8
XFILLER_7_316 VPWR VGND sg13g2_fill_1
Xfanout1312 net1314 net1312 VPWR VGND sg13g2_buf_1
Xfanout1301 net1302 net1301 VPWR VGND sg13g2_buf_8
Xfanout1323 net1324 net1323 VPWR VGND sg13g2_buf_8
Xfanout1356 net1357 net1356 VPWR VGND sg13g2_buf_8
Xfanout1345 net1351 net1345 VPWR VGND sg13g2_buf_1
Xfanout1334 _2774_ net1334 VPWR VGND sg13g2_buf_8
XFILLER_47_710 VPWR VGND sg13g2_decap_8
XFILLER_4_1013 VPWR VGND sg13g2_decap_8
Xfanout1367 net1369 net1367 VPWR VGND sg13g2_buf_8
Xfanout1378 net1383 net1378 VPWR VGND sg13g2_buf_8
Xfanout1389 _2742_ net1389 VPWR VGND sg13g2_buf_8
XFILLER_46_231 VPWR VGND sg13g2_decap_4
XFILLER_47_787 VPWR VGND sg13g2_decap_8
XFILLER_28_990 VPWR VGND sg13g2_decap_8
XFILLER_42_470 VPWR VGND sg13g2_decap_8
X_4580_ _2079_ net999 _2078_ VPWR VGND sg13g2_nand2_1
X_6559__285 VPWR VGND net285 sg13g2_tiehi
X_3600_ net1380 _1121_ _1199_ VPWR VGND sg13g2_nor2_1
X_3531_ VGND VPWR net1201 _1131_ _1133_ _1132_ sg13g2_a21oi_1
X_3462_ _1071_ VPWR _1076_ VGND _1062_ _1070_ sg13g2_o21ai_1
X_6250_ VGND VPWR net1254 _0784_ _0787_ _0786_ sg13g2_a21oi_1
X_5201_ net1023 net1151 _2640_ VPWR VGND sg13g2_nor2b_1
X_6181_ s0.data_out\[18\]\[5\] s0.data_out\[17\]\[5\] net1258 _0730_ VPWR VGND sg13g2_mux2_1
X_3393_ _1005_ net1215 _1006_ _1007_ VPWR VGND sg13g2_a21o_1
X_5132_ net1031 VPWR _2574_ VGND net1392 net1022 sg13g2_o21ai_1
X_5063_ _2512_ net1030 _2513_ _2514_ VPWR VGND sg13g2_a21o_1
X_4014_ _1566_ net1391 net1435 VPWR VGND sg13g2_nand2_1
XFILLER_25_404 VPWR VGND sg13g2_fill_1
XFILLER_40_407 VPWR VGND sg13g2_fill_1
X_5965_ net1003 _2795_ _0535_ VPWR VGND sg13g2_nor2_1
X_5896_ s0.data_out\[20\]\[0\] s0.data_out\[19\]\[0\] net1283 _0469_ VPWR VGND sg13g2_mux2_1
XFILLER_21_610 VPWR VGND sg13g2_fill_2
X_4916_ net1036 net1173 _2379_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_470 VPWR VGND sg13g2_fill_1
X_4847_ _2310_ _2321_ _2322_ VPWR VGND sg13g2_nor2_1
XFILLER_21_676 VPWR VGND sg13g2_decap_8
X_4778_ net1049 net1163 _2253_ VPWR VGND sg13g2_nor2b_1
X_6517_ net34 VGND VPWR _0027_ s0.genblk1\[20\].modules.bubble clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_3729_ _0128_ _1313_ _1314_ _2827_ net1379 VPWR VGND sg13g2_a22oi_1
X_6448_ VPWR _0089_ _0971_ VGND sg13g2_inv_1
X_6379_ _0902_ net1226 _0903_ _0904_ VPWR VGND sg13g2_a21o_1
XFILLER_0_558 VPWR VGND sg13g2_decap_8
XFILLER_29_721 VPWR VGND sg13g2_decap_4
XFILLER_28_286 VPWR VGND sg13g2_fill_2
XFILLER_32_919 VPWR VGND sg13g2_fill_1
XFILLER_19_1021 VPWR VGND sg13g2_decap_8
XFILLER_12_643 VPWR VGND sg13g2_fill_1
XFILLER_40_974 VPWR VGND sg13g2_decap_8
XFILLER_8_636 VPWR VGND sg13g2_fill_1
XFILLER_8_625 VPWR VGND sg13g2_fill_2
XFILLER_7_135 VPWR VGND sg13g2_decap_8
XFILLER_4_831 VPWR VGND sg13g2_decap_8
XFILLER_3_363 VPWR VGND sg13g2_decap_4
Xfanout1120 s0.valid_out\[8\][0] net1120 VPWR VGND sg13g2_buf_8
Xfanout1131 net1133 net1131 VPWR VGND sg13g2_buf_8
XFILLER_39_529 VPWR VGND sg13g2_fill_1
XFILLER_39_518 VPWR VGND sg13g2_fill_1
Xfanout1153 net1155 net1153 VPWR VGND sg13g2_buf_8
Xfanout1142 net1146 net1142 VPWR VGND sg13g2_buf_8
Xfanout1164 net1165 net1164 VPWR VGND sg13g2_buf_8
Xfanout1175 net1176 net1175 VPWR VGND sg13g2_buf_8
Xfanout1197 net1200 net1197 VPWR VGND sg13g2_buf_8
Xfanout1186 s0.shift_out\[11\][0] net1186 VPWR VGND sg13g2_buf_8
X_5750_ net1472 net338 _0027_ VPWR VGND sg13g2_and2_1
X_5681_ s0.data_out\[21\]\[4\] s0.data_out\[22\]\[4\] net1321 _3075_ VPWR VGND sg13g2_mux2_1
XFILLER_33_1007 VPWR VGND sg13g2_decap_8
X_4701_ _2188_ net1067 s0.data_out\[4\]\[4\] VPWR VGND sg13g2_nand2_1
X_4632_ net1088 VPWR _2123_ VGND _2058_ _2122_ sg13g2_o21ai_1
XFILLER_31_985 VPWR VGND sg13g2_decap_8
X_4563_ VGND VPWR net1088 _2059_ _2062_ _2061_ sg13g2_a21oi_1
X_4494_ _1972_ _1999_ net1479 _2000_ VPWR VGND sg13g2_nand3_1
X_6302_ VGND VPWR net1251 _0836_ _0839_ _0838_ sg13g2_a21oi_1
X_6572__271 VPWR VGND net271 sg13g2_tiehi
X_3514_ _1116_ net1212 net457 VPWR VGND sg13g2_nand2_1
X_6233_ net1250 VPWR _0773_ VGND net1394 net1236 sg13g2_o21ai_1
X_3445_ _1059_ s0.data_out\[14\]\[5\] net1234 VPWR VGND sg13g2_nand2b_1
X_6164_ net1249 net1148 _0713_ VPWR VGND sg13g2_nor2b_1
X_5115_ VGND VPWR net1009 _2526_ _2561_ net1349 sg13g2_a21oi_1
X_6095_ net1352 _0618_ _0651_ VPWR VGND sg13g2_nor2_1
X_5046_ _2497_ s0.data_out\[1\]\[3\] net1043 VPWR VGND sg13g2_nand2b_1
XFILLER_26_713 VPWR VGND sg13g2_decap_8
XFILLER_38_584 VPWR VGND sg13g2_fill_2
XFILLER_41_705 VPWR VGND sg13g2_decap_4
XFILLER_25_267 VPWR VGND sg13g2_fill_1
X_5948_ net1418 _0518_ _0521_ VPWR VGND sg13g2_nor2_1
XFILLER_40_248 VPWR VGND sg13g2_fill_2
X_5879_ net1352 _0447_ _0038_ VPWR VGND sg13g2_nor2_1
X_6763__64 VPWR VGND net64 sg13g2_tiehi
XFILLER_4_105 VPWR VGND sg13g2_fill_1
XFILLER_49_1003 VPWR VGND sg13g2_decap_8
XFILLER_4_116 VPWR VGND sg13g2_fill_1
XFILLER_1_856 VPWR VGND sg13g2_decap_8
XFILLER_49_849 VPWR VGND sg13g2_decap_8
XFILLER_48_337 VPWR VGND sg13g2_decap_8
XFILLER_29_540 VPWR VGND sg13g2_fill_1
XFILLER_29_584 VPWR VGND sg13g2_fill_1
XFILLER_17_71 VPWR VGND sg13g2_decap_8
XFILLER_44_576 VPWR VGND sg13g2_decap_4
XFILLER_13_952 VPWR VGND sg13g2_decap_8
XFILLER_9_989 VPWR VGND sg13g2_decap_8
X_6556__288 VPWR VGND net288 sg13g2_tiehi
XFILLER_4_683 VPWR VGND sg13g2_decap_8
XFILLER_48_893 VPWR VGND sg13g2_decap_8
XFILLER_35_554 VPWR VGND sg13g2_fill_2
X_5802_ VGND VPWR _0387_ _0385_ net1407 sg13g2_or2_1
X_3994_ VPWR _0155_ _1552_ VGND sg13g2_inv_1
X_6782_ net104 VGND VPWR _0292_ s0.data_out\[0\]\[4\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_5733_ _0023_ _0321_ _0322_ _2765_ net1340 VPWR VGND sg13g2_a22oi_1
XFILLER_31_771 VPWR VGND sg13g2_decap_8
X_5664_ VGND VPWR net1313 _3055_ _3058_ _3057_ sg13g2_a21oi_1
X_5595_ _0008_ net399 _2996_ _2771_ net1340 VPWR VGND sg13g2_a22oi_1
X_4615_ net1370 _2040_ _2110_ VPWR VGND sg13g2_nor2_1
X_4546_ net1074 net1165 _2045_ VPWR VGND sg13g2_nor2b_1
X_4477_ _1930_ _1986_ net1479 _1987_ VPWR VGND sg13g2_nand3_1
X_3428_ VGND VPWR net1229 _1039_ _1042_ _1041_ sg13g2_a21oi_1
X_6216_ net1252 s0.data_out\[17\]\[4\] _0760_ VPWR VGND sg13g2_and2_1
X_6147_ _0696_ net1259 net689 VPWR VGND sg13g2_nand2_1
X_6078_ _0637_ VPWR _0638_ VGND _2755_ _0636_ sg13g2_o21ai_1
XFILLER_39_893 VPWR VGND sg13g2_fill_1
XFILLER_38_381 VPWR VGND sg13g2_fill_1
X_5029_ _2480_ net1009 _2479_ VPWR VGND sg13g2_nand2_1
XFILLER_26_554 VPWR VGND sg13g2_decap_4
XFILLER_14_716 VPWR VGND sg13g2_fill_2
XFILLER_10_966 VPWR VGND sg13g2_decap_8
XFILLER_1_653 VPWR VGND sg13g2_decap_8
XFILLER_0_141 VPWR VGND sg13g2_decap_8
XFILLER_0_152 VPWR VGND sg13g2_fill_2
XFILLER_49_646 VPWR VGND sg13g2_decap_8
XFILLER_45_874 VPWR VGND sg13g2_fill_1
XFILLER_44_340 VPWR VGND sg13g2_fill_1
XFILLER_44_384 VPWR VGND sg13g2_fill_2
X_4400_ s0.data_out\[7\]\[2\] s0.data_out\[6\]\[2\] net1092 _1911_ VPWR VGND sg13g2_mux2_1
X_5380_ VPWR _2798_ net436 VGND sg13g2_inv_1
X_4331_ s0.data_out\[8\]\[5\] s0.data_out\[7\]\[5\] net1108 _1854_ VPWR VGND sg13g2_mux2_1
X_4262_ net1125 VPWR _1789_ VGND _1728_ _1788_ sg13g2_o21ai_1
X_6001_ _0562_ net1271 net428 VPWR VGND sg13g2_nand2_1
X_4193_ net1116 net1145 _1728_ VPWR VGND sg13g2_nor2b_1
XFILLER_48_690 VPWR VGND sg13g2_decap_8
XFILLER_39_178 VPWR VGND sg13g2_decap_4
XFILLER_39_1024 VPWR VGND sg13g2_decap_4
XFILLER_36_896 VPWR VGND sg13g2_fill_1
XFILLER_35_373 VPWR VGND sg13g2_decap_4
X_6765_ net49 VGND VPWR _0275_ s0.shift_out\[1\][0] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_3977_ net1014 _2840_ _1539_ VPWR VGND sg13g2_nor2_1
X_5716_ net1007 _2781_ _0309_ VPWR VGND sg13g2_nor2_1
X_6696_ net137 VGND VPWR net454 s0.data_out\[7\]\[2\] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_5647_ net1303 net1162 _3041_ VPWR VGND sg13g2_nor2b_1
XFILLER_3_929 VPWR VGND sg13g2_decap_8
X_5578_ VGND VPWR _2984_ net1329 net335 sg13g2_or2_1
Xhold241 s0.data_out\[15\]\[7\] VPWR VGND net561 sg13g2_dlygate4sd3_1
Xhold230 s0.data_out\[13\]\[6\] VPWR VGND net550 sg13g2_dlygate4sd3_1
Xhold252 s0.data_out\[9\]\[1\] VPWR VGND net572 sg13g2_dlygate4sd3_1
X_4529_ _2028_ net997 _2027_ VPWR VGND sg13g2_nand2_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
Xhold285 s0.data_out\[1\]\[6\] VPWR VGND net605 sg13g2_dlygate4sd3_1
Xhold263 s0.data_out\[2\]\[4\] VPWR VGND net583 sg13g2_dlygate4sd3_1
XFILLER_6_8 VPWR VGND sg13g2_fill_2
Xhold274 _0023_ VPWR VGND net594 sg13g2_dlygate4sd3_1
Xhold296 s0.data_out\[12\]\[5\] VPWR VGND net616 sg13g2_dlygate4sd3_1
XFILLER_46_616 VPWR VGND sg13g2_fill_2
XFILLER_45_115 VPWR VGND sg13g2_fill_2
XFILLER_14_513 VPWR VGND sg13g2_fill_1
XFILLER_26_384 VPWR VGND sg13g2_decap_8
XFILLER_10_774 VPWR VGND sg13g2_decap_4
XFILLER_5_255 VPWR VGND sg13g2_decap_4
XFILLER_5_299 VPWR VGND sg13g2_fill_2
XFILLER_2_973 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_49_476 VPWR VGND sg13g2_decap_8
XFILLER_17_351 VPWR VGND sg13g2_fill_2
XFILLER_18_896 VPWR VGND sg13g2_fill_1
X_4880_ net1054 s0.data_out\[3\]\[6\] _2348_ VPWR VGND sg13g2_and2_1
X_3900_ _1466_ _2745_ net489 VPWR VGND sg13g2_nand2_1
X_3831_ VGND VPWR _1410_ _1409_ _1408_ sg13g2_or2_1
X_6550_ net295 VGND VPWR _0060_ s0.data_out\[19\]\[7\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3762_ _1339_ net1178 _1340_ _1341_ VPWR VGND sg13g2_a21o_1
XFILLER_32_376 VPWR VGND sg13g2_fill_1
X_5501_ net1325 _2905_ _2906_ _2907_ VPWR VGND sg13g2_nor3_1
X_6481_ VGND VPWR net1337 net1235 _0997_ net1229 sg13g2_a21oi_1
X_3693_ _1283_ net1198 net631 VPWR VGND sg13g2_nand2_1
X_5432_ VPWR _2850_ net670 VGND sg13g2_inv_1
X_5363_ VPWR _2781_ net519 VGND sg13g2_inv_1
X_4314_ _1837_ net627 net1120 VPWR VGND sg13g2_nand2b_1
X_5294_ VGND VPWR _2718_ _2719_ _0287_ _2720_ sg13g2_a21oi_1
X_4245_ net1375 _1715_ _1776_ VPWR VGND sg13g2_nor2_1
X_4176_ _1710_ VPWR _1711_ VGND net1119 _2844_ sg13g2_o21ai_1
XFILLER_27_115 VPWR VGND sg13g2_decap_4
XFILLER_36_660 VPWR VGND sg13g2_fill_1
X_6748_ net81 VGND VPWR _0258_ s0.data_out\[3\]\[6\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_6617__222 VPWR VGND net222 sg13g2_tiehi
X_6679_ net155 VGND VPWR _0189_ s0.valid_out\[8\][0] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_3_726 VPWR VGND sg13g2_decap_8
XFILLER_2_225 VPWR VGND sg13g2_decap_8
XFILLER_2_269 VPWR VGND sg13g2_fill_2
XFILLER_47_969 VPWR VGND sg13g2_decap_8
XFILLER_18_137 VPWR VGND sg13g2_decap_8
XFILLER_18_148 VPWR VGND sg13g2_fill_1
XFILLER_33_118 VPWR VGND sg13g2_decap_4
XFILLER_14_332 VPWR VGND sg13g2_fill_2
XFILLER_30_814 VPWR VGND sg13g2_decap_4
XFILLER_10_560 VPWR VGND sg13g2_decap_8
XFILLER_6_531 VPWR VGND sg13g2_decap_4
XFILLER_6_564 VPWR VGND sg13g2_fill_2
XFILLER_29_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_770 VPWR VGND sg13g2_decap_8
X_4030_ net1124 net1171 _1577_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_262 VPWR VGND sg13g2_fill_1
X_5981_ net1273 s0.data_out\[19\]\[6\] _0547_ VPWR VGND sg13g2_and2_1
X_4932_ _2395_ net1045 net512 VPWR VGND sg13g2_nand2_1
XFILLER_21_803 VPWR VGND sg13g2_fill_1
X_6602_ net238 VGND VPWR _0112_ s0.shift_out\[14\][0] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_4863_ net1060 VPWR _2335_ VGND _2253_ _2334_ sg13g2_o21ai_1
XFILLER_32_162 VPWR VGND sg13g2_fill_1
XFILLER_32_173 VPWR VGND sg13g2_decap_8
X_4794_ _2269_ net1060 _2268_ VPWR VGND sg13g2_nand2b_1
X_3814_ _1393_ net1188 net373 VPWR VGND sg13g2_nand2_1
X_6533_ net313 VGND VPWR net425 s0.data_out\[20\]\[2\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_3745_ net1207 VPWR _1327_ VGND _1260_ _1326_ sg13g2_o21ai_1
X_6464_ _0093_ _0982_ _0983_ _2810_ net1367 VPWR VGND sg13g2_a22oi_1
X_3676_ s0.data_out\[13\]\[6\] s0.data_out\[12\]\[6\] net1199 _1266_ VPWR VGND sg13g2_mux2_1
X_5415_ VPWR _2833_ net442 VGND sg13g2_inv_1
X_6395_ _0920_ s0.data_out\[15\]\[3\] net1248 VPWR VGND sg13g2_nand2b_1
X_5346_ VPWR _2764_ net438 VGND sg13g2_inv_1
X_5277_ net385 net1024 net1021 _2704_ VPWR VGND sg13g2_a21o_1
X_4228_ VGND VPWR _1763_ net1332 net336 sg13g2_or2_1
X_4159_ VGND VPWR _1694_ _1693_ net1446 sg13g2_or2_1
XFILLER_44_939 VPWR VGND sg13g2_decap_8
XFILLER_37_980 VPWR VGND sg13g2_decap_8
XFILLER_16_608 VPWR VGND sg13g2_fill_1
XFILLER_43_438 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_35_clk clknet_3_1__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_24_652 VPWR VGND sg13g2_fill_2
XFILLER_3_545 VPWR VGND sg13g2_decap_4
Xfanout1313 net1314 net1313 VPWR VGND sg13g2_buf_8
Xfanout1302 net347 net1302 VPWR VGND sg13g2_buf_2
XFILLER_3_589 VPWR VGND sg13g2_fill_1
Xfanout1324 net398 net1324 VPWR VGND sg13g2_buf_8
Xfanout1357 net1364 net1357 VPWR VGND sg13g2_buf_8
Xfanout1335 _2774_ net1335 VPWR VGND sg13g2_buf_8
Xfanout1346 net1350 net1346 VPWR VGND sg13g2_buf_8
Xfanout1368 net1369 net1368 VPWR VGND sg13g2_buf_1
Xfanout1379 net1383 net1379 VPWR VGND sg13g2_buf_8
XFILLER_47_766 VPWR VGND sg13g2_decap_8
XFILLER_46_287 VPWR VGND sg13g2_fill_2
X_6698__135 VPWR VGND net135 sg13g2_tiehi
XFILLER_36_81 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_26_clk clknet_3_6__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_15_696 VPWR VGND sg13g2_fill_1
XFILLER_30_611 VPWR VGND sg13g2_decap_8
XFILLER_30_622 VPWR VGND sg13g2_decap_4
X_3530_ net1201 net1172 _1132_ VPWR VGND sg13g2_nor2b_1
X_3461_ _1055_ _1072_ _1073_ _1074_ _1075_ VPWR VGND sg13g2_nor4_1
X_5200_ s0.data_out\[1\]\[5\] s0.data_out\[0\]\[5\] net1025 _2639_ VPWR VGND sg13g2_mux2_1
X_6180_ _0729_ net1257 net368 VPWR VGND sg13g2_nand2_1
X_3392_ net1213 net1164 _1006_ VPWR VGND sg13g2_nor2b_1
X_5131_ _0271_ _2572_ _2573_ _2880_ net1349 VPWR VGND sg13g2_a22oi_1
X_5062_ net1032 net1147 _2513_ VPWR VGND sg13g2_nor2b_1
XFILLER_42_1020 VPWR VGND sg13g2_decap_8
X_4013_ VGND VPWR net1390 net1334 _0161_ _1565_ sg13g2_a21oi_1
XFILLER_26_906 VPWR VGND sg13g2_fill_2
XFILLER_38_788 VPWR VGND sg13g2_fill_1
XFILLER_41_909 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_17_clk clknet_3_6__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
X_5964_ _0042_ _0533_ _0534_ _2790_ net1354 VPWR VGND sg13g2_a22oi_1
X_5895_ VGND VPWR net1294 _0465_ _0468_ _0467_ sg13g2_a21oi_1
X_4915_ s0.data_out\[3\]\[0\] s0.data_out\[2\]\[0\] net1043 _2378_ VPWR VGND sg13g2_mux2_1
XFILLER_33_460 VPWR VGND sg13g2_fill_1
X_4846_ VGND VPWR _2306_ _2308_ _2321_ net1428 sg13g2_a21oi_1
X_6516_ net35 VGND VPWR _0026_ s0.valid_out\[21\][0] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_4777_ s0.data_out\[4\]\[2\] s0.data_out\[3\]\[2\] net1057 _2252_ VPWR VGND sg13g2_mux2_1
XFILLER_10_1008 VPWR VGND sg13g2_decap_8
X_3728_ net1379 _1254_ _1314_ VPWR VGND sg13g2_nor2_1
X_6614__225 VPWR VGND net225 sg13g2_tiehi
X_6447_ _0970_ VPWR _0971_ VGND net1483 net662 sg13g2_o21ai_1
X_3659_ _1249_ net1197 net467 VPWR VGND sg13g2_nand2_1
X_6378_ net1226 net1168 _0903_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_537 VPWR VGND sg13g2_decap_8
X_5329_ _2747_ net1131 VPWR VGND sg13g2_inv_2
XFILLER_29_755 VPWR VGND sg13g2_decap_8
XFILLER_17_906 VPWR VGND sg13g2_decap_4
XFILLER_17_928 VPWR VGND sg13g2_fill_1
X_6621__218 VPWR VGND net218 sg13g2_tiehi
XFILLER_43_235 VPWR VGND sg13g2_fill_2
XFILLER_19_1000 VPWR VGND sg13g2_decap_8
XFILLER_25_994 VPWR VGND sg13g2_decap_8
XFILLER_40_953 VPWR VGND sg13g2_decap_8
XFILLER_24_493 VPWR VGND sg13g2_fill_2
XFILLER_11_143 VPWR VGND sg13g2_fill_1
XFILLER_11_176 VPWR VGND sg13g2_decap_8
XFILLER_4_810 VPWR VGND sg13g2_decap_8
XFILLER_22_72 VPWR VGND sg13g2_decap_8
XFILLER_4_887 VPWR VGND sg13g2_decap_8
Xfanout1121 s0.valid_out\[8\][0] net1121 VPWR VGND sg13g2_buf_8
Xfanout1132 net1133 net1132 VPWR VGND sg13g2_buf_8
Xfanout1110 net1112 net1110 VPWR VGND sg13g2_buf_8
Xfanout1165 s0.data_new_delayed\[2\] net1165 VPWR VGND sg13g2_buf_8
Xfanout1154 net1155 net1154 VPWR VGND sg13g2_buf_8
Xfanout1143 net1146 net1143 VPWR VGND sg13g2_buf_8
XFILLER_19_221 VPWR VGND sg13g2_fill_2
Xfanout1198 net1200 net1198 VPWR VGND sg13g2_buf_8
Xfanout1187 net1190 net1187 VPWR VGND sg13g2_buf_8
Xfanout1176 net1177 net1176 VPWR VGND sg13g2_buf_8
XFILLER_15_460 VPWR VGND sg13g2_fill_2
XFILLER_16_994 VPWR VGND sg13g2_decap_8
X_5680_ _3074_ net1314 _3073_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_964 VPWR VGND sg13g2_decap_8
X_4700_ net1062 net1157 _2187_ VPWR VGND sg13g2_nor2b_1
X_4631_ net1079 net488 _2122_ VPWR VGND sg13g2_and2_1
XFILLER_8_85 VPWR VGND sg13g2_decap_4
XFILLER_8_63 VPWR VGND sg13g2_fill_1
X_4562_ VGND VPWR _1949_ _2060_ _2061_ net1088 sg13g2_a21oi_1
X_4493_ net1097 VPWR _1999_ VGND _1967_ _1998_ sg13g2_o21ai_1
X_6301_ VGND VPWR _0729_ _0837_ _0838_ net1251 sg13g2_a21oi_1
X_3513_ net1485 net343 _0111_ VPWR VGND sg13g2_and2_1
XFILLER_6_191 VPWR VGND sg13g2_fill_2
X_6232_ _0072_ _0771_ _0772_ _2797_ net1365 VPWR VGND sg13g2_a22oi_1
X_3444_ _1056_ net1215 _1057_ _1058_ VPWR VGND sg13g2_a21o_1
Xclkbuf_leaf_6_clk clknet_3_3__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
XFILLER_40_0 VPWR VGND sg13g2_fill_1
X_6163_ s0.data_out\[18\]\[6\] s0.data_out\[17\]\[6\] net1258 _0712_ VPWR VGND sg13g2_mux2_1
X_5114_ VGND VPWR net1028 s0.data_out\[1\]\[4\] _2560_ _2522_ sg13g2_a21oi_1
X_6094_ net1278 VPWR _0650_ VGND _0615_ _0649_ sg13g2_o21ai_1
X_5045_ _2494_ net1028 _2495_ _2496_ VPWR VGND sg13g2_a21o_1
XFILLER_25_246 VPWR VGND sg13g2_decap_4
X_5947_ net1437 _0483_ _0520_ VPWR VGND sg13g2_nor2_1
XFILLER_25_279 VPWR VGND sg13g2_fill_2
X_5878_ VGND VPWR _0449_ _0452_ _0037_ _0453_ sg13g2_a21oi_1
XFILLER_21_441 VPWR VGND sg13g2_decap_8
X_4829_ s0.data_out\[4\]\[4\] s0.data_out\[3\]\[4\] net1057 _2304_ VPWR VGND sg13g2_mux2_1
XFILLER_1_835 VPWR VGND sg13g2_decap_8
XFILLER_0_323 VPWR VGND sg13g2_decap_8
XFILLER_49_828 VPWR VGND sg13g2_decap_8
X_6549__296 VPWR VGND net296 sg13g2_tiehi
XFILLER_29_530 VPWR VGND sg13g2_fill_2
XFILLER_29_552 VPWR VGND sg13g2_decap_8
XFILLER_44_522 VPWR VGND sg13g2_fill_1
XFILLER_1_1017 VPWR VGND sg13g2_decap_8
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
X_6695__138 VPWR VGND net138 sg13g2_tiehi
XFILLER_9_902 VPWR VGND sg13g2_fill_2
XFILLER_40_794 VPWR VGND sg13g2_fill_1
XFILLER_40_783 VPWR VGND sg13g2_decap_8
XFILLER_9_968 VPWR VGND sg13g2_decap_8
XFILLER_33_71 VPWR VGND sg13g2_fill_2
XFILLER_8_467 VPWR VGND sg13g2_fill_2
XFILLER_4_662 VPWR VGND sg13g2_decap_8
Xhold1 s0.genblk1\[4\].modules.bubble VPWR VGND net321 sg13g2_dlygate4sd3_1
XFILLER_48_872 VPWR VGND sg13g2_decap_8
XFILLER_35_533 VPWR VGND sg13g2_fill_1
XFILLER_35_577 VPWR VGND sg13g2_fill_2
X_5801_ _0386_ _0385_ net1407 _0378_ net1398 VPWR VGND sg13g2_a22oi_1
X_6781_ net117 VGND VPWR net403 s0.data_out\[0\]\[3\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_3993_ _1551_ VPWR _1552_ VGND net1491 net697 sg13g2_o21ai_1
X_5732_ net1340 _3064_ _0322_ VPWR VGND sg13g2_nor2_1
X_5663_ VGND VPWR _2943_ _3056_ _3057_ net1313 sg13g2_a21oi_1
X_5594_ net1340 net355 _2996_ VPWR VGND sg13g2_nor2_1
X_4614_ net1091 VPWR _2109_ VGND _2037_ _2108_ sg13g2_o21ai_1
X_6760__68 VPWR VGND net68 sg13g2_tiehi
X_4545_ s0.data_out\[6\]\[2\] s0.data_out\[5\]\[2\] net1081 _2044_ VPWR VGND sg13g2_mux2_1
X_4476_ net1096 VPWR _1986_ VGND _1926_ _1985_ sg13g2_o21ai_1
X_3427_ VGND VPWR _0932_ _1040_ _1041_ net1229 sg13g2_a21oi_1
X_6215_ _0068_ _0758_ _0759_ _2800_ net1357 VPWR VGND sg13g2_a22oi_1
X_6146_ _0679_ _0693_ _0694_ _0695_ VPWR VGND sg13g2_nor3_1
X_6077_ VGND VPWR net1003 _0581_ _0637_ net1355 sg13g2_a21oi_1
X_5028_ s0.data_out\[1\]\[0\] s0.data_out\[2\]\[0\] net1043 _2479_ VPWR VGND sg13g2_mux2_1
XFILLER_10_945 VPWR VGND sg13g2_decap_8
XFILLER_6_949 VPWR VGND sg13g2_decap_8
XFILLER_1_632 VPWR VGND sg13g2_decap_8
XFILLER_49_625 VPWR VGND sg13g2_decap_8
XFILLER_17_500 VPWR VGND sg13g2_fill_1
X_6562__282 VPWR VGND net282 sg13g2_tiehi
XFILLER_17_555 VPWR VGND sg13g2_decap_4
XFILLER_45_886 VPWR VGND sg13g2_decap_8
XFILLER_17_599 VPWR VGND sg13g2_decap_4
XFILLER_32_536 VPWR VGND sg13g2_decap_8
XFILLER_9_732 VPWR VGND sg13g2_decap_4
XFILLER_9_787 VPWR VGND sg13g2_fill_1
X_4330_ _1853_ net1107 net470 VPWR VGND sg13g2_nand2_1
XFILLER_5_42 VPWR VGND sg13g2_fill_2
X_4261_ net1000 _2848_ _1788_ VPWR VGND sg13g2_nor2_1
X_6000_ net1470 net337 _0051_ VPWR VGND sg13g2_and2_1
X_4192_ s0.data_out\[9\]\[7\] s0.data_out\[8\]\[7\] net1121 _1727_ VPWR VGND sg13g2_mux2_1
XFILLER_36_831 VPWR VGND sg13g2_fill_2
XFILLER_39_1003 VPWR VGND sg13g2_decap_8
X_6764_ net62 VGND VPWR _0274_ s0.genblk1\[19\].modules.bubble clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_23_569 VPWR VGND sg13g2_fill_2
X_3976_ _0151_ _1537_ _1538_ _2837_ net1385 VPWR VGND sg13g2_a22oi_1
X_5715_ VPWR _0019_ _0308_ VGND sg13g2_inv_1
X_6695_ net138 VGND VPWR net409 s0.data_out\[7\]\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_5646_ s0.data_out\[22\]\[2\] s0.data_out\[21\]\[2\] net1310 _3040_ VPWR VGND sg13g2_mux2_1
XFILLER_3_908 VPWR VGND sg13g2_decap_8
X_5577_ _2983_ net1390 net1464 VPWR VGND sg13g2_nand2_1
Xhold220 s0.data_out\[3\]\[0\] VPWR VGND net540 sg13g2_dlygate4sd3_1
Xhold242 _0108_ VPWR VGND net562 sg13g2_dlygate4sd3_1
Xhold231 _1325_ VPWR VGND net551 sg13g2_dlygate4sd3_1
Xhold253 _0181_ VPWR VGND net573 sg13g2_dlygate4sd3_1
X_4528_ net571 net692 net1092 _2027_ VPWR VGND sg13g2_mux2_1
X_4459_ _1970_ net1097 _1969_ VPWR VGND sg13g2_nand2b_1
Xhold264 _2563_ VPWR VGND net584 sg13g2_dlygate4sd3_1
Xhold275 s0.data_out\[12\]\[7\] VPWR VGND net595 sg13g2_dlygate4sd3_1
X_6497__56 VPWR VGND net56 sg13g2_tiehi
Xhold286 s0.data_out\[5\]\[2\] VPWR VGND net606 sg13g2_dlygate4sd3_1
Xhold297 _1438_ VPWR VGND net617 sg13g2_dlygate4sd3_1
X_6129_ VGND VPWR net1268 _0675_ _0678_ _0677_ sg13g2_a21oi_1
XFILLER_45_149 VPWR VGND sg13g2_fill_1
X_6546__299 VPWR VGND net299 sg13g2_tiehi
XFILLER_27_853 VPWR VGND sg13g2_decap_4
XFILLER_42_823 VPWR VGND sg13g2_decap_8
XFILLER_41_311 VPWR VGND sg13g2_fill_1
XFILLER_10_742 VPWR VGND sg13g2_fill_2
XFILLER_2_952 VPWR VGND sg13g2_decap_8
XFILLER_1_451 VPWR VGND sg13g2_decap_4
XFILLER_7_1023 VPWR VGND sg13g2_decap_4
XFILLER_39_81 VPWR VGND sg13g2_fill_1
XFILLER_39_70 VPWR VGND sg13g2_fill_1
XFILLER_44_160 VPWR VGND sg13g2_fill_1
X_3830_ VGND VPWR _1403_ _1405_ _1409_ net1423 sg13g2_a21oi_1
XFILLER_33_878 VPWR VGND sg13g2_fill_1
XFILLER_20_539 VPWR VGND sg13g2_fill_2
X_3761_ net1178 net1168 _1340_ VPWR VGND sg13g2_nor2b_1
XFILLER_9_551 VPWR VGND sg13g2_decap_8
X_5500_ net1328 s0.data_out\[22\]\[2\] _2906_ VPWR VGND sg13g2_nor2_1
X_6480_ _0994_ _0995_ _0996_ VPWR VGND sg13g2_nor2_1
X_3692_ _1279_ _1281_ net1423 _1282_ VPWR VGND sg13g2_nand3_1
X_5431_ VPWR _2849_ net687 VGND sg13g2_inv_1
X_5362_ VPWR _2780_ net650 VGND sg13g2_inv_1
X_4313_ _1834_ net1102 _1835_ _1836_ VPWR VGND sg13g2_a21o_1
X_5293_ VGND VPWR _2720_ net1329 net333 sg13g2_or2_1
X_6494__59 VPWR VGND net59 sg13g2_tiehi
X_4244_ net1123 VPWR _1775_ VGND _1712_ _1774_ sg13g2_o21ai_1
X_4175_ _1710_ net1119 net637 VPWR VGND sg13g2_nand2_1
XFILLER_23_322 VPWR VGND sg13g2_decap_4
XFILLER_24_823 VPWR VGND sg13g2_fill_2
XFILLER_24_856 VPWR VGND sg13g2_decap_8
X_6747_ net82 VGND VPWR _0257_ s0.data_out\[3\]\[5\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_23_399 VPWR VGND sg13g2_fill_1
X_3959_ _1503_ _1524_ _1525_ VPWR VGND sg13g2_nor2b_1
X_6678_ net157 VGND VPWR net359 s0.was_valid_out\[8\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5629_ VGND VPWR net1317 _3020_ _3023_ _3022_ sg13g2_a21oi_1
XFILLER_3_705 VPWR VGND sg13g2_decap_8
X_6552__292 VPWR VGND net292 sg13g2_tiehi
XFILLER_47_948 VPWR VGND sg13g2_decap_8
XFILLER_42_642 VPWR VGND sg13g2_fill_2
XFILLER_15_889 VPWR VGND sg13g2_fill_2
XFILLER_41_152 VPWR VGND sg13g2_fill_2
XFILLER_30_826 VPWR VGND sg13g2_fill_2
XFILLER_1_281 VPWR VGND sg13g2_fill_2
XFILLER_37_414 VPWR VGND sg13g2_fill_1
XFILLER_37_447 VPWR VGND sg13g2_fill_1
XFILLER_46_981 VPWR VGND sg13g2_decap_8
XFILLER_37_469 VPWR VGND sg13g2_fill_2
X_5980_ _0046_ _0545_ _0546_ _2786_ net1352 VPWR VGND sg13g2_a22oi_1
XFILLER_24_108 VPWR VGND sg13g2_decap_4
X_4931_ VPWR VGND net1438 _2386_ _2393_ net1444 _2394_ _2369_ sg13g2_a221oi_1
X_4862_ net1049 net434 _2334_ VPWR VGND sg13g2_and2_1
XFILLER_33_653 VPWR VGND sg13g2_fill_1
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
X_6601_ net239 VGND VPWR _0111_ s0.genblk1\[13\].modules.bubble clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_3813_ net1183 net1158 _1392_ VPWR VGND sg13g2_nor2b_1
X_4793_ VGND VPWR net1049 _2266_ _2268_ _2267_ sg13g2_a21oi_1
XFILLER_9_370 VPWR VGND sg13g2_fill_2
X_3744_ net1015 _2830_ _1326_ VPWR VGND sg13g2_nor2_1
X_6532_ net314 VGND VPWR net634 s0.data_out\[20\]\[1\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_6463_ net1367 _0950_ _0983_ VPWR VGND sg13g2_nor2_1
X_3675_ _1265_ net1199 net619 VPWR VGND sg13g2_nand2_1
X_5414_ VPWR _2832_ net467 VGND sg13g2_inv_1
X_6394_ _0917_ net1225 _0918_ _0919_ VPWR VGND sg13g2_a21o_1
XFILLER_0_719 VPWR VGND sg13g2_decap_8
X_5345_ VPWR _2763_ net377 VGND sg13g2_inv_1
X_5276_ _2703_ _2702_ net1436 _2696_ net1443 VPWR VGND sg13g2_a22oi_1
X_4227_ _1680_ _1760_ _1761_ _1762_ VPWR VGND sg13g2_nor3_1
XFILLER_29_904 VPWR VGND sg13g2_decap_8
XFILLER_28_436 VPWR VGND sg13g2_fill_2
XFILLER_29_959 VPWR VGND sg13g2_decap_8
X_4158_ VGND VPWR net1122 _1690_ _1693_ _1692_ sg13g2_a21oi_1
XFILLER_44_918 VPWR VGND sg13g2_decap_8
X_4089_ s0.data_out\[9\]\[5\] s0.data_out\[10\]\[5\] net1175 _1636_ VPWR VGND sg13g2_mux2_1
XFILLER_43_428 VPWR VGND sg13g2_fill_1
XFILLER_12_804 VPWR VGND sg13g2_fill_2
XFILLER_11_336 VPWR VGND sg13g2_fill_2
XFILLER_11_41 VPWR VGND sg13g2_fill_1
Xfanout1314 s0.shift_out\[22\][0] net1314 VPWR VGND sg13g2_buf_2
Xfanout1303 net1304 net1303 VPWR VGND sg13g2_buf_2
Xfanout1336 net1338 net1336 VPWR VGND sg13g2_buf_8
Xfanout1325 net1326 net1325 VPWR VGND sg13g2_buf_8
Xfanout1347 net1350 net1347 VPWR VGND sg13g2_buf_1
Xfanout1369 net1377 net1369 VPWR VGND sg13g2_buf_8
Xfanout1358 net1362 net1358 VPWR VGND sg13g2_buf_8
XFILLER_47_745 VPWR VGND sg13g2_decap_8
XFILLER_15_620 VPWR VGND sg13g2_decap_8
XFILLER_15_653 VPWR VGND sg13g2_decap_8
XFILLER_43_984 VPWR VGND sg13g2_decap_8
X_3460_ _1074_ _1070_ _1062_ VPWR VGND sg13g2_nand2b_1
XFILLER_42_4 VPWR VGND sg13g2_fill_1
X_3391_ s0.data_out\[15\]\[2\] s0.data_out\[14\]\[2\] net1219 _1005_ VPWR VGND sg13g2_mux2_1
X_5130_ net1349 _2510_ _2573_ VPWR VGND sg13g2_nor2_1
X_5061_ s0.data_out\[2\]\[6\] s0.data_out\[1\]\[6\] net1034 _2512_ VPWR VGND sg13g2_mux2_1
XFILLER_38_723 VPWR VGND sg13g2_decap_8
X_4012_ net1390 net1162 _1565_ VPWR VGND sg13g2_nor2_1
X_6607__233 VPWR VGND net233 sg13g2_tiehi
XFILLER_37_244 VPWR VGND sg13g2_fill_1
XFILLER_26_929 VPWR VGND sg13g2_decap_8
XFILLER_37_299 VPWR VGND sg13g2_decap_8
X_5963_ net1354 _0467_ _0534_ VPWR VGND sg13g2_nor2_1
X_4914_ VGND VPWR net1047 _2374_ _2377_ _2376_ sg13g2_a21oi_1
X_5894_ VGND VPWR _0336_ _0466_ _0467_ net1294 sg13g2_a21oi_1
XFILLER_34_984 VPWR VGND sg13g2_decap_8
X_4845_ _2318_ _2319_ _2320_ VPWR VGND sg13g2_nor2b_1
X_4776_ _2251_ net1056 net434 VPWR VGND sg13g2_nand2_1
X_6515_ net37 VGND VPWR _0025_ s0.was_valid_out\[21\][0] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3727_ net1209 VPWR _1313_ VGND _1251_ _1312_ sg13g2_o21ai_1
X_3658_ _1233_ VPWR _1248_ VGND net1454 _1240_ sg13g2_o21ai_1
X_6446_ _0913_ _0969_ net1477 _0970_ VPWR VGND sg13g2_nand3_1
X_6377_ _0901_ VPWR _0902_ VGND net1232 _2813_ sg13g2_o21ai_1
X_3589_ VGND VPWR net1201 s0.data_out\[13\]\[0\] _1190_ _1132_ sg13g2_a21oi_1
X_5328_ _2746_ net1138 VPWR VGND sg13g2_inv_2
XFILLER_0_516 VPWR VGND sg13g2_decap_8
X_5259_ net1489 net336 _0286_ VPWR VGND sg13g2_and2_1
XFILLER_29_767 VPWR VGND sg13g2_decap_8
XFILLER_28_288 VPWR VGND sg13g2_fill_1
XFILLER_25_973 VPWR VGND sg13g2_decap_8
XFILLER_40_932 VPWR VGND sg13g2_decap_8
XFILLER_4_866 VPWR VGND sg13g2_decap_8
Xfanout1100 net1101 net1100 VPWR VGND sg13g2_buf_8
XFILLER_26_1027 VPWR VGND sg13g2_fill_2
Xfanout1111 net1112 net1111 VPWR VGND sg13g2_buf_1
Xfanout1122 net1123 net1122 VPWR VGND sg13g2_buf_8
Xfanout1133 net1134 net1133 VPWR VGND sg13g2_buf_8
Xfanout1155 net708 net1155 VPWR VGND sg13g2_buf_8
Xfanout1144 net1146 net1144 VPWR VGND sg13g2_buf_8
Xfanout1177 s0.valid_out\[10\][0] net1177 VPWR VGND sg13g2_buf_8
Xfanout1166 net702 net1166 VPWR VGND sg13g2_buf_8
Xfanout1199 net1200 net1199 VPWR VGND sg13g2_buf_2
Xfanout1188 net1190 net1188 VPWR VGND sg13g2_buf_8
XFILLER_47_553 VPWR VGND sg13g2_decap_8
XFILLER_19_244 VPWR VGND sg13g2_decap_8
XFILLER_19_288 VPWR VGND sg13g2_fill_2
XFILLER_16_973 VPWR VGND sg13g2_decap_8
XFILLER_15_494 VPWR VGND sg13g2_fill_2
X_4630_ _0222_ _2120_ _2121_ _2861_ net1372 VPWR VGND sg13g2_a22oi_1
X_4561_ _2060_ s0.data_out\[5\]\[7\] net1094 VPWR VGND sg13g2_nand2b_1
X_6300_ _0837_ net475 net1258 VPWR VGND sg13g2_nand2b_1
X_3512_ net1381 _1110_ _0110_ VPWR VGND sg13g2_nor2_1
X_4492_ net1087 s0.data_out\[6\]\[4\] _1998_ VPWR VGND sg13g2_and2_1
X_6231_ net1365 _0709_ _0772_ VPWR VGND sg13g2_nor2_1
X_3443_ net1215 net1154 _1057_ VPWR VGND sg13g2_nor2b_1
X_6162_ _0711_ net1257 net664 VPWR VGND sg13g2_nand2_1
XFILLER_33_0 VPWR VGND sg13g2_decap_4
X_5113_ _0267_ _2558_ _2559_ _2882_ net1348 VPWR VGND sg13g2_a22oi_1
X_6093_ net1266 net440 _0649_ VPWR VGND sg13g2_and2_1
XFILLER_38_531 VPWR VGND sg13g2_decap_8
X_5044_ net1028 net1161 _2495_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_726 VPWR VGND sg13g2_decap_4
X_5946_ _0519_ _0518_ net1418 _0511_ net1427 VPWR VGND sg13g2_a22oi_1
X_5877_ net1472 VPWR _0453_ VGND net649 _0447_ sg13g2_o21ai_1
XFILLER_22_987 VPWR VGND sg13g2_decap_8
XFILLER_33_291 VPWR VGND sg13g2_decap_4
X_4828_ _2303_ net1056 net387 VPWR VGND sg13g2_nand2_1
X_4759_ net996 _2869_ _2238_ VPWR VGND sg13g2_nor2_1
X_6429_ s0.data_out\[16\]\[5\] s0.data_out\[15\]\[5\] net1233 _0954_ VPWR VGND sg13g2_mux2_1
X_6688__146 VPWR VGND net146 sg13g2_tiehi
XFILLER_1_814 VPWR VGND sg13g2_decap_8
XFILLER_49_807 VPWR VGND sg13g2_decap_8
XFILLER_12_431 VPWR VGND sg13g2_fill_2
XFILLER_12_453 VPWR VGND sg13g2_fill_1
XFILLER_13_987 VPWR VGND sg13g2_decap_8
XFILLER_24_291 VPWR VGND sg13g2_fill_2
XFILLER_9_947 VPWR VGND sg13g2_decap_8
XFILLER_32_1020 VPWR VGND sg13g2_decap_8
XFILLER_3_151 VPWR VGND sg13g2_decap_8
XFILLER_0_880 VPWR VGND sg13g2_decap_8
Xhold2 s0.genblk1\[17\].modules.bubble VPWR VGND net322 sg13g2_dlygate4sd3_1
XFILLER_48_851 VPWR VGND sg13g2_decap_8
XFILLER_35_523 VPWR VGND sg13g2_fill_2
XFILLER_35_556 VPWR VGND sg13g2_fill_1
X_6604__236 VPWR VGND net236 sg13g2_tiehi
X_3992_ _1550_ net1491 _1551_ VPWR VGND _1498_ sg13g2_nand3b_1
X_5800_ VGND VPWR net1301 _0382_ _0385_ _0384_ sg13g2_a21oi_1
X_6780_ net130 VGND VPWR _0290_ s0.data_out\[0\]\[2\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_5731_ net1313 VPWR _0321_ VGND _3061_ _0320_ sg13g2_o21ai_1
XFILLER_31_751 VPWR VGND sg13g2_fill_2
X_5662_ _3056_ s0.data_out\[21\]\[7\] net1318 VPWR VGND sg13g2_nand2b_1
X_5593_ net1326 VPWR _2995_ VGND _2935_ _2994_ sg13g2_o21ai_1
XFILLER_30_294 VPWR VGND sg13g2_decap_8
X_4613_ net1075 s0.data_out\[5\]\[3\] _2108_ VPWR VGND sg13g2_and2_1
X_4544_ _2043_ net1080 s0.data_out\[5\]\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_7_490 VPWR VGND sg13g2_fill_1
X_6214_ net1357 _0701_ _0759_ VPWR VGND sg13g2_nor2_1
X_6611__229 VPWR VGND net229 sg13g2_tiehi
X_4475_ net997 _2864_ _1985_ VPWR VGND sg13g2_nor2_1
X_3426_ _1040_ s0.data_out\[14\]\[7\] net1234 VPWR VGND sg13g2_nand2b_1
X_6145_ VPWR VGND _0692_ net1460 _0690_ net1452 _0694_ _0686_ sg13g2_a221oi_1
X_6076_ VGND VPWR net1265 s0.data_out\[18\]\[0\] _0636_ _0578_ sg13g2_a21oi_1
X_5027_ VGND VPWR net1038 _2475_ _2478_ _2477_ sg13g2_a21oi_1
XFILLER_14_718 VPWR VGND sg13g2_fill_1
X_5929_ VGND VPWR _0502_ _0492_ net1400 sg13g2_or2_1
XFILLER_16_1015 VPWR VGND sg13g2_decap_8
XFILLER_22_773 VPWR VGND sg13g2_fill_1
XFILLER_6_928 VPWR VGND sg13g2_decap_8
XFILLER_5_449 VPWR VGND sg13g2_fill_2
XFILLER_1_611 VPWR VGND sg13g2_decap_8
XFILLER_49_604 VPWR VGND sg13g2_decap_8
XFILLER_1_688 VPWR VGND sg13g2_decap_8
XFILLER_23_1008 VPWR VGND sg13g2_decap_8
XFILLER_28_83 VPWR VGND sg13g2_fill_1
XFILLER_45_843 VPWR VGND sg13g2_decap_8
XFILLER_44_386 VPWR VGND sg13g2_fill_1
XFILLER_13_740 VPWR VGND sg13g2_decap_8
XFILLER_40_581 VPWR VGND sg13g2_fill_1
XFILLER_13_784 VPWR VGND sg13g2_fill_1
XFILLER_5_983 VPWR VGND sg13g2_decap_8
X_4260_ _0186_ _1786_ _1787_ _2847_ net1384 VPWR VGND sg13g2_a22oi_1
X_4191_ _1726_ net1120 net371 VPWR VGND sg13g2_nand2_1
XFILLER_39_147 VPWR VGND sg13g2_fill_1
XFILLER_39_136 VPWR VGND sg13g2_fill_1
XFILLER_36_843 VPWR VGND sg13g2_fill_2
XFILLER_35_331 VPWR VGND sg13g2_decap_8
XFILLER_36_876 VPWR VGND sg13g2_decap_4
XFILLER_35_342 VPWR VGND sg13g2_fill_1
XFILLER_24_19 VPWR VGND sg13g2_decap_8
X_6763_ net64 VGND VPWR _0273_ s0.valid_out\[1\][0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3975_ net1385 _1459_ _1538_ VPWR VGND sg13g2_nor2_1
X_5714_ _0307_ VPWR _0308_ VGND net1463 net646 sg13g2_o21ai_1
X_6694_ net139 VGND VPWR _0204_ s0.data_out\[7\]\[0\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_5645_ net1435 _3038_ _3039_ VPWR VGND sg13g2_nor2_1
XFILLER_40_29 VPWR VGND sg13g2_fill_2
X_5576_ _2898_ _2980_ _2981_ _2982_ VPWR VGND sg13g2_nor3_1
Xhold210 s0.data_out\[15\]\[1\] VPWR VGND net530 sg13g2_dlygate4sd3_1
Xhold232 s0.was_valid_out\[7\][0] VPWR VGND net552 sg13g2_dlygate4sd3_1
Xhold243 s0.shift_out\[7\][0] VPWR VGND net563 sg13g2_dlygate4sd3_1
X_4527_ VGND VPWR net1085 _2023_ _2026_ _2025_ sg13g2_a21oi_1
Xhold221 s0.data_out\[1\]\[3\] VPWR VGND net541 sg13g2_dlygate4sd3_1
Xhold265 s0.shift_out\[3\][0] VPWR VGND net585 sg13g2_dlygate4sd3_1
Xhold287 s0.data_out\[15\]\[0\] VPWR VGND net607 sg13g2_dlygate4sd3_1
Xhold276 s0.data_out\[9\]\[0\] VPWR VGND net596 sg13g2_dlygate4sd3_1
Xhold254 s0.data_out\[3\]\[3\] VPWR VGND net574 sg13g2_dlygate4sd3_1
X_4458_ VGND VPWR net1087 _1968_ _1969_ _1967_ sg13g2_a21oi_1
XFILLER_49_49 VPWR VGND sg13g2_fill_2
X_6685__149 VPWR VGND net149 sg13g2_tiehi
X_3409_ s0.data_out\[14\]\[0\] s0.data_out\[15\]\[0\] net1232 _1023_ VPWR VGND sg13g2_mux2_1
Xhold298 s0.data_out\[11\]\[5\] VPWR VGND net618 sg13g2_dlygate4sd3_1
X_4389_ _1903_ _1902_ _1901_ VPWR VGND sg13g2_nand2b_1
X_6128_ VGND VPWR _0562_ _0676_ _0677_ net1268 sg13g2_a21oi_1
XFILLER_45_117 VPWR VGND sg13g2_fill_1
XFILLER_39_681 VPWR VGND sg13g2_fill_1
X_6059_ _0620_ net1272 s0.data_out\[18\]\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_26_320 VPWR VGND sg13g2_decap_4
XFILLER_42_846 VPWR VGND sg13g2_decap_8
XFILLER_42_879 VPWR VGND sg13g2_fill_2
XFILLER_10_710 VPWR VGND sg13g2_fill_1
XFILLER_14_41 VPWR VGND sg13g2_fill_1
XFILLER_14_63 VPWR VGND sg13g2_decap_8
XFILLER_14_96 VPWR VGND sg13g2_fill_2
XFILLER_22_581 VPWR VGND sg13g2_fill_2
XFILLER_5_202 VPWR VGND sg13g2_fill_2
XFILLER_2_931 VPWR VGND sg13g2_decap_8
XFILLER_30_84 VPWR VGND sg13g2_decap_4
XFILLER_7_1002 VPWR VGND sg13g2_decap_8
XFILLER_49_467 VPWR VGND sg13g2_decap_4
XFILLER_49_456 VPWR VGND sg13g2_decap_8
XFILLER_17_353 VPWR VGND sg13g2_fill_1
X_6601__239 VPWR VGND net239 sg13g2_tiehi
XFILLER_32_345 VPWR VGND sg13g2_fill_1
X_3760_ s0.data_out\[12\]\[1\] s0.data_out\[11\]\[1\] net1187 _1339_ VPWR VGND sg13g2_mux2_1
X_5430_ VPWR _2848_ net371 VGND sg13g2_inv_1
XFILLER_9_563 VPWR VGND sg13g2_decap_8
XFILLER_9_574 VPWR VGND sg13g2_fill_2
X_3691_ _1281_ _1280_ net1207 VPWR VGND sg13g2_nand2b_1
X_5361_ VPWR _2779_ net527 VGND sg13g2_inv_1
X_5292_ VGND VPWR net1399 _2716_ _2719_ net1393 sg13g2_a21oi_1
X_4312_ net1103 net1149 _1835_ VPWR VGND sg13g2_nor2b_1
X_4243_ net1000 _2851_ _1774_ VPWR VGND sg13g2_nor2_1
X_4174_ VPWR VGND _1707_ net1459 _1705_ net1455 _1709_ _1701_ sg13g2_a221oi_1
XFILLER_36_695 VPWR VGND sg13g2_decap_4
X_6746_ net83 VGND VPWR _0256_ s0.data_out\[3\]\[4\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_6691__142 VPWR VGND net142 sg13g2_tiehi
XFILLER_32_890 VPWR VGND sg13g2_fill_1
X_3958_ _1520_ VPWR _1524_ VGND _1510_ _1518_ sg13g2_o21ai_1
X_6677_ net158 VGND VPWR _0187_ s0.data_out\[9\]\[7\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_3889_ s0.data_out\[11\]\[2\] s0.data_out\[10\]\[2\] net1174 _1455_ VPWR VGND sg13g2_mux2_1
X_5628_ VGND VPWR _2915_ _3021_ _3022_ net1316 sg13g2_a21oi_1
X_5559_ _2963_ net1311 _2964_ _2965_ VPWR VGND sg13g2_a21o_1
XFILLER_47_927 VPWR VGND sg13g2_decap_8
X_6493__60 VPWR VGND net60 sg13g2_tiehi
XFILLER_42_621 VPWR VGND sg13g2_fill_1
XFILLER_42_610 VPWR VGND sg13g2_decap_8
XFILLER_26_172 VPWR VGND sg13g2_fill_2
XFILLER_41_131 VPWR VGND sg13g2_decap_8
X_6774__228 VPWR VGND net228 sg13g2_tiehi
XFILLER_41_164 VPWR VGND sg13g2_decap_8
XFILLER_14_367 VPWR VGND sg13g2_decap_8
XFILLER_10_551 VPWR VGND sg13g2_decap_4
XFILLER_41_61 VPWR VGND sg13g2_fill_2
XFILLER_37_7 VPWR VGND sg13g2_fill_1
XFILLER_38_905 VPWR VGND sg13g2_fill_1
XFILLER_49_297 VPWR VGND sg13g2_decap_4
XFILLER_38_949 VPWR VGND sg13g2_decap_8
XFILLER_2_99 VPWR VGND sg13g2_fill_1
XFILLER_46_960 VPWR VGND sg13g2_decap_8
XFILLER_17_150 VPWR VGND sg13g2_decap_4
X_4930_ VGND VPWR net1048 _2390_ _2393_ _2392_ sg13g2_a21oi_1
XFILLER_36_1007 VPWR VGND sg13g2_decap_8
X_4861_ _0241_ _2332_ _2333_ _2873_ net1359 VPWR VGND sg13g2_a22oi_1
XFILLER_33_632 VPWR VGND sg13g2_decap_8
X_6600_ net240 VGND VPWR _0110_ s0.valid_out\[14\][0] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_3812_ _1388_ _1389_ _1391_ VPWR VGND _1390_ sg13g2_nand3b_1
X_4792_ net1050 net1170 _2267_ VPWR VGND sg13g2_nor2b_1
X_3743_ VPWR _0131_ net551 VGND sg13g2_inv_1
X_6531_ net315 VGND VPWR _0041_ s0.data_out\[20\]\[0\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_6462_ net1240 VPWR _0982_ VGND _0947_ _0981_ sg13g2_o21ai_1
X_3674_ VGND VPWR net1207 _1261_ _1264_ _1263_ sg13g2_a21oi_1
X_6393_ net1226 net994 _0918_ VPWR VGND sg13g2_nor2_1
X_5413_ VPWR _2831_ net619 VGND sg13g2_inv_1
X_5344_ _2762_ net1066 VPWR VGND sg13g2_inv_2
X_5275_ VPWR _2702_ _2701_ VGND sg13g2_inv_1
X_4226_ _1733_ _1735_ _1761_ VPWR VGND sg13g2_nor2_1
XFILLER_28_404 VPWR VGND sg13g2_fill_1
X_4157_ VGND VPWR _1583_ _1691_ _1692_ net1122 sg13g2_a21oi_1
X_4088_ _1635_ net1138 _1634_ VPWR VGND sg13g2_nand2b_1
XFILLER_24_687 VPWR VGND sg13g2_fill_2
XFILLER_23_186 VPWR VGND sg13g2_fill_1
X_6729_ net101 VGND VPWR _0239_ s0.shift_out\[4\][0] clknet_leaf_13_clk sg13g2_dfrbpq_2
XFILLER_20_893 VPWR VGND sg13g2_fill_2
XFILLER_11_75 VPWR VGND sg13g2_decap_8
XFILLER_11_86 VPWR VGND sg13g2_fill_1
Xfanout1304 net1306 net1304 VPWR VGND sg13g2_buf_1
Xfanout1337 net1338 net1337 VPWR VGND sg13g2_buf_8
Xfanout1326 net398 net1326 VPWR VGND sg13g2_buf_8
Xfanout1315 net1317 net1315 VPWR VGND sg13g2_buf_8
Xfanout1348 net1350 net1348 VPWR VGND sg13g2_buf_8
Xfanout1359 net1362 net1359 VPWR VGND sg13g2_buf_1
XFILLER_47_724 VPWR VGND sg13g2_decap_8
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
XFILLER_19_437 VPWR VGND sg13g2_fill_2
XFILLER_43_963 VPWR VGND sg13g2_decap_8
XFILLER_42_451 VPWR VGND sg13g2_fill_2
XFILLER_42_484 VPWR VGND sg13g2_decap_4
XFILLER_7_886 VPWR VGND sg13g2_decap_8
XFILLER_6_352 VPWR VGND sg13g2_decap_4
XFILLER_7_897 VPWR VGND sg13g2_decap_8
X_3390_ _1004_ net1220 net548 VPWR VGND sg13g2_nand2_1
XFILLER_35_4 VPWR VGND sg13g2_fill_1
X_5060_ VGND VPWR net1039 _2508_ _2511_ _2510_ sg13g2_a21oi_1
X_4011_ net1166 net1450 net1390 _0160_ VPWR VGND sg13g2_mux2_1
XFILLER_26_908 VPWR VGND sg13g2_fill_1
XFILLER_26_919 VPWR VGND sg13g2_decap_4
XFILLER_37_278 VPWR VGND sg13g2_decap_4
X_5962_ net1294 VPWR _0533_ VGND _0464_ _0532_ sg13g2_o21ai_1
XFILLER_19_993 VPWR VGND sg13g2_decap_8
XFILLER_25_429 VPWR VGND sg13g2_decap_4
X_4913_ VGND VPWR _2259_ _2375_ _2376_ net1047 sg13g2_a21oi_1
XFILLER_34_963 VPWR VGND sg13g2_decap_8
X_5893_ _0466_ _2753_ s0.data_out\[19\]\[1\] VPWR VGND sg13g2_nand2_1
X_4844_ _2315_ _2317_ net1419 _2319_ VPWR VGND sg13g2_nand3_1
X_4775_ net1473 net340 _0238_ VPWR VGND sg13g2_and2_1
XFILLER_21_657 VPWR VGND sg13g2_decap_8
X_6514_ net38 VGND VPWR _0024_ s0.data_out\[22\]\[7\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_3726_ net1016 _2832_ _1312_ VPWR VGND sg13g2_nor2_1
X_3657_ VPWR VGND _1246_ net1459 _1244_ net1454 _1247_ _1240_ sg13g2_a221oi_1
X_6445_ net1243 VPWR _0969_ VGND _0909_ _0968_ sg13g2_o21ai_1
X_3588_ VGND VPWR _1186_ _1188_ _0112_ _1189_ sg13g2_a21oi_1
X_6376_ _0901_ net1232 net530 VPWR VGND sg13g2_nand2_1
X_5327_ _2745_ net1187 VPWR VGND sg13g2_inv_2
X_5258_ net1392 _2686_ _0285_ VPWR VGND sg13g2_nor2_1
X_5189_ _2625_ _2626_ _2624_ _2628_ VPWR VGND sg13g2_nand3_1
X_4209_ _1741_ _1743_ net1424 _1744_ VPWR VGND sg13g2_nand3_1
XFILLER_25_952 VPWR VGND sg13g2_decap_8
XFILLER_12_602 VPWR VGND sg13g2_decap_8
XFILLER_40_988 VPWR VGND sg13g2_decap_8
XFILLER_22_41 VPWR VGND sg13g2_decap_4
XFILLER_7_149 VPWR VGND sg13g2_decap_4
XFILLER_4_845 VPWR VGND sg13g2_decap_8
XFILLER_3_344 VPWR VGND sg13g2_fill_2
Xfanout1101 net1104 net1101 VPWR VGND sg13g2_buf_2
Xfanout1112 net1113 net1112 VPWR VGND sg13g2_buf_8
XFILLER_26_1006 VPWR VGND sg13g2_decap_8
Xfanout1134 s0.valid_out\[9\][0] net1134 VPWR VGND sg13g2_buf_8
Xfanout1123 net1127 net1123 VPWR VGND sg13g2_buf_8
Xfanout1156 net1160 net1156 VPWR VGND sg13g2_buf_8
Xfanout1145 net1146 net1145 VPWR VGND sg13g2_buf_8
Xfanout1167 s0.data_new_delayed\[1\] net1167 VPWR VGND sg13g2_buf_1
Xfanout1178 net1180 net1178 VPWR VGND sg13g2_buf_8
Xfanout1189 net1190 net1189 VPWR VGND sg13g2_buf_1
XFILLER_16_930 VPWR VGND sg13g2_fill_2
XFILLER_34_237 VPWR VGND sg13g2_decap_4
XFILLER_15_462 VPWR VGND sg13g2_fill_1
XFILLER_31_922 VPWR VGND sg13g2_fill_2
XFILLER_30_465 VPWR VGND sg13g2_decap_8
X_4560_ _2057_ net1078 _2058_ _2059_ VPWR VGND sg13g2_a21o_1
XFILLER_31_999 VPWR VGND sg13g2_decap_8
X_3511_ _1114_ _1115_ _0109_ VPWR VGND sg13g2_nor2_1
X_4491_ _0207_ _1996_ _1997_ _2857_ net1371 VPWR VGND sg13g2_a22oi_1
XFILLER_6_193 VPWR VGND sg13g2_fill_1
X_6230_ net1263 VPWR _0771_ VGND _0706_ _0770_ sg13g2_o21ai_1
X_3442_ s0.data_out\[15\]\[5\] s0.data_out\[14\]\[5\] net1219 _1056_ VPWR VGND sg13g2_mux2_1
X_6161_ VGND VPWR net1262 _0707_ _0710_ _0709_ sg13g2_a21oi_1
X_5112_ net1348 _2498_ _2559_ VPWR VGND sg13g2_nor2_1
X_6092_ _0056_ _0647_ _0648_ _2794_ net1355 VPWR VGND sg13g2_a22oi_1
X_5043_ s0.data_out\[2\]\[3\] s0.data_out\[1\]\[3\] net1035 _2494_ VPWR VGND sg13g2_mux2_1
XFILLER_43_29 VPWR VGND sg13g2_fill_1
X_5945_ VGND VPWR net1288 _0515_ _0518_ _0517_ sg13g2_a21oi_1
X_5876_ _0450_ _0451_ _0452_ VPWR VGND sg13g2_nor2_1
XFILLER_21_410 VPWR VGND sg13g2_decap_4
XFILLER_22_966 VPWR VGND sg13g2_decap_8
X_4827_ net1050 net1157 _2302_ VPWR VGND sg13g2_nor2b_1
X_4758_ _0234_ _2236_ _2237_ _2868_ net1363 VPWR VGND sg13g2_a22oi_1
XFILLER_5_609 VPWR VGND sg13g2_fill_1
X_4689_ _2176_ net1069 net492 VPWR VGND sg13g2_nand2_1
X_3709_ _1272_ _1274_ _1299_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_1017 VPWR VGND sg13g2_decap_8
X_6428_ _0953_ net1234 net430 VPWR VGND sg13g2_nand2_1
X_6359_ _0885_ _0886_ _0887_ VPWR VGND sg13g2_nor2_1
XFILLER_0_358 VPWR VGND sg13g2_decap_4
XFILLER_17_705 VPWR VGND sg13g2_decap_8
XFILLER_29_532 VPWR VGND sg13g2_fill_1
XFILLER_29_565 VPWR VGND sg13g2_fill_2
XFILLER_44_535 VPWR VGND sg13g2_decap_8
XFILLER_16_226 VPWR VGND sg13g2_fill_2
XFILLER_40_730 VPWR VGND sg13g2_fill_2
XFILLER_9_904 VPWR VGND sg13g2_fill_1
XFILLER_13_966 VPWR VGND sg13g2_decap_8
XFILLER_33_84 VPWR VGND sg13g2_fill_2
XFILLER_8_469 VPWR VGND sg13g2_fill_1
XFILLER_4_697 VPWR VGND sg13g2_decap_8
XFILLER_3_196 VPWR VGND sg13g2_fill_1
XFILLER_48_830 VPWR VGND sg13g2_decap_8
Xhold3 s0.genblk1\[15\].modules.bubble VPWR VGND net323 sg13g2_dlygate4sd3_1
X_3991_ net1184 VPWR _1550_ VGND _1495_ _1549_ sg13g2_o21ai_1
XFILLER_35_579 VPWR VGND sg13g2_fill_1
X_5730_ net1008 _2780_ _0320_ VPWR VGND sg13g2_nor2_1
XFILLER_16_793 VPWR VGND sg13g2_fill_1
X_5661_ _3053_ net1300 _3054_ _3055_ VPWR VGND sg13g2_a21o_1
X_5592_ net1011 _2770_ _2994_ VPWR VGND sg13g2_nor2_1
X_4612_ VPWR _0218_ _2107_ VGND sg13g2_inv_1
X_4543_ net1439 _2041_ _2042_ VPWR VGND sg13g2_nor2_1
X_4474_ VGND VPWR _1979_ _1983_ _0203_ _1984_ sg13g2_a21oi_1
X_6213_ net1267 VPWR _0758_ VGND _0698_ _0757_ sg13g2_o21ai_1
X_3425_ _1037_ net1217 _1038_ _1039_ VPWR VGND sg13g2_a21o_1
X_6144_ net1452 _0686_ _0693_ VPWR VGND sg13g2_nor2_1
X_6075_ net327 net1330 _0635_ _0052_ VPWR VGND sg13g2_nor3_1
XFILLER_38_340 VPWR VGND sg13g2_decap_4
X_5026_ VGND VPWR _2371_ _2476_ _2477_ net1038 sg13g2_a21oi_1
XFILLER_41_549 VPWR VGND sg13g2_fill_2
X_5928_ VPWR _0501_ _0500_ VGND sg13g2_inv_1
XFILLER_13_229 VPWR VGND sg13g2_decap_8
XFILLER_22_763 VPWR VGND sg13g2_fill_2
X_5859_ VPWR _0034_ _0437_ VGND sg13g2_inv_1
XFILLER_6_907 VPWR VGND sg13g2_decap_8
XFILLER_0_122 VPWR VGND sg13g2_fill_2
XFILLER_1_667 VPWR VGND sg13g2_decap_8
XFILLER_0_188 VPWR VGND sg13g2_decap_8
XFILLER_0_177 VPWR VGND sg13g2_decap_4
XFILLER_0_166 VPWR VGND sg13g2_fill_1
XFILLER_45_811 VPWR VGND sg13g2_fill_2
XFILLER_45_800 VPWR VGND sg13g2_decap_8
XFILLER_28_73 VPWR VGND sg13g2_decap_4
XFILLER_17_524 VPWR VGND sg13g2_decap_8
XFILLER_17_568 VPWR VGND sg13g2_fill_2
XFILLER_13_752 VPWR VGND sg13g2_fill_2
XFILLER_8_266 VPWR VGND sg13g2_decap_8
XFILLER_5_962 VPWR VGND sg13g2_decap_8
XFILLER_5_44 VPWR VGND sg13g2_fill_1
X_6610__230 VPWR VGND net230 sg13g2_tiehi
X_4190_ VGND VPWR net1126 _1722_ _1725_ _1724_ sg13g2_a21oi_1
XFILLER_39_159 VPWR VGND sg13g2_fill_2
XFILLER_36_833 VPWR VGND sg13g2_fill_1
XFILLER_23_505 VPWR VGND sg13g2_decap_8
XFILLER_23_516 VPWR VGND sg13g2_fill_1
X_6762_ net66 VGND VPWR net517 s0.was_valid_out\[1\][0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_6678__157 VPWR VGND net157 sg13g2_tiehi
X_3974_ net1181 VPWR _1537_ VGND _1456_ _1536_ sg13g2_o21ai_1
X_6693_ net140 VGND VPWR _0203_ s0.shift_out\[7\][0] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5713_ _3044_ _0306_ net1476 _0307_ VPWR VGND sg13g2_nand3_1
X_5644_ VGND VPWR net1316 _3035_ _3038_ _3037_ sg13g2_a21oi_1
X_5575_ _2956_ _2957_ _2981_ VPWR VGND sg13g2_nor2_1
Xhold200 _0032_ VPWR VGND net520 sg13g2_dlygate4sd3_1
Xhold211 _0102_ VPWR VGND net531 sg13g2_dlygate4sd3_1
Xhold244 s0.data_out\[22\]\[5\] VPWR VGND net564 sg13g2_dlygate4sd3_1
Xhold233 s0.data_out\[15\]\[3\] VPWR VGND net553 sg13g2_dlygate4sd3_1
X_4526_ VGND VPWR _1918_ _2024_ _2025_ net1085 sg13g2_a21oi_1
Xhold222 _2668_ VPWR VGND net542 sg13g2_dlygate4sd3_1
XFILLER_49_28 VPWR VGND sg13g2_decap_8
XFILLER_46_1009 VPWR VGND sg13g2_decap_8
Xhold266 s0.data_out\[22\]\[3\] VPWR VGND net586 sg13g2_dlygate4sd3_1
Xhold277 s0.data_out\[19\]\[0\] VPWR VGND net597 sg13g2_dlygate4sd3_1
Xhold255 _0255_ VPWR VGND net575 sg13g2_dlygate4sd3_1
X_4457_ s0.data_out\[7\]\[4\] s0.data_out\[6\]\[4\] net1092 _1968_ VPWR VGND sg13g2_mux2_1
Xhold288 s0.shift_out\[4\][0] VPWR VGND net608 sg13g2_dlygate4sd3_1
X_3408_ _1022_ net1228 _1021_ VPWR VGND sg13g2_nand2b_1
Xhold299 s0.data_out\[12\]\[6\] VPWR VGND net619 sg13g2_dlygate4sd3_1
X_4388_ _1902_ net1337 net1094 VPWR VGND sg13g2_nand2_1
X_6127_ _0676_ s0.data_out\[17\]\[2\] net1271 VPWR VGND sg13g2_nand2b_1
X_6058_ VGND VPWR net1278 _0616_ _0619_ _0618_ sg13g2_a21oi_1
X_5009_ net1039 VPWR _2463_ VGND net1392 net1030 sg13g2_o21ai_1
XFILLER_14_538 VPWR VGND sg13g2_decap_8
XFILLER_26_398 VPWR VGND sg13g2_fill_1
XFILLER_5_269 VPWR VGND sg13g2_fill_2
XFILLER_5_247 VPWR VGND sg13g2_decap_4
XFILLER_2_910 VPWR VGND sg13g2_decap_8
XFILLER_49_424 VPWR VGND sg13g2_fill_2
XFILLER_2_987 VPWR VGND sg13g2_decap_8
XFILLER_49_435 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_4
XFILLER_17_310 VPWR VGND sg13g2_decap_8
XFILLER_18_822 VPWR VGND sg13g2_fill_2
XFILLER_17_332 VPWR VGND sg13g2_fill_2
XFILLER_44_195 VPWR VGND sg13g2_fill_1
X_3690_ s0.data_out\[12\]\[5\] s0.data_out\[13\]\[5\] net1212 _1280_ VPWR VGND sg13g2_mux2_1
X_5360_ _2778_ net379 VPWR VGND sg13g2_inv_2
X_4311_ s0.data_out\[8\]\[6\] s0.data_out\[7\]\[6\] net1108 _1834_ VPWR VGND sg13g2_mux2_1
X_5291_ _2713_ _2710_ _2717_ _2718_ VPWR VGND sg13g2_a21o_1
X_4242_ _0182_ _1772_ _1773_ _2845_ net1376 VPWR VGND sg13g2_a22oi_1
X_4173_ _1694_ VPWR _1708_ VGND net1455 _1701_ sg13g2_o21ai_1
X_6684__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_36_674 VPWR VGND sg13g2_fill_1
X_3957_ _1523_ _1485_ _1522_ VPWR VGND sg13g2_nand2_1
X_6745_ net84 VGND VPWR net575 s0.data_out\[3\]\[3\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_6676_ net159 VGND VPWR net510 s0.data_out\[9\]\[6\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_3888_ net1490 net329 _0147_ VPWR VGND sg13g2_and2_1
XFILLER_13_1008 VPWR VGND sg13g2_decap_8
X_5627_ _3021_ net557 net1320 VPWR VGND sg13g2_nand2b_1
X_5558_ net1312 net1156 _2964_ VPWR VGND sg13g2_nor2b_1
X_4509_ _0211_ _2010_ _2011_ _2855_ net1373 VPWR VGND sg13g2_a22oi_1
X_5489_ _2896_ VPWR _2898_ VGND net1324 _2897_ sg13g2_o21ai_1
XFILLER_47_906 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_38_clk clknet_3_1__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_15_836 VPWR VGND sg13g2_decap_4
XFILLER_27_685 VPWR VGND sg13g2_fill_2
XFILLER_42_633 VPWR VGND sg13g2_fill_1
XFILLER_41_154 VPWR VGND sg13g2_fill_1
X_6600__240 VPWR VGND net240 sg13g2_tiehi
XFILLER_10_574 VPWR VGND sg13g2_fill_1
XFILLER_29_1015 VPWR VGND sg13g2_decap_8
X_6668__167 VPWR VGND net167 sg13g2_tiehi
XFILLER_2_784 VPWR VGND sg13g2_decap_8
XFILLER_49_221 VPWR VGND sg13g2_decap_4
XFILLER_37_405 VPWR VGND sg13g2_decap_8
XFILLER_2_45 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_29_clk clknet_3_5__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
X_4860_ net1358 _2264_ _2333_ VPWR VGND sg13g2_nor2_1
XFILLER_32_110 VPWR VGND sg13g2_fill_1
X_3811_ net1404 _1380_ _1390_ VPWR VGND sg13g2_nor2_1
X_6530_ net316 VGND VPWR _0040_ s0.shift_out\[20\][0] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_4791_ s0.data_out\[4\]\[0\] s0.data_out\[3\]\[0\] net1057 _2266_ VPWR VGND sg13g2_mux2_1
XFILLER_32_187 VPWR VGND sg13g2_fill_1
X_3742_ _1324_ VPWR _1325_ VGND net1486 net550 sg13g2_o21ai_1
X_6461_ net1223 s0.data_out\[15\]\[4\] _0981_ VPWR VGND sg13g2_and2_1
X_3673_ VGND VPWR _1148_ _1262_ _1263_ net1206 sg13g2_a21oi_1
X_6392_ _0916_ VPWR _0917_ VGND net1232 _2811_ sg13g2_o21ai_1
X_5412_ VPWR _2830_ net595 VGND sg13g2_inv_1
X_5343_ VPWR _2761_ net1088 VGND sg13g2_inv_1
X_5274_ VGND VPWR net1019 net993 _2701_ _2700_ sg13g2_a21oi_1
X_4225_ _1760_ _1733_ _1736_ _1759_ VPWR VGND sg13g2_and3_1
X_4156_ _1691_ s0.data_out\[8\]\[2\] net1131 VPWR VGND sg13g2_nand2b_1
XFILLER_46_29 VPWR VGND sg13g2_fill_1
X_4087_ VGND VPWR net1128 _1632_ _1634_ _1633_ sg13g2_a21oi_1
XFILLER_37_994 VPWR VGND sg13g2_decap_8
XFILLER_36_493 VPWR VGND sg13g2_fill_1
XFILLER_36_482 VPWR VGND sg13g2_fill_2
XFILLER_24_633 VPWR VGND sg13g2_decap_4
XFILLER_12_806 VPWR VGND sg13g2_fill_1
XFILLER_11_338 VPWR VGND sg13g2_fill_1
X_4989_ net1048 VPWR _2448_ VGND _2389_ _2447_ sg13g2_o21ai_1
X_6728_ net102 VGND VPWR _0238_ s0.genblk1\[3\].modules.bubble clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
XFILLER_11_349 VPWR VGND sg13g2_fill_2
X_6659_ net177 VGND VPWR net490 s0.data_out\[10\]\[1\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_3_537 VPWR VGND sg13g2_fill_1
XFILLER_3_559 VPWR VGND sg13g2_fill_2
XFILLER_11_98 VPWR VGND sg13g2_fill_2
Xfanout1305 net1306 net1305 VPWR VGND sg13g2_buf_8
Xfanout1338 _2743_ net1338 VPWR VGND sg13g2_buf_8
Xfanout1327 s0.valid_out\[23\][0] net1327 VPWR VGND sg13g2_buf_8
Xfanout1316 net1317 net1316 VPWR VGND sg13g2_buf_8
XFILLER_4_1006 VPWR VGND sg13g2_decap_8
Xfanout1349 net1350 net1349 VPWR VGND sg13g2_buf_2
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_28_983 VPWR VGND sg13g2_decap_8
XFILLER_43_942 VPWR VGND sg13g2_decap_8
XFILLER_15_644 VPWR VGND sg13g2_fill_2
XFILLER_7_810 VPWR VGND sg13g2_fill_1
XFILLER_10_382 VPWR VGND sg13g2_decap_8
XFILLER_2_570 VPWR VGND sg13g2_decap_8
XFILLER_38_703 VPWR VGND sg13g2_decap_4
X_4010_ net1170 net1458 net1391 _0159_ VPWR VGND sg13g2_mux2_1
XFILLER_28_4 VPWR VGND sg13g2_fill_2
X_6681__153 VPWR VGND net153 sg13g2_tiehi
XFILLER_38_747 VPWR VGND sg13g2_fill_2
XFILLER_38_769 VPWR VGND sg13g2_decap_4
X_5961_ net1003 _2796_ _0532_ VPWR VGND sg13g2_nor2_1
XFILLER_19_972 VPWR VGND sg13g2_decap_8
X_4912_ _2375_ s0.data_out\[2\]\[1\] net1056 VPWR VGND sg13g2_nand2b_1
XFILLER_34_942 VPWR VGND sg13g2_decap_8
X_5892_ _0463_ net1276 _0464_ _0465_ VPWR VGND sg13g2_a21o_1
X_4843_ VGND VPWR _2315_ _2317_ _2318_ net1419 sg13g2_a21oi_1
X_4774_ net1361 _2243_ _2244_ _0237_ VPWR VGND sg13g2_nor3_1
X_6513_ net39 VGND VPWR net594 s0.data_out\[22\]\[6\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_3725_ _0127_ _1310_ _1311_ _2828_ net1379 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_9_clk clknet_3_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_6444_ net1226 s0.data_out\[15\]\[0\] _0968_ VPWR VGND sg13g2_and2_1
X_3656_ _1246_ _1245_ net1201 VPWR VGND sg13g2_nand2b_1
X_3587_ VGND VPWR _1189_ net1332 net328 sg13g2_or2_1
X_6375_ VGND VPWR _0900_ _0899_ net1446 sg13g2_or2_1
X_5326_ _2744_ net1195 VPWR VGND sg13g2_inv_2
X_5257_ _2685_ _2686_ _0284_ VPWR VGND sg13g2_nor2_1
X_4208_ _1743_ _1742_ net1125 VPWR VGND sg13g2_nand2b_1
X_5188_ _2627_ _2624_ _2625_ _2626_ VPWR VGND sg13g2_and3_1
X_4139_ net1126 VPWR _1677_ VGND net1396 net1117 sg13g2_o21ai_1
XFILLER_28_268 VPWR VGND sg13g2_decap_4
XFILLER_19_1014 VPWR VGND sg13g2_decap_8
XFILLER_11_113 VPWR VGND sg13g2_fill_1
XFILLER_40_967 VPWR VGND sg13g2_decap_8
XFILLER_8_618 VPWR VGND sg13g2_decap_8
XFILLER_7_128 VPWR VGND sg13g2_fill_2
XFILLER_7_117 VPWR VGND sg13g2_fill_1
XFILLER_4_824 VPWR VGND sg13g2_decap_8
XFILLER_3_367 VPWR VGND sg13g2_fill_1
Xfanout1113 s0.shift_out\[8\][0] net1113 VPWR VGND sg13g2_buf_1
Xfanout1102 net1104 net1102 VPWR VGND sg13g2_buf_8
Xfanout1146 net707 net1146 VPWR VGND sg13g2_buf_8
Xfanout1135 net1136 net1135 VPWR VGND sg13g2_buf_8
Xfanout1124 net1127 net1124 VPWR VGND sg13g2_buf_8
Xfanout1168 net1169 net1168 VPWR VGND sg13g2_buf_8
Xfanout1157 net1160 net1157 VPWR VGND sg13g2_buf_8
Xfanout1179 net1180 net1179 VPWR VGND sg13g2_buf_1
XFILLER_47_50 VPWR VGND sg13g2_decap_8
XFILLER_19_235 VPWR VGND sg13g2_decap_4
XFILLER_42_260 VPWR VGND sg13g2_decap_4
XFILLER_15_496 VPWR VGND sg13g2_fill_1
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_30_400 VPWR VGND sg13g2_decap_8
XFILLER_30_444 VPWR VGND sg13g2_fill_2
XFILLER_31_978 VPWR VGND sg13g2_decap_8
X_6509__43 VPWR VGND net43 sg13g2_tiehi
X_3510_ net1485 VPWR _1115_ VGND net615 _1110_ sg13g2_o21ai_1
XFILLER_7_640 VPWR VGND sg13g2_fill_1
XFILLER_10_190 VPWR VGND sg13g2_fill_2
X_4490_ net1371 net390 _1997_ VPWR VGND sg13g2_nor2_1
X_3441_ _1051_ _1052_ _1050_ _1055_ VPWR VGND sg13g2_nand3_1
X_6160_ VGND VPWR _0594_ _0708_ _0709_ net1262 sg13g2_a21oi_1
X_5111_ net1038 VPWR _2558_ VGND _2495_ _2557_ sg13g2_o21ai_1
X_6091_ net1355 _0590_ _0648_ VPWR VGND sg13g2_nor2_1
X_5042_ _2493_ net1334 _2491_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_577 VPWR VGND sg13g2_fill_1
XFILLER_25_216 VPWR VGND sg13g2_fill_1
X_5944_ VGND VPWR _0398_ _0516_ _0517_ net1288 sg13g2_a21oi_1
XFILLER_34_761 VPWR VGND sg13g2_fill_2
X_5875_ VGND VPWR _2738_ _2753_ _0451_ net1288 sg13g2_a21oi_1
XFILLER_33_271 VPWR VGND sg13g2_decap_4
X_4826_ _2301_ _2297_ _2298_ _2300_ VPWR VGND sg13g2_and3_1
X_4757_ net1363 _2174_ _2237_ VPWR VGND sg13g2_nor2_1
X_4688_ VGND VPWR net1076 _2172_ _2175_ _2174_ sg13g2_a21oi_1
X_3708_ _1275_ _1297_ _1298_ VPWR VGND sg13g2_and2_1
X_6427_ _0952_ net1430 _0951_ VPWR VGND sg13g2_nand2_1
X_3639_ _1227_ net1193 _1228_ _1229_ VPWR VGND sg13g2_a21o_1
X_6729__101 VPWR VGND net101 sg13g2_tiehi
X_6358_ VGND VPWR net1337 net1247 _0886_ net1240 sg13g2_a21oi_1
X_5309_ net1466 net361 _2728_ VPWR VGND sg13g2_nor2_1
XFILLER_0_337 VPWR VGND sg13g2_fill_2
XFILLER_1_849 VPWR VGND sg13g2_decap_8
X_6289_ VGND VPWR net1250 _0823_ _0826_ _0825_ sg13g2_a21oi_1
XFILLER_17_728 VPWR VGND sg13g2_decap_4
XFILLER_16_238 VPWR VGND sg13g2_fill_2
XFILLER_17_739 VPWR VGND sg13g2_decap_4
XFILLER_40_742 VPWR VGND sg13g2_fill_2
XFILLER_33_41 VPWR VGND sg13g2_fill_2
X_6506__46 VPWR VGND net46 sg13g2_tiehi
XFILLER_4_676 VPWR VGND sg13g2_decap_8
Xhold4 s0.genblk1\[8\].modules.bubble VPWR VGND net324 sg13g2_dlygate4sd3_1
XFILLER_48_886 VPWR VGND sg13g2_decap_8
XFILLER_47_363 VPWR VGND sg13g2_fill_2
XFILLER_35_547 VPWR VGND sg13g2_decap_8
XFILLER_35_525 VPWR VGND sg13g2_fill_1
X_3990_ net1013 _2842_ _1549_ VPWR VGND sg13g2_nor2_1
X_5660_ net1300 net1142 _3054_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_753 VPWR VGND sg13g2_fill_1
X_4611_ _2106_ VPWR _2107_ VGND net1479 net682 sg13g2_o21ai_1
X_5591_ _0007_ _2992_ _2993_ _2773_ net1341 VPWR VGND sg13g2_a22oi_1
XFILLER_8_982 VPWR VGND sg13g2_decap_8
X_4542_ VGND VPWR net1087 _2038_ _2041_ _2040_ sg13g2_a21oi_1
X_4473_ VGND VPWR _1984_ net1331 net344 sg13g2_or2_1
X_3424_ net1217 net1145 _1038_ VPWR VGND sg13g2_nor2b_1
X_6212_ _2757_ _2805_ _0757_ VPWR VGND sg13g2_nor2_1
X_6143_ _0692_ _0691_ net1267 VPWR VGND sg13g2_nand2b_1
X_6074_ VPWR VGND _0612_ _0634_ _0633_ _0593_ _0635_ _0632_ sg13g2_a221oi_1
XFILLER_38_330 VPWR VGND sg13g2_decap_4
X_5025_ _2476_ net494 net1043 VPWR VGND sg13g2_nand2b_1
XFILLER_38_363 VPWR VGND sg13g2_fill_1
XFILLER_0_1020 VPWR VGND sg13g2_decap_8
X_5927_ _0500_ _0499_ net1409 _0492_ net1400 VPWR VGND sg13g2_a22oi_1
XFILLER_22_720 VPWR VGND sg13g2_fill_1
X_5858_ _0436_ VPWR _0437_ VGND net1462 net659 sg13g2_o21ai_1
X_4809_ s0.data_out\[4\]\[7\] s0.data_out\[3\]\[7\] net1059 _2284_ VPWR VGND sg13g2_mux2_1
X_5789_ net1286 net1142 _0374_ VPWR VGND sg13g2_nor2b_1
XFILLER_10_959 VPWR VGND sg13g2_decap_8
XFILLER_0_134 VPWR VGND sg13g2_decap_8
XFILLER_1_646 VPWR VGND sg13g2_decap_8
XFILLER_49_639 VPWR VGND sg13g2_decap_8
XFILLER_29_330 VPWR VGND sg13g2_fill_1
XFILLER_5_941 VPWR VGND sg13g2_decap_8
XFILLER_4_484 VPWR VGND sg13g2_fill_1
XFILLER_48_683 VPWR VGND sg13g2_decap_8
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_1017 VPWR VGND sg13g2_decap_8
X_6761_ net67 VGND VPWR net513 s0.data_out\[2\]\[7\] clknet_leaf_11_clk sg13g2_dfrbpq_2
XFILLER_35_388 VPWR VGND sg13g2_fill_2
X_5712_ net1316 VPWR _0306_ VGND _3041_ _0305_ sg13g2_o21ai_1
X_3973_ net1136 s0.data_out\[10\]\[2\] _1536_ VPWR VGND sg13g2_and2_1
X_6692_ net141 VGND VPWR _0202_ s0.genblk1\[6\].modules.bubble clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
XFILLER_31_561 VPWR VGND sg13g2_fill_2
X_5643_ VGND VPWR _2933_ _3036_ _3037_ net1316 sg13g2_a21oi_1
XFILLER_31_583 VPWR VGND sg13g2_fill_2
X_5574_ _2959_ _2974_ _2976_ _2980_ VPWR VGND sg13g2_nor3_1
XFILLER_8_790 VPWR VGND sg13g2_fill_1
X_4525_ _2024_ s0.data_out\[5\]\[1\] net1092 VPWR VGND sg13g2_nand2b_1
Xhold201 s0.data_out\[7\]\[0\] VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold223 s0.was_valid_out\[18\][0] VPWR VGND net543 sg13g2_dlygate4sd3_1
Xhold234 _0104_ VPWR VGND net554 sg13g2_dlygate4sd3_1
Xhold212 s0.data_out\[13\]\[3\] VPWR VGND net532 sg13g2_dlygate4sd3_1
Xhold256 s0.data_out\[2\]\[5\] VPWR VGND net576 sg13g2_dlygate4sd3_1
X_4456_ net1087 net1158 _1967_ VPWR VGND sg13g2_nor2b_1
Xhold245 _0319_ VPWR VGND net565 sg13g2_dlygate4sd3_1
Xhold267 _0020_ VPWR VGND net587 sg13g2_dlygate4sd3_1
Xhold278 _0639_ VPWR VGND net598 sg13g2_dlygate4sd3_1
X_4387_ net1100 VPWR _1901_ VGND net1394 net1089 sg13g2_o21ai_1
Xhold289 s0.data_out\[21\]\[4\] VPWR VGND net609 sg13g2_dlygate4sd3_1
X_3407_ VGND VPWR net1213 _1019_ _1021_ _1020_ sg13g2_a21oi_1
X_6126_ _0673_ net1252 _0674_ _0675_ VPWR VGND sg13g2_a21o_1
X_6057_ VGND VPWR _0505_ _0617_ _0618_ net1277 sg13g2_a21oi_1
X_5008_ _0259_ _2461_ _2462_ _2874_ net1348 VPWR VGND sg13g2_a22oi_1
XFILLER_26_333 VPWR VGND sg13g2_fill_1
XFILLER_26_344 VPWR VGND sg13g2_fill_1
XFILLER_26_377 VPWR VGND sg13g2_decap_8
XFILLER_5_204 VPWR VGND sg13g2_fill_1
XFILLER_10_767 VPWR VGND sg13g2_decap_8
XFILLER_10_778 VPWR VGND sg13g2_fill_1
XFILLER_5_237 VPWR VGND sg13g2_fill_1
XFILLER_10_789 VPWR VGND sg13g2_decap_4
XFILLER_5_259 VPWR VGND sg13g2_fill_1
XFILLER_2_966 VPWR VGND sg13g2_decap_8
XFILLER_39_95 VPWR VGND sg13g2_fill_2
X_4310_ _1833_ net1107 net627 VPWR VGND sg13g2_nand2_1
X_5290_ _2714_ VPWR _2717_ VGND net1399 _2716_ sg13g2_o21ai_1
X_4241_ net1376 _1692_ _1773_ VPWR VGND sg13g2_nor2_1
X_4172_ _1707_ _1706_ net1122 VPWR VGND sg13g2_nand2b_1
XFILLER_27_108 VPWR VGND sg13g2_decap_8
XFILLER_27_119 VPWR VGND sg13g2_fill_1
XFILLER_36_642 VPWR VGND sg13g2_fill_1
XFILLER_35_185 VPWR VGND sg13g2_fill_1
X_6744_ net85 VGND VPWR net435 s0.data_out\[3\]\[2\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_3956_ _1503_ _1510_ _1517_ _1521_ _1522_ VPWR VGND sg13g2_nor4_1
X_6675_ net160 VGND VPWR _0185_ s0.data_out\[9\]\[5\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_5626_ _3018_ net1303 _3019_ _3020_ VPWR VGND sg13g2_a21o_1
X_3887_ net1490 net341 _0146_ VPWR VGND sg13g2_and2_1
X_5557_ s0.data_out\[23\]\[4\] s0.data_out\[22\]\[4\] net1318 _2963_ VPWR VGND sg13g2_mux2_1
XFILLER_3_719 VPWR VGND sg13g2_decap_8
X_4508_ net1372 _1954_ _2011_ VPWR VGND sg13g2_nor2_1
XFILLER_2_218 VPWR VGND sg13g2_decap_8
X_5488_ net1392 _2750_ _2897_ VPWR VGND sg13g2_nor2_1
X_4439_ s0.data_out\[7\]\[7\] s0.data_out\[6\]\[7\] net1095 _1950_ VPWR VGND sg13g2_mux2_1
X_6109_ _0060_ _0660_ _0661_ _2791_ net1356 VPWR VGND sg13g2_a22oi_1
XFILLER_25_75 VPWR VGND sg13g2_decap_4
XFILLER_30_807 VPWR VGND sg13g2_decap_8
XFILLER_22_391 VPWR VGND sg13g2_fill_1
XFILLER_6_535 VPWR VGND sg13g2_fill_1
XFILLER_6_524 VPWR VGND sg13g2_decap_8
XFILLER_41_85 VPWR VGND sg13g2_decap_4
XFILLER_6_557 VPWR VGND sg13g2_decap_8
XFILLER_2_763 VPWR VGND sg13g2_decap_8
XFILLER_38_929 VPWR VGND sg13g2_fill_2
XFILLER_37_428 VPWR VGND sg13g2_decap_4
XFILLER_46_995 VPWR VGND sg13g2_decap_8
XFILLER_17_174 VPWR VGND sg13g2_fill_2
X_3810_ VGND VPWR _1389_ _1387_ net1413 sg13g2_or2_1
X_4790_ VGND VPWR net1060 _2262_ _2265_ _2264_ sg13g2_a21oi_1
X_3741_ _1323_ net1486 _1324_ VPWR VGND _1270_ sg13g2_nand3b_1
X_3672_ _1262_ s0.data_out\[12\]\[7\] net1212 VPWR VGND sg13g2_nand2b_1
X_6460_ _0092_ _0979_ _0980_ _2811_ net1369 VPWR VGND sg13g2_a22oi_1
X_6391_ _0916_ net1232 net553 VPWR VGND sg13g2_nand2_1
X_5411_ VPWR _2829_ net481 VGND sg13g2_inv_1
X_5342_ VPWR _2760_ net1107 VGND sg13g2_inv_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_5_590 VPWR VGND sg13g2_fill_1
X_5273_ VGND VPWR net1026 net402 _2700_ net1019 sg13g2_a21oi_1
X_4224_ _1744_ VPWR _1759_ VGND _1745_ _1753_ sg13g2_o21ai_1
XFILLER_29_918 VPWR VGND sg13g2_decap_4
X_4155_ _1688_ net1113 _1689_ _1690_ VPWR VGND sg13g2_a21o_1
X_4086_ net1128 net1153 _1633_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_973 VPWR VGND sg13g2_decap_8
XFILLER_23_100 VPWR VGND sg13g2_decap_4
XFILLER_23_111 VPWR VGND sg13g2_fill_1
X_6773__241 VPWR VGND net241 sg13g2_tiehi
X_4988_ net1009 _2882_ _2447_ VPWR VGND sg13g2_nor2_1
X_6727_ net103 VGND VPWR _0237_ s0.valid_out\[4\][0] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3939_ net1140 net1153 _1505_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_862 VPWR VGND sg13g2_decap_8
X_6658_ net178 VGND VPWR _0168_ s0.data_out\[10\]\[0\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_5609_ net1323 VPWR _3007_ VGND _2945_ _3006_ sg13g2_o21ai_1
X_6589_ net252 VGND VPWR _0099_ s0.genblk1\[14\].modules.bubble clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_3_549 VPWR VGND sg13g2_fill_1
Xfanout1339 net1340 net1339 VPWR VGND sg13g2_buf_8
Xfanout1306 net347 net1306 VPWR VGND sg13g2_buf_2
Xfanout1317 s0.shift_out\[22\][0] net1317 VPWR VGND sg13g2_buf_8
Xfanout1328 s0.valid_out\[23\][0] net1328 VPWR VGND sg13g2_buf_8
XFILLER_47_759 VPWR VGND sg13g2_decap_8
XFILLER_28_962 VPWR VGND sg13g2_decap_8
XFILLER_43_921 VPWR VGND sg13g2_decap_8
XFILLER_14_111 VPWR VGND sg13g2_fill_2
XFILLER_15_634 VPWR VGND sg13g2_fill_2
XFILLER_42_464 VPWR VGND sg13g2_fill_2
XFILLER_42_453 VPWR VGND sg13g2_fill_1
XFILLER_30_604 VPWR VGND sg13g2_decap_8
XFILLER_43_998 VPWR VGND sg13g2_decap_8
XFILLER_30_637 VPWR VGND sg13g2_fill_2
XFILLER_30_659 VPWR VGND sg13g2_decap_4
X_6674__161 VPWR VGND net161 sg13g2_tiehi
XFILLER_11_873 VPWR VGND sg13g2_fill_1
XFILLER_42_1013 VPWR VGND sg13g2_decap_8
XFILLER_38_737 VPWR VGND sg13g2_decap_4
X_5960_ VPWR _0041_ _0531_ VGND sg13g2_inv_1
XFILLER_46_792 VPWR VGND sg13g2_decap_8
X_5891_ net1277 net1166 _0464_ VPWR VGND sg13g2_nor2b_1
X_4911_ _2372_ net1036 _2373_ _2374_ VPWR VGND sg13g2_a21o_1
XFILLER_34_921 VPWR VGND sg13g2_decap_8
XFILLER_34_932 VPWR VGND sg13g2_fill_1
X_4842_ _2317_ net996 _2316_ VPWR VGND sg13g2_nand2_1
XFILLER_34_998 VPWR VGND sg13g2_decap_8
X_4773_ _0236_ net1473 _2246_ _2250_ VPWR VGND sg13g2_and3_1
X_6538__308 VPWR VGND net308 sg13g2_tiehi
X_6512_ net40 VGND VPWR _0022_ s0.data_out\[22\]\[5\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_3724_ net1379 _1231_ _1311_ VPWR VGND sg13g2_nor2_1
X_6443_ net326 net1331 _0967_ _0088_ VPWR VGND sg13g2_nor3_1
X_3655_ s0.data_out\[12\]\[0\] s0.data_out\[13\]\[0\] net1210 _1245_ VPWR VGND sg13g2_mux2_1
X_3586_ VPWR VGND _1187_ _1110_ _1166_ _1163_ _1188_ _1165_ sg13g2_a221oi_1
X_6374_ VGND VPWR net1242 _0896_ _0899_ _0898_ sg13g2_a21oi_1
X_5325_ VPWR _2743_ net1394 VGND sg13g2_inv_1
X_5256_ net1466 VPWR _2686_ VGND net1025 net1023 sg13g2_o21ai_1
X_4207_ _1631_ VPWR _1742_ VGND net1132 _2849_ sg13g2_o21ai_1
X_5187_ VGND VPWR _2626_ _2617_ net1399 sg13g2_or2_1
XFILLER_28_214 VPWR VGND sg13g2_fill_1
XFILLER_29_715 VPWR VGND sg13g2_fill_2
X_4138_ _0175_ _1675_ _1676_ _2841_ net1387 VPWR VGND sg13g2_a22oi_1
X_4069_ _1616_ net509 net1175 VPWR VGND sg13g2_nand2b_1
XFILLER_25_910 VPWR VGND sg13g2_decap_4
XFILLER_24_431 VPWR VGND sg13g2_decap_8
XFILLER_25_987 VPWR VGND sg13g2_decap_8
XFILLER_40_946 VPWR VGND sg13g2_decap_8
XFILLER_24_486 VPWR VGND sg13g2_decap_8
X_6658__178 VPWR VGND net178 sg13g2_tiehi
X_6518__33 VPWR VGND net33 sg13g2_tiehi
XFILLER_22_10 VPWR VGND sg13g2_decap_8
XFILLER_4_803 VPWR VGND sg13g2_decap_4
XFILLER_3_346 VPWR VGND sg13g2_fill_1
Xfanout1103 net1104 net1103 VPWR VGND sg13g2_buf_1
Xfanout1125 net1126 net1125 VPWR VGND sg13g2_buf_2
Xfanout1114 net1117 net1114 VPWR VGND sg13g2_buf_8
Xfanout1147 net1150 net1147 VPWR VGND sg13g2_buf_8
Xfanout1136 net1137 net1136 VPWR VGND sg13g2_buf_8
Xfanout1158 net1160 net1158 VPWR VGND sg13g2_buf_8
Xfanout1169 s0.data_new_delayed\[1\] net1169 VPWR VGND sg13g2_buf_8
XFILLER_15_453 VPWR VGND sg13g2_decap_8
XFILLER_16_987 VPWR VGND sg13g2_decap_8
XFILLER_31_957 VPWR VGND sg13g2_decap_8
XFILLER_8_89 VPWR VGND sg13g2_fill_1
XFILLER_6_173 VPWR VGND sg13g2_fill_1
X_3440_ _1054_ _1050_ _1051_ _1052_ VPWR VGND sg13g2_and3_1
XFILLER_3_880 VPWR VGND sg13g2_decap_8
X_6090_ net1279 VPWR _0647_ VGND _0587_ _0646_ sg13g2_o21ai_1
X_5110_ net1028 s0.data_out\[1\]\[3\] _2557_ VPWR VGND sg13g2_and2_1
X_5041_ VGND VPWR _2492_ _2491_ net1334 sg13g2_or2_1
XFILLER_38_545 VPWR VGND sg13g2_decap_4
X_6544__301 VPWR VGND net301 sg13g2_tiehi
XFILLER_25_239 VPWR VGND sg13g2_decap_8
X_5943_ _0516_ _2753_ net352 VPWR VGND sg13g2_nand2_1
X_5874_ net1273 _0444_ _0450_ VPWR VGND sg13g2_nor2_1
X_4825_ VGND VPWR _2300_ _2289_ net1401 sg13g2_or2_1
XFILLER_21_434 VPWR VGND sg13g2_decap_8
X_4756_ net1076 VPWR _2236_ VGND _2171_ _2235_ sg13g2_o21ai_1
X_4687_ VGND VPWR _2063_ _2173_ _2174_ net1076 sg13g2_a21oi_1
X_3707_ _1282_ VPWR _1297_ VGND _1290_ _1293_ sg13g2_o21ai_1
X_6426_ VGND VPWR net1240 _0948_ _0951_ _0950_ sg13g2_a21oi_1
X_3638_ net1193 net1165 _1228_ VPWR VGND sg13g2_nor2b_1
X_6357_ VGND VPWR net1337 net1233 _0885_ _0884_ sg13g2_a21oi_1
X_3569_ s0.data_out\[13\]\[5\] s0.data_out\[14\]\[5\] net1221 _1171_ VPWR VGND sg13g2_mux2_1
X_5308_ VGND VPWR net1466 _2712_ _0294_ _2727_ sg13g2_a21oi_1
XFILLER_0_316 VPWR VGND sg13g2_decap_8
XFILLER_1_828 VPWR VGND sg13g2_decap_8
X_6288_ VGND VPWR _0711_ _0824_ _0825_ net1250 sg13g2_a21oi_1
X_5239_ VPWR _0280_ _2672_ VGND sg13g2_inv_1
XFILLER_29_523 VPWR VGND sg13g2_decap_8
XFILLER_29_545 VPWR VGND sg13g2_decap_8
XFILLER_16_206 VPWR VGND sg13g2_decap_4
XFILLER_16_228 VPWR VGND sg13g2_fill_1
XFILLER_40_710 VPWR VGND sg13g2_fill_2
XFILLER_25_773 VPWR VGND sg13g2_decap_4
XFILLER_40_732 VPWR VGND sg13g2_fill_1
X_6671__164 VPWR VGND net164 sg13g2_tiehi
XFILLER_4_633 VPWR VGND sg13g2_fill_2
XFILLER_3_110 VPWR VGND sg13g2_fill_1
X_6782__104 VPWR VGND net104 sg13g2_tiehi
X_6528__318 VPWR VGND net318 sg13g2_tiehi
Xhold5 s0.genblk1\[1\].modules.bubble VPWR VGND net325 sg13g2_dlygate4sd3_1
XFILLER_0_894 VPWR VGND sg13g2_decap_8
XFILLER_12_8 VPWR VGND sg13g2_fill_1
XFILLER_48_865 VPWR VGND sg13g2_decap_8
X_4610_ _2105_ VPWR _2106_ VGND net997 _2104_ sg13g2_o21ai_1
X_5590_ net1341 _2907_ _2993_ VPWR VGND sg13g2_nor2_1
XFILLER_8_961 VPWR VGND sg13g2_decap_8
X_4541_ VGND VPWR _1934_ _2039_ _2040_ net1091 sg13g2_a21oi_1
X_4472_ _1904_ _1981_ _1982_ _1983_ VPWR VGND sg13g2_nor3_1
X_3423_ s0.data_out\[15\]\[7\] s0.data_out\[14\]\[7\] net1221 _1037_ VPWR VGND sg13g2_mux2_1
X_6211_ _0067_ _0755_ _0756_ _2801_ net1355 VPWR VGND sg13g2_a22oi_1
X_6142_ s0.data_out\[17\]\[0\] s0.data_out\[18\]\[0\] net1270 _0691_ VPWR VGND sg13g2_mux2_1
XFILLER_31_0 VPWR VGND sg13g2_fill_2
XFILLER_39_810 VPWR VGND sg13g2_fill_1
X_6073_ _0556_ VPWR _0634_ VGND _0608_ _0611_ sg13g2_o21ai_1
X_6648__188 VPWR VGND net188 sg13g2_tiehi
X_5024_ _2473_ net1027 _2474_ _2475_ VPWR VGND sg13g2_a21o_1
X_5926_ VGND VPWR net1287 _0496_ _0499_ _0498_ sg13g2_a21oi_1
X_5857_ _0435_ VPWR _0436_ VGND net1008 _0434_ sg13g2_o21ai_1
X_4808_ _2283_ net1058 net484 VPWR VGND sg13g2_nand2_1
X_5788_ s0.data_out\[21\]\[7\] s0.data_out\[20\]\[7\] net1296 _0373_ VPWR VGND sg13g2_mux2_1
XFILLER_10_938 VPWR VGND sg13g2_decap_8
X_4739_ _2222_ VPWR _2223_ VGND net1474 net606 sg13g2_o21ai_1
X_6409_ net1224 net1144 _0934_ VPWR VGND sg13g2_nor2b_1
XFILLER_1_625 VPWR VGND sg13g2_decap_8
XFILLER_49_618 VPWR VGND sg13g2_decap_8
XFILLER_45_879 VPWR VGND sg13g2_decap_8
XFILLER_45_857 VPWR VGND sg13g2_decap_4
XFILLER_17_548 VPWR VGND sg13g2_decap_8
XFILLER_9_736 VPWR VGND sg13g2_fill_2
XFILLER_5_920 VPWR VGND sg13g2_decap_8
XFILLER_5_997 VPWR VGND sg13g2_decap_8
XFILLER_0_691 VPWR VGND sg13g2_decap_8
XFILLER_48_662 VPWR VGND sg13g2_decap_8
X_6541__304 VPWR VGND net304 sg13g2_tiehi
XFILLER_35_356 VPWR VGND sg13g2_fill_2
X_6760_ net68 VGND VPWR net581 s0.data_out\[2\]\[6\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_5711_ net1304 s0.data_out\[21\]\[2\] _0305_ VPWR VGND sg13g2_and2_1
X_6719__112 VPWR VGND net112 sg13g2_tiehi
X_3972_ _0150_ _1534_ _1535_ _2838_ net1385 VPWR VGND sg13g2_a22oi_1
X_6691_ net142 VGND VPWR _0201_ s0.valid_out\[7\][0] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5642_ _3036_ net519 net1320 VPWR VGND sg13g2_nand2b_1
X_5573_ _2978_ VPWR _2979_ VGND _2930_ _2939_ sg13g2_o21ai_1
Xhold202 s0.data_out\[14\]\[4\] VPWR VGND net522 sg13g2_dlygate4sd3_1
X_4524_ _2021_ net1074 _2022_ _2023_ VPWR VGND sg13g2_a21o_1
Xhold235 s0.data_out\[7\]\[7\] VPWR VGND net555 sg13g2_dlygate4sd3_1
Xhold224 _0061_ VPWR VGND net544 sg13g2_dlygate4sd3_1
Xhold213 _0128_ VPWR VGND net533 sg13g2_dlygate4sd3_1
Xhold257 _2567_ VPWR VGND net577 sg13g2_dlygate4sd3_1
X_4455_ _1966_ net1421 _1965_ VPWR VGND sg13g2_nand2_1
Xhold246 s0.was_valid_out\[13\][0] VPWR VGND net566 sg13g2_dlygate4sd3_1
Xhold268 s0.data_out\[11\]\[1\] VPWR VGND net588 sg13g2_dlygate4sd3_1
X_4386_ _0199_ net556 _1900_ _2848_ net1375 VPWR VGND sg13g2_a22oi_1
Xhold279 s0.data_out\[16\]\[6\] VPWR VGND net599 sg13g2_dlygate4sd3_1
X_3406_ net1213 net1171 _1020_ VPWR VGND sg13g2_nor2b_1
X_6726__105 VPWR VGND net105 sg13g2_tiehi
X_6125_ net1252 net1165 _0674_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_651 VPWR VGND sg13g2_fill_2
X_6056_ _0617_ net440 net1284 VPWR VGND sg13g2_nand2b_1
XFILLER_22_1022 VPWR VGND sg13g2_decap_8
X_5007_ net1360 _2400_ _2462_ VPWR VGND sg13g2_nor2_1
X_5909_ VGND VPWR _0359_ _0481_ _0482_ net1293 sg13g2_a21oi_1
XFILLER_14_55 VPWR VGND sg13g2_decap_4
XFILLER_30_76 VPWR VGND sg13g2_fill_2
XFILLER_2_945 VPWR VGND sg13g2_decap_8
XFILLER_7_1016 VPWR VGND sg13g2_decap_8
XFILLER_49_426 VPWR VGND sg13g2_fill_1
XFILLER_7_1027 VPWR VGND sg13g2_fill_2
XFILLER_29_172 VPWR VGND sg13g2_fill_2
XFILLER_17_334 VPWR VGND sg13g2_fill_1
XFILLER_9_544 VPWR VGND sg13g2_decap_8
XFILLER_40_392 VPWR VGND sg13g2_decap_8
X_4240_ net1123 VPWR _1772_ VGND _1689_ _1771_ sg13g2_o21ai_1
X_4171_ _1578_ VPWR _1706_ VGND net1131 _2854_ sg13g2_o21ai_1
XFILLER_49_982 VPWR VGND sg13g2_decap_8
XFILLER_24_816 VPWR VGND sg13g2_decap_8
XFILLER_23_315 VPWR VGND sg13g2_decap_8
X_6743_ net86 VGND VPWR net401 s0.data_out\[3\]\[1\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_3955_ _1519_ _1520_ _1518_ _1521_ VPWR VGND sg13g2_nand3_1
X_6674_ net161 VGND VPWR _0184_ s0.data_out\[9\]\[4\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_5625_ net1303 net1166 _3019_ VPWR VGND sg13g2_nor2b_1
X_3886_ net1386 _1448_ _0145_ VPWR VGND sg13g2_nor2_1
X_5556_ net1324 _2960_ _2961_ _2962_ VPWR VGND sg13g2_nor3_1
X_4507_ net1100 VPWR _2010_ VGND _1951_ _2009_ sg13g2_o21ai_1
X_5487_ _2896_ _2895_ _2894_ VPWR VGND sg13g2_nand2b_1
X_4438_ _1949_ net1094 net404 VPWR VGND sg13g2_nand2_1
X_4369_ _0195_ _1886_ _1887_ _2851_ net1374 VPWR VGND sg13g2_a22oi_1
X_6108_ net1356 _0599_ _0661_ VPWR VGND sg13g2_nor2_1
X_6039_ VGND VPWR net1274 _0597_ _0600_ _0599_ sg13g2_a21oi_1
XFILLER_27_621 VPWR VGND sg13g2_fill_1
XFILLER_15_805 VPWR VGND sg13g2_fill_2
XFILLER_26_142 VPWR VGND sg13g2_decap_4
XFILLER_41_145 VPWR VGND sg13g2_fill_1
XFILLER_41_178 VPWR VGND sg13g2_fill_2
XFILLER_22_370 VPWR VGND sg13g2_fill_2
XFILLER_6_503 VPWR VGND sg13g2_fill_2
XFILLER_2_742 VPWR VGND sg13g2_decap_8
XFILLER_46_974 VPWR VGND sg13g2_decap_8
XFILLER_21_819 VPWR VGND sg13g2_fill_2
X_3740_ net1207 VPWR _1323_ VGND _1267_ _1322_ sg13g2_o21ai_1
XFILLER_20_307 VPWR VGND sg13g2_fill_2
XFILLER_32_167 VPWR VGND sg13g2_fill_2
X_6716__115 VPWR VGND net115 sg13g2_tiehi
XFILLER_9_341 VPWR VGND sg13g2_fill_1
XFILLER_12_1010 VPWR VGND sg13g2_decap_8
X_3671_ _1259_ net1194 _1260_ _1261_ VPWR VGND sg13g2_a21o_1
X_6390_ _0900_ VPWR _0915_ VGND net1456 _0907_ sg13g2_o21ai_1
X_5410_ VPWR _2828_ net457 VGND sg13g2_inv_1
X_5341_ _2759_ net1112 VPWR VGND sg13g2_inv_2
X_5272_ _2694_ _2697_ _2698_ _2699_ VPWR VGND sg13g2_or3_1
X_4223_ _1733_ _1736_ _1718_ _1758_ VPWR VGND _1757_ sg13g2_nand4_1
X_4154_ net1113 net1164 _1689_ VPWR VGND sg13g2_nor2b_1
X_6723__108 VPWR VGND net108 sg13g2_tiehi
X_4085_ s0.data_out\[10\]\[5\] s0.data_out\[9\]\[5\] net1134 _1632_ VPWR VGND sg13g2_mux2_1
XFILLER_28_418 VPWR VGND sg13g2_decap_4
XFILLER_28_429 VPWR VGND sg13g2_decap_8
XFILLER_37_952 VPWR VGND sg13g2_decap_8
XFILLER_36_484 VPWR VGND sg13g2_fill_1
X_6726_ net105 VGND VPWR _0236_ s0.was_valid_out\[4\][0] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4987_ _0254_ _2445_ _2446_ _2878_ net1358 VPWR VGND sg13g2_a22oi_1
X_3938_ s0.data_out\[11\]\[5\] s0.data_out\[10\]\[5\] net1176 _1504_ VPWR VGND sg13g2_mux2_1
X_6657_ net179 VGND VPWR _0167_ s0.shift_out\[10\][0] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3869_ net1381 _1386_ _1441_ VPWR VGND sg13g2_nor2_1
X_6588_ net253 VGND VPWR _0098_ s0.valid_out\[15\][0] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5608_ net1012 _2763_ _3006_ VPWR VGND sg13g2_nor2_1
X_5539_ net1311 net1142 _2945_ VPWR VGND sg13g2_nor2b_1
Xfanout1318 net1322 net1318 VPWR VGND sg13g2_buf_8
Xfanout1307 net1310 net1307 VPWR VGND sg13g2_buf_8
Xfanout1329 net1333 net1329 VPWR VGND sg13g2_buf_8
XFILLER_47_738 VPWR VGND sg13g2_decap_8
XFILLER_19_407 VPWR VGND sg13g2_decap_4
XFILLER_43_900 VPWR VGND sg13g2_decap_8
XFILLER_15_613 VPWR VGND sg13g2_decap_8
XFILLER_43_977 VPWR VGND sg13g2_decap_8
XFILLER_15_646 VPWR VGND sg13g2_fill_1
X_6784__78 VPWR VGND net78 sg13g2_tiehi
XFILLER_10_373 VPWR VGND sg13g2_decap_4
XFILLER_10_395 VPWR VGND sg13g2_decap_8
XFILLER_2_561 VPWR VGND sg13g2_decap_4
XFILLER_28_6 VPWR VGND sg13g2_fill_1
XFILLER_46_771 VPWR VGND sg13g2_decap_8
XFILLER_18_462 VPWR VGND sg13g2_decap_8
X_5890_ _0462_ VPWR _0463_ VGND net1283 _2790_ sg13g2_o21ai_1
X_4910_ net1036 net1167 _2373_ VPWR VGND sg13g2_nor2b_1
XFILLER_45_292 VPWR VGND sg13g2_fill_2
X_4841_ _2195_ VPWR _2316_ VGND net1069 _2875_ sg13g2_o21ai_1
XFILLER_34_977 VPWR VGND sg13g2_decap_8
X_4772_ _2248_ _2249_ _2247_ _2250_ VPWR VGND sg13g2_nand3_1
X_6511_ net41 VGND VPWR _0021_ s0.data_out\[22\]\[4\] clknet_leaf_0_clk sg13g2_dfrbpq_2
X_3723_ net1204 VPWR _1310_ VGND _1228_ _1309_ sg13g2_o21ai_1
X_6442_ VPWR VGND _0943_ _0966_ _0965_ _0924_ _0967_ _0964_ sg13g2_a221oi_1
X_3654_ _1244_ net1201 _1243_ VPWR VGND sg13g2_nand2b_1
X_3585_ _1173_ VPWR _1187_ VGND _1175_ _1183_ sg13g2_o21ai_1
X_6373_ VGND VPWR _0781_ _0897_ _0898_ net1242 sg13g2_a21oi_1
XFILLER_0_509 VPWR VGND sg13g2_decap_8
X_5324_ VPWR _2742_ net1471 VGND sg13g2_inv_1
X_5255_ VGND VPWR net427 net1001 _2685_ net1392 sg13g2_a21oi_1
X_4206_ _1741_ net1125 _1740_ VPWR VGND sg13g2_nand2b_1
X_5186_ VGND VPWR _2625_ _2623_ net1408 sg13g2_or2_1
X_4137_ net1386 _1610_ _1676_ VPWR VGND sg13g2_nor2_1
X_4068_ _1613_ net1128 _1614_ _1615_ VPWR VGND sg13g2_a21o_1
XFILLER_25_900 VPWR VGND sg13g2_fill_1
XFILLER_25_966 VPWR VGND sg13g2_decap_8
X_6709_ net123 VGND VPWR net448 s0.data_out\[6\]\[3\] clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_4_859 VPWR VGND sg13g2_decap_8
XFILLER_0_4 VPWR VGND sg13g2_decap_8
Xfanout1104 net563 net1104 VPWR VGND sg13g2_buf_8
Xfanout1115 net1117 net1115 VPWR VGND sg13g2_buf_1
Xfanout1126 net1127 net1126 VPWR VGND sg13g2_buf_8
Xfanout1137 net1141 net1137 VPWR VGND sg13g2_buf_8
XFILLER_47_513 VPWR VGND sg13g2_fill_2
XFILLER_19_204 VPWR VGND sg13g2_fill_2
Xfanout1148 net1150 net1148 VPWR VGND sg13g2_buf_8
Xfanout1159 net1160 net1159 VPWR VGND sg13g2_buf_8
XFILLER_16_966 VPWR VGND sg13g2_decap_8
XFILLER_42_240 VPWR VGND sg13g2_decap_8
XFILLER_7_631 VPWR VGND sg13g2_decap_8
XFILLER_6_163 VPWR VGND sg13g2_fill_1
XFILLER_2_380 VPWR VGND sg13g2_fill_2
X_5040_ _2490_ VPWR _2491_ VGND net1009 _2488_ sg13g2_o21ai_1
XFILLER_38_524 VPWR VGND sg13g2_decap_8
X_5942_ _0513_ net1273 _0514_ _0515_ VPWR VGND sg13g2_a21o_1
XFILLER_46_590 VPWR VGND sg13g2_fill_2
X_5873_ VGND VPWR _0449_ _0448_ _0446_ sg13g2_or2_1
X_4824_ net1401 _2289_ _2299_ VPWR VGND sg13g2_nor2_1
XFILLER_33_295 VPWR VGND sg13g2_fill_2
X_4755_ net996 _2870_ _2235_ VPWR VGND sg13g2_nor2_1
X_3706_ _1275_ _1295_ _1257_ _1296_ VPWR VGND sg13g2_nand3_1
X_4686_ _2173_ s0.data_out\[4\]\[6\] net1082 VPWR VGND sg13g2_nand2b_1
X_6515__37 VPWR VGND net37 sg13g2_tiehi
X_6425_ VGND VPWR _0842_ _0949_ _0950_ net1240 sg13g2_a21oi_1
X_3637_ s0.data_out\[13\]\[2\] s0.data_out\[12\]\[2\] net1200 _1227_ VPWR VGND sg13g2_mux2_1
X_6356_ net1240 VPWR _0884_ VGND net1394 net1223 sg13g2_o21ai_1
XFILLER_1_807 VPWR VGND sg13g2_decap_8
X_3568_ _1170_ net1218 _1169_ VPWR VGND sg13g2_nand2b_1
X_5307_ net1466 net394 _2727_ VPWR VGND sg13g2_nor2_1
XFILLER_0_306 VPWR VGND sg13g2_decap_4
X_6287_ _0824_ net599 net1257 VPWR VGND sg13g2_nand2b_1
X_3499_ net1380 _1041_ _1105_ VPWR VGND sg13g2_nor2_1
X_5238_ _2671_ VPWR _2672_ VGND net1467 net677 sg13g2_o21ai_1
X_6664__172 VPWR VGND net172 sg13g2_tiehi
X_5169_ net1005 _2607_ _2608_ VPWR VGND sg13g2_nor2_1
XFILLER_44_516 VPWR VGND sg13g2_fill_1
XFILLER_17_33 VPWR VGND sg13g2_fill_1
XFILLER_25_752 VPWR VGND sg13g2_decap_4
XFILLER_24_262 VPWR VGND sg13g2_fill_1
XFILLER_33_43 VPWR VGND sg13g2_fill_1
XFILLER_8_428 VPWR VGND sg13g2_decap_4
XFILLER_32_1013 VPWR VGND sg13g2_decap_8
XFILLER_4_612 VPWR VGND sg13g2_fill_2
XFILLER_3_144 VPWR VGND sg13g2_decap_8
XFILLER_3_177 VPWR VGND sg13g2_fill_2
XFILLER_0_873 VPWR VGND sg13g2_decap_8
XFILLER_48_844 VPWR VGND sg13g2_decap_8
XFILLER_47_321 VPWR VGND sg13g2_fill_1
Xhold6 s0.genblk1\[16\].modules.bubble VPWR VGND net326 sg13g2_dlygate4sd3_1
XFILLER_47_365 VPWR VGND sg13g2_fill_1
XFILLER_43_582 VPWR VGND sg13g2_fill_2
XFILLER_8_940 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_10_clk clknet_3_2__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_4540_ _2039_ s0.data_out\[5\]\[3\] net1093 VPWR VGND sg13g2_nand2b_1
X_4471_ _1956_ _1958_ _1982_ VPWR VGND sg13g2_nor2b_1
XFILLER_7_483 VPWR VGND sg13g2_decap_8
X_6210_ net1357 _0677_ _0756_ VPWR VGND sg13g2_nor2_1
X_3422_ _1036_ net1222 net612 VPWR VGND sg13g2_nand2_1
X_6141_ _0690_ net1267 _0689_ VPWR VGND sg13g2_nand2b_1
X_6072_ _0627_ _0630_ _0633_ VPWR VGND sg13g2_nor2_1
X_5023_ net1027 net1166 _2474_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_855 VPWR VGND sg13g2_fill_2
Xfanout1490 net1492 net1490 VPWR VGND sg13g2_buf_8
XFILLER_38_387 VPWR VGND sg13g2_fill_2
X_5925_ VGND VPWR _0379_ _0497_ _0498_ net1287 sg13g2_a21oi_1
XFILLER_22_700 VPWR VGND sg13g2_fill_1
XFILLER_22_711 VPWR VGND sg13g2_decap_8
X_5856_ VGND VPWR net1008 _0403_ _0435_ net1344 sg13g2_a21oi_1
XFILLER_16_1008 VPWR VGND sg13g2_decap_8
X_4807_ _2281_ VPWR _2282_ VGND _2272_ _2273_ sg13g2_o21ai_1
X_5787_ _0372_ net1296 net473 VPWR VGND sg13g2_nand2_1
X_4738_ _2154_ _2221_ net1474 _2222_ VPWR VGND sg13g2_nand3_1
X_4669_ _2156_ net1068 net444 VPWR VGND sg13g2_nand2_1
X_6408_ s0.data_out\[16\]\[7\] s0.data_out\[15\]\[7\] net1233 _0933_ VPWR VGND sg13g2_mux2_1
XFILLER_1_604 VPWR VGND sg13g2_decap_8
X_6339_ VGND VPWR net1002 _0846_ _0871_ net1365 sg13g2_a21oi_1
XFILLER_0_158 VPWR VGND sg13g2_fill_2
XFILLER_29_321 VPWR VGND sg13g2_decap_8
XFILLER_45_836 VPWR VGND sg13g2_decap_8
XFILLER_17_505 VPWR VGND sg13g2_fill_1
XFILLER_29_398 VPWR VGND sg13g2_decap_8
XFILLER_13_700 VPWR VGND sg13g2_fill_1
XFILLER_12_210 VPWR VGND sg13g2_fill_2
XFILLER_8_236 VPWR VGND sg13g2_fill_2
X_6534__312 VPWR VGND net312 sg13g2_tiehi
XFILLER_5_976 VPWR VGND sg13g2_decap_8
XFILLER_5_69 VPWR VGND sg13g2_fill_2
X_6502__51 VPWR VGND net51 sg13g2_tiehi
XFILLER_39_107 VPWR VGND sg13g2_decap_4
XFILLER_0_670 VPWR VGND sg13g2_decap_8
XFILLER_48_641 VPWR VGND sg13g2_decap_8
X_3971_ net1385 _1467_ _1535_ VPWR VGND sg13g2_nor2_1
X_5710_ _0018_ _0303_ _0304_ _2775_ net1342 VPWR VGND sg13g2_a22oi_1
X_6690_ net144 VGND VPWR _0200_ s0.was_valid_out\[7\][0] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5641_ _3033_ net1303 _3034_ _3035_ VPWR VGND sg13g2_a21o_1
X_5572_ _2959_ _2975_ _2976_ _2977_ _2978_ VPWR VGND sg13g2_nor4_1
X_6654__182 VPWR VGND net182 sg13g2_tiehi
X_4523_ net1074 net1169 _2022_ VPWR VGND sg13g2_nor2b_1
Xhold214 s0.data_out\[18\]\[6\] VPWR VGND net534 sg13g2_dlygate4sd3_1
Xhold225 s0.data_out\[14\]\[6\] VPWR VGND net545 sg13g2_dlygate4sd3_1
Xhold203 _1206_ VPWR VGND net523 sg13g2_dlygate4sd3_1
Xhold258 s0.data_out\[6\]\[6\] VPWR VGND net578 sg13g2_dlygate4sd3_1
Xhold236 _1899_ VPWR VGND net556 sg13g2_dlygate4sd3_1
X_4454_ VGND VPWR net1101 _1962_ _1965_ _1964_ sg13g2_a21oi_1
Xhold269 s0.data_out\[9\]\[3\] VPWR VGND net589 sg13g2_dlygate4sd3_1
Xhold247 _0121_ VPWR VGND net567 sg13g2_dlygate4sd3_1
X_4385_ net1375 _1845_ _1900_ VPWR VGND sg13g2_nor2_1
X_3405_ s0.data_out\[15\]\[0\] s0.data_out\[14\]\[0\] net1219 _1019_ VPWR VGND sg13g2_mux2_1
X_6124_ s0.data_out\[18\]\[2\] s0.data_out\[17\]\[2\] net1259 _0673_ VPWR VGND sg13g2_mux2_1
X_6055_ _0614_ net1266 _0615_ _0616_ VPWR VGND sg13g2_a21o_1
X_5006_ net1052 VPWR _2461_ VGND _2397_ _2460_ sg13g2_o21ai_1
XFILLER_22_1001 VPWR VGND sg13g2_decap_8
XFILLER_27_803 VPWR VGND sg13g2_decap_4
XFILLER_26_313 VPWR VGND sg13g2_decap_8
X_6661__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_26_324 VPWR VGND sg13g2_fill_1
X_5908_ _0481_ _2753_ s0.data_out\[19\]\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_34_390 VPWR VGND sg13g2_fill_2
XFILLER_10_725 VPWR VGND sg13g2_fill_2
X_5839_ net1345 _0341_ _0422_ VPWR VGND sg13g2_nor2_1
XFILLER_22_596 VPWR VGND sg13g2_fill_2
XFILLER_2_924 VPWR VGND sg13g2_decap_8
XFILLER_30_88 VPWR VGND sg13g2_fill_1
XFILLER_49_449 VPWR VGND sg13g2_decap_8
XFILLER_39_97 VPWR VGND sg13g2_fill_1
XFILLER_17_324 VPWR VGND sg13g2_fill_1
XFILLER_32_327 VPWR VGND sg13g2_fill_2
XFILLER_41_883 VPWR VGND sg13g2_fill_2
XFILLER_9_523 VPWR VGND sg13g2_fill_2
XFILLER_9_589 VPWR VGND sg13g2_decap_4
X_6638__199 VPWR VGND net199 sg13g2_tiehi
XFILLER_45_1012 VPWR VGND sg13g2_decap_8
X_4170_ _1705_ net1122 _1704_ VPWR VGND sg13g2_nand2b_1
XFILLER_49_961 VPWR VGND sg13g2_decap_8
XFILLER_36_688 VPWR VGND sg13g2_decap_8
XFILLER_36_699 VPWR VGND sg13g2_fill_2
XFILLER_16_390 VPWR VGND sg13g2_fill_1
X_6742_ net87 VGND VPWR _0252_ s0.data_out\[3\]\[0\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_3954_ _1507_ _1509_ net1424 _1520_ VPWR VGND sg13g2_nand3_1
X_6673_ net162 VGND VPWR net590 s0.data_out\[9\]\[3\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3885_ VGND VPWR _1450_ _1453_ _0144_ _1454_ sg13g2_a21oi_1
XFILLER_32_883 VPWR VGND sg13g2_fill_2
X_5624_ s0.data_out\[22\]\[1\] s0.data_out\[21\]\[1\] net1307 _3018_ VPWR VGND sg13g2_mux2_1
X_5555_ net1327 s0.data_out\[22\]\[4\] _2961_ VPWR VGND sg13g2_nor2_1
X_4506_ net998 _2860_ _2009_ VPWR VGND sg13g2_nor2_1
X_5486_ _2895_ net1336 net1318 VPWR VGND sg13g2_nand2_1
X_4437_ VGND VPWR net1100 _1945_ _1948_ _1947_ sg13g2_a21oi_1
X_4368_ net1374 _1829_ _1887_ VPWR VGND sg13g2_nor2_1
X_6107_ net1274 VPWR _0660_ VGND _0596_ _0659_ sg13g2_o21ai_1
X_4299_ VPWR VGND _1821_ net1459 _1819_ net1456 _1822_ _1814_ sg13g2_a221oi_1
XFILLER_39_460 VPWR VGND sg13g2_fill_2
X_6038_ VGND VPWR _0486_ _0598_ _0599_ net1274 sg13g2_a21oi_1
XFILLER_39_482 VPWR VGND sg13g2_decap_8
XFILLER_14_305 VPWR VGND sg13g2_fill_1
XFILLER_41_10 VPWR VGND sg13g2_decap_8
XFILLER_10_544 VPWR VGND sg13g2_decap_8
XFILLER_10_555 VPWR VGND sg13g2_fill_1
X_6531__315 VPWR VGND net315 sg13g2_tiehi
XFILLER_2_721 VPWR VGND sg13g2_decap_8
XFILLER_2_798 VPWR VGND sg13g2_decap_8
X_6709__123 VPWR VGND net123 sg13g2_tiehi
XFILLER_49_279 VPWR VGND sg13g2_decap_8
XFILLER_46_953 VPWR VGND sg13g2_decap_8
XFILLER_18_677 VPWR VGND sg13g2_fill_1
XFILLER_21_809 VPWR VGND sg13g2_fill_1
XFILLER_14_861 VPWR VGND sg13g2_fill_1
XFILLER_40_190 VPWR VGND sg13g2_decap_4
X_3670_ net1194 net1145 _1260_ VPWR VGND sg13g2_nor2b_1
X_5340_ VPWR _2758_ net1023 VGND sg13g2_inv_1
X_5271_ net1449 _2691_ _2698_ VPWR VGND sg13g2_nor2_1
X_6651__185 VPWR VGND net185 sg13g2_tiehi
X_4222_ _1754_ _1755_ _1756_ _1757_ VPWR VGND sg13g2_nor3_1
X_4153_ s0.data_out\[9\]\[2\] s0.data_out\[8\]\[2\] net1119 _1688_ VPWR VGND sg13g2_mux2_1
X_4084_ _1631_ net1132 s0.data_out\[9\]\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_36_430 VPWR VGND sg13g2_fill_2
XFILLER_24_658 VPWR VGND sg13g2_fill_1
X_4986_ net1358 _2368_ _2446_ VPWR VGND sg13g2_nor2_1
X_6725_ net106 VGND VPWR _0235_ s0.data_out\[5\]\[7\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_3937_ _1502_ _1500_ _1503_ VPWR VGND _1501_ sg13g2_nand3b_1
XFILLER_20_886 VPWR VGND sg13g2_decap_8
X_6656_ net180 VGND VPWR _0166_ s0.data_new_delayed\[7\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3868_ net1195 VPWR _1440_ VGND _1383_ _1439_ sg13g2_o21ai_1
X_6587_ net255 VGND VPWR net363 s0.was_valid_out\[15\][0] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_5607_ _0011_ _3004_ _3005_ _2766_ net1339 VPWR VGND sg13g2_a22oi_1
X_3799_ _1378_ net451 net1199 VPWR VGND sg13g2_nand2b_1
X_5538_ s0.data_out\[23\]\[7\] s0.data_out\[22\]\[7\] net1318 _2944_ VPWR VGND sg13g2_mux2_1
X_5469_ _2886_ VPWR net2 VGND _2778_ net992 sg13g2_o21ai_1
Xfanout1308 net1310 net1308 VPWR VGND sg13g2_buf_8
Xfanout1319 net1322 net1319 VPWR VGND sg13g2_buf_1
XFILLER_47_717 VPWR VGND sg13g2_decap_8
XFILLER_27_463 VPWR VGND sg13g2_fill_2
XFILLER_15_636 VPWR VGND sg13g2_fill_1
XFILLER_28_997 VPWR VGND sg13g2_decap_8
XFILLER_43_956 VPWR VGND sg13g2_decap_8
XFILLER_42_488 VPWR VGND sg13g2_fill_1
XFILLER_42_477 VPWR VGND sg13g2_decap_8
XFILLER_6_301 VPWR VGND sg13g2_fill_2
XFILLER_7_879 VPWR VGND sg13g2_decap_8
XFILLER_2_584 VPWR VGND sg13g2_decap_4
XFILLER_46_750 VPWR VGND sg13g2_decap_8
XFILLER_37_249 VPWR VGND sg13g2_decap_4
XFILLER_19_986 VPWR VGND sg13g2_decap_8
XFILLER_34_912 VPWR VGND sg13g2_decap_4
X_4840_ _2315_ net1064 _2314_ VPWR VGND sg13g2_nand2b_1
XFILLER_34_956 VPWR VGND sg13g2_decap_8
XFILLER_21_617 VPWR VGND sg13g2_decap_4
X_4771_ net996 VPWR _2249_ VGND net524 net1069 sg13g2_o21ai_1
XFILLER_14_691 VPWR VGND sg13g2_fill_1
X_6510_ net42 VGND VPWR net587 s0.data_out\[22\]\[3\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_6527__24 VPWR VGND net24 sg13g2_tiehi
X_3722_ net1193 s0.data_out\[12\]\[2\] _1309_ VPWR VGND sg13g2_and2_1
X_6441_ _0887_ VPWR _0966_ VGND _0939_ _0942_ sg13g2_o21ai_1
X_3653_ VGND VPWR net1192 _1241_ _1243_ _1242_ sg13g2_a21oi_1
X_6372_ _0897_ net420 net1248 VPWR VGND sg13g2_nand2b_1
X_5323_ _2741_ net1217 VPWR VGND sg13g2_inv_2
X_3584_ _1166_ _1185_ _1147_ _1186_ VPWR VGND sg13g2_nand3_1
X_5254_ VPWR _0283_ _2684_ VGND sg13g2_inv_1
X_5185_ _2624_ _2623_ net1408 _2617_ net1399 VPWR VGND sg13g2_a22oi_1
X_4205_ VGND VPWR net1116 _1738_ _1740_ _1739_ sg13g2_a21oi_1
X_4136_ net1139 VPWR _1675_ VGND _1607_ _1674_ sg13g2_o21ai_1
XFILLER_3_1020 VPWR VGND sg13g2_decap_8
XFILLER_44_709 VPWR VGND sg13g2_fill_2
X_4067_ net1129 net1149 _1614_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_271 VPWR VGND sg13g2_fill_1
XFILLER_24_400 VPWR VGND sg13g2_fill_2
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
X_4969_ _2419_ VPWR _2432_ VGND _2421_ _2428_ sg13g2_o21ai_1
XFILLER_7_109 VPWR VGND sg13g2_fill_2
X_6708_ net124 VGND VPWR _0218_ s0.data_out\[6\]\[2\] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_6639_ net198 VGND VPWR _0149_ s0.data_out\[11\]\[0\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_4_838 VPWR VGND sg13g2_decap_8
Xfanout1116 net1117 net1116 VPWR VGND sg13g2_buf_8
Xfanout1127 s0.shift_out\[9\][0] net1127 VPWR VGND sg13g2_buf_8
Xfanout1138 net1141 net1138 VPWR VGND sg13g2_buf_8
Xfanout1105 net1109 net1105 VPWR VGND sg13g2_buf_8
XFILLER_47_503 VPWR VGND sg13g2_fill_1
Xfanout1149 net1150 net1149 VPWR VGND sg13g2_buf_8
X_6706__126 VPWR VGND net126 sg13g2_tiehi
XFILLER_35_709 VPWR VGND sg13g2_fill_1
XFILLER_31_915 VPWR VGND sg13g2_decap_8
XFILLER_30_414 VPWR VGND sg13g2_decap_4
XFILLER_8_69 VPWR VGND sg13g2_fill_2
XFILLER_11_672 VPWR VGND sg13g2_decap_4
X_6713__119 VPWR VGND net119 sg13g2_tiehi
XFILLER_6_142 VPWR VGND sg13g2_decap_4
X_6524__27 VPWR VGND net27 sg13g2_tiehi
XFILLER_2_392 VPWR VGND sg13g2_fill_1
XFILLER_26_4 VPWR VGND sg13g2_fill_2
X_5941_ net1275 net1152 _0514_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_230 VPWR VGND sg13g2_fill_1
XFILLER_34_731 VPWR VGND sg13g2_decap_4
X_5872_ net366 net1281 _0448_ VPWR VGND sg13g2_nor2_1
X_4823_ VGND VPWR _2298_ _2296_ net1409 sg13g2_or2_1
XFILLER_22_959 VPWR VGND sg13g2_decap_8
XFILLER_34_797 VPWR VGND sg13g2_fill_2
X_4754_ VPWR _0233_ _2234_ VGND sg13g2_inv_1
X_3705_ _1291_ _1292_ _1293_ _1294_ _1295_ VPWR VGND sg13g2_nor4_1
X_4685_ _2170_ net1065 _2171_ _2172_ VPWR VGND sg13g2_a21o_1
X_6424_ _0949_ s0.data_out\[15\]\[4\] net1247 VPWR VGND sg13g2_nand2b_1
X_3636_ net1490 net342 _0123_ VPWR VGND sg13g2_and2_1
X_6355_ _0084_ _0882_ _0883_ _2803_ net1365 VPWR VGND sg13g2_a22oi_1
X_3567_ VGND VPWR net1205 _1167_ _1169_ _1168_ sg13g2_a21oi_1
X_5306_ VGND VPWR net1466 _2688_ _0293_ _2726_ sg13g2_a21oi_1
X_6286_ _0821_ net1237 _0822_ _0823_ VPWR VGND sg13g2_a21o_1
X_5237_ _2670_ VPWR _2671_ VGND net1005 _2669_ sg13g2_o21ai_1
X_3498_ net1229 VPWR _1104_ VGND _1038_ _1103_ sg13g2_o21ai_1
XFILLER_29_536 VPWR VGND sg13g2_decap_4
X_5168_ VGND VPWR net1021 _2605_ _2607_ _2606_ sg13g2_a21oi_1
X_5099_ _2548_ VPWR _2549_ VGND net1468 net663 sg13g2_o21ai_1
X_4119_ net1384 _1597_ _1662_ VPWR VGND sg13g2_nor2_1
XFILLER_44_528 VPWR VGND sg13g2_decap_8
XFILLER_17_78 VPWR VGND sg13g2_decap_4
XFILLER_13_959 VPWR VGND sg13g2_decap_8
XFILLER_21_992 VPWR VGND sg13g2_decap_8
XFILLER_3_167 VPWR VGND sg13g2_fill_1
XFILLER_3_189 VPWR VGND sg13g2_decap_8
XFILLER_0_852 VPWR VGND sg13g2_decap_8
XFILLER_48_823 VPWR VGND sg13g2_decap_8
Xhold7 s0.genblk1\[19\].modules.bubble VPWR VGND net327 sg13g2_dlygate4sd3_1
XFILLER_16_731 VPWR VGND sg13g2_decap_8
XFILLER_15_241 VPWR VGND sg13g2_decap_8
XFILLER_30_255 VPWR VGND sg13g2_fill_1
X_4470_ _1959_ _1980_ _1981_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_996 VPWR VGND sg13g2_decap_8
X_3421_ _1034_ VPWR _1035_ VGND _1025_ _1026_ sg13g2_o21ai_1
X_6140_ VGND VPWR net1252 _0687_ _0689_ _0688_ sg13g2_a21oi_1
XFILLER_31_2 VPWR VGND sg13g2_fill_1
X_6071_ _0612_ _0627_ _0629_ _0631_ _0632_ VPWR VGND sg13g2_and4_1
X_5022_ s0.data_out\[2\]\[1\] s0.data_out\[1\]\[1\] net1033 _2473_ VPWR VGND sg13g2_mux2_1
Xfanout1480 net1482 net1480 VPWR VGND sg13g2_buf_1
Xfanout1491 net1492 net1491 VPWR VGND sg13g2_buf_1
XFILLER_17_0 VPWR VGND sg13g2_fill_2
X_5924_ _0497_ s0.data_out\[19\]\[6\] net1296 VPWR VGND sg13g2_nand2b_1
X_5855_ VGND VPWR net1289 net468 _0434_ _0400_ sg13g2_a21oi_1
XFILLER_22_756 VPWR VGND sg13g2_decap_8
X_4806_ _2281_ _2280_ net1437 _2257_ net1444 VPWR VGND sg13g2_a22oi_1
X_5786_ _0368_ _0370_ _0371_ VPWR VGND sg13g2_nor2_1
X_4737_ net1072 VPWR _2221_ VGND _2150_ _2220_ sg13g2_o21ai_1
X_4668_ VGND VPWR _2152_ _2154_ _2155_ net1447 sg13g2_a21oi_1
X_6407_ _0932_ net1234 net561 VPWR VGND sg13g2_nand2_1
X_3619_ _0119_ _1212_ _1213_ _2820_ net1381 VPWR VGND sg13g2_a22oi_1
X_4599_ VGND VPWR _2092_ _2096_ _0215_ _2097_ sg13g2_a21oi_1
X_6338_ VGND VPWR net1237 net525 _0870_ _0841_ sg13g2_a21oi_1
XFILLER_0_115 VPWR VGND sg13g2_decap_8
X_6511__41 VPWR VGND net41 sg13g2_tiehi
XFILLER_0_148 VPWR VGND sg13g2_decap_4
X_6269_ net1238 net994 _0806_ VPWR VGND sg13g2_nor2_1
XFILLER_28_11 VPWR VGND sg13g2_decap_4
XFILLER_44_303 VPWR VGND sg13g2_fill_2
X_6703__129 VPWR VGND net129 sg13g2_tiehi
XFILLER_17_517 VPWR VGND sg13g2_decap_8
XFILLER_28_77 VPWR VGND sg13g2_fill_1
XFILLER_29_377 VPWR VGND sg13g2_fill_1
XFILLER_12_233 VPWR VGND sg13g2_fill_2
XFILLER_13_767 VPWR VGND sg13g2_fill_2
XFILLER_5_955 VPWR VGND sg13g2_decap_8
XFILLER_4_443 VPWR VGND sg13g2_fill_1
X_6647__190 VPWR VGND net190 sg13g2_tiehi
XFILLER_48_697 VPWR VGND sg13g2_decap_8
X_3970_ net1178 VPWR _1534_ VGND _1464_ _1533_ sg13g2_o21ai_1
XFILLER_15_1020 VPWR VGND sg13g2_decap_8
X_5640_ net1303 net1161 _3034_ VPWR VGND sg13g2_nor2b_1
X_5571_ _2974_ VPWR _2977_ VGND net1426 _2966_ sg13g2_o21ai_1
X_4522_ s0.data_out\[6\]\[1\] s0.data_out\[5\]\[1\] net1081 _2021_ VPWR VGND sg13g2_mux2_1
Xhold204 s0.was_valid_out\[3\][0] VPWR VGND net524 sg13g2_dlygate4sd3_1
X_4453_ VGND VPWR _1853_ _1963_ _1964_ net1101 sg13g2_a21oi_1
Xhold215 _0769_ VPWR VGND net535 sg13g2_dlygate4sd3_1
Xhold226 _0119_ VPWR VGND net546 sg13g2_dlygate4sd3_1
Xhold248 s0.data_out\[5\]\[5\] VPWR VGND net568 sg13g2_dlygate4sd3_1
Xhold259 s0.data_out\[1\]\[5\] VPWR VGND net579 sg13g2_dlygate4sd3_1
X_3404_ VGND VPWR net1227 _1015_ _1018_ _1017_ sg13g2_a21oi_1
Xhold237 s0.data_out\[21\]\[1\] VPWR VGND net557 sg13g2_dlygate4sd3_1
X_4384_ net1115 VPWR _1899_ VGND _1842_ _1898_ sg13g2_o21ai_1
X_6123_ _0672_ net1260 net511 VPWR VGND sg13g2_nand2_1
X_6054_ net1266 net1156 _0615_ VPWR VGND sg13g2_nor2b_1
X_5005_ net1010 _2880_ _2460_ VPWR VGND sg13g2_nor2_1
XFILLER_39_653 VPWR VGND sg13g2_fill_1
XFILLER_38_130 VPWR VGND sg13g2_decap_4
XFILLER_39_664 VPWR VGND sg13g2_decap_8
X_5907_ _0478_ net1276 _0479_ _0480_ VPWR VGND sg13g2_a21o_1
XFILLER_22_520 VPWR VGND sg13g2_decap_8
X_5838_ net1306 VPWR _0421_ VGND _0338_ _0420_ sg13g2_o21ai_1
X_5769_ s0.data_out\[20\]\[2\] s0.data_out\[21\]\[2\] net1309 _0354_ VPWR VGND sg13g2_mux2_1
XFILLER_30_12 VPWR VGND sg13g2_fill_1
XFILLER_2_903 VPWR VGND sg13g2_decap_8
XFILLER_30_78 VPWR VGND sg13g2_fill_1
XFILLER_39_32 VPWR VGND sg13g2_fill_2
XFILLER_39_21 VPWR VGND sg13g2_fill_2
XFILLER_39_54 VPWR VGND sg13g2_decap_4
XFILLER_44_122 VPWR VGND sg13g2_fill_2
XFILLER_45_667 VPWR VGND sg13g2_decap_4
XFILLER_26_881 VPWR VGND sg13g2_fill_1
XFILLER_13_520 VPWR VGND sg13g2_fill_2
XFILLER_25_391 VPWR VGND sg13g2_fill_2
XFILLER_9_502 VPWR VGND sg13g2_fill_1
XFILLER_49_940 VPWR VGND sg13g2_decap_8
XFILLER_35_111 VPWR VGND sg13g2_fill_2
X_6741_ net88 VGND VPWR _0251_ s0.shift_out\[3\][0] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_3953_ VGND VPWR _1519_ _1483_ net1441 sg13g2_or2_1
XFILLER_31_361 VPWR VGND sg13g2_decap_8
X_3884_ net1490 VPWR _1454_ VGND net644 _1448_ sg13g2_o21ai_1
X_6672_ net163 VGND VPWR net466 s0.data_out\[9\]\[2\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_5623_ _3017_ net1309 net557 VPWR VGND sg13g2_nand2_1
X_5554_ net416 net1327 _2960_ VPWR VGND sg13g2_nor2b_1
X_4505_ VPWR _0210_ _2008_ VGND sg13g2_inv_1
X_5485_ net1324 VPWR _2894_ VGND net1392 net1312 sg13g2_o21ai_1
X_4436_ VGND VPWR _1833_ _1946_ _1947_ net1100 sg13g2_a21oi_1
X_4367_ net1112 VPWR _1886_ VGND _1826_ _1885_ sg13g2_o21ai_1
X_6106_ net1261 net499 _0659_ VPWR VGND sg13g2_and2_1
X_4298_ _1821_ net1000 _1820_ VPWR VGND sg13g2_nand2_1
X_6037_ _0598_ net499 net1281 VPWR VGND sg13g2_nand2b_1
XFILLER_15_807 VPWR VGND sg13g2_fill_1
XFILLER_42_626 VPWR VGND sg13g2_decap_8
XFILLER_10_512 VPWR VGND sg13g2_fill_2
XFILLER_22_372 VPWR VGND sg13g2_fill_1
XFILLER_23_895 VPWR VGND sg13g2_fill_2
XFILLER_41_55 VPWR VGND sg13g2_fill_1
XFILLER_10_567 VPWR VGND sg13g2_decap_8
XFILLER_2_700 VPWR VGND sg13g2_decap_8
XFILLER_29_1008 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
XFILLER_2_777 VPWR VGND sg13g2_decap_8
XFILLER_49_225 VPWR VGND sg13g2_fill_2
XFILLER_49_258 VPWR VGND sg13g2_decap_4
XFILLER_46_932 VPWR VGND sg13g2_decap_8
X_6644__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_41_670 VPWR VGND sg13g2_decap_4
XFILLER_9_310 VPWR VGND sg13g2_fill_2
XFILLER_14_884 VPWR VGND sg13g2_decap_4
XFILLER_20_309 VPWR VGND sg13g2_fill_1
XFILLER_14_895 VPWR VGND sg13g2_fill_2
X_5270_ net1443 _2696_ _2697_ VPWR VGND sg13g2_nor2_1
X_4221_ _1756_ _1753_ _1745_ VPWR VGND sg13g2_nand2b_1
X_4152_ _1687_ net1118 net518 VPWR VGND sg13g2_nand2_1
X_4083_ _1627_ _1629_ net1433 _1630_ VPWR VGND sg13g2_nand3_1
XFILLER_37_987 VPWR VGND sg13g2_decap_8
XFILLER_36_464 VPWR VGND sg13g2_decap_4
XFILLER_24_637 VPWR VGND sg13g2_fill_2
X_4985_ net1047 VPWR _2445_ VGND _2365_ _2444_ sg13g2_o21ai_1
X_6724_ net107 VGND VPWR net450 s0.data_out\[5\]\[6\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_3936_ VGND VPWR _1502_ _1492_ net1405 sg13g2_or2_1
X_3867_ net1182 s0.data_out\[11\]\[6\] _1439_ VPWR VGND sg13g2_and2_1
X_6655_ net181 VGND VPWR _0165_ s0.data_new_delayed\[6\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_6586_ net256 VGND VPWR net504 s0.data_out\[16\]\[7\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_5606_ net1339 _2950_ _3005_ VPWR VGND sg13g2_nor2_1
X_3798_ _1375_ net1182 _1376_ _1377_ VPWR VGND sg13g2_a21o_1
X_5537_ _2943_ net1319 net377 VPWR VGND sg13g2_nand2_1
XFILLER_11_58 VPWR VGND sg13g2_fill_2
X_5468_ _2886_ net1458 net992 VPWR VGND sg13g2_nand2_1
X_5399_ VPWR _2817_ net420 VGND sg13g2_inv_1
Xfanout1309 net1310 net1309 VPWR VGND sg13g2_buf_8
X_4419_ _1930_ _1929_ net1096 VPWR VGND sg13g2_nand2b_1
XFILLER_46_239 VPWR VGND sg13g2_fill_1
XFILLER_46_217 VPWR VGND sg13g2_decap_8
XFILLER_28_976 VPWR VGND sg13g2_decap_8
XFILLER_43_935 VPWR VGND sg13g2_decap_8
XFILLER_42_401 VPWR VGND sg13g2_fill_1
XFILLER_36_77 VPWR VGND sg13g2_decap_4
X_6598__243 VPWR VGND net243 sg13g2_tiehi
XFILLER_35_1023 VPWR VGND sg13g2_decap_4
XFILLER_11_810 VPWR VGND sg13g2_fill_2
XFILLER_7_847 VPWR VGND sg13g2_fill_1
XFILLER_42_1027 VPWR VGND sg13g2_fill_2
XFILLER_38_707 VPWR VGND sg13g2_fill_1
XFILLER_45_261 VPWR VGND sg13g2_fill_2
X_4770_ VGND VPWR _2248_ _2241_ net1054 sg13g2_or2_1
XFILLER_20_139 VPWR VGND sg13g2_fill_1
X_6783__91 VPWR VGND net91 sg13g2_tiehi
X_3721_ _0126_ _1307_ _1308_ _2829_ net1378 VPWR VGND sg13g2_a22oi_1
X_6440_ _0961_ VPWR _0965_ VGND _0952_ _0960_ sg13g2_o21ai_1
X_3652_ net1191 net1171 _1242_ VPWR VGND sg13g2_nor2b_1
X_6371_ _0894_ net1225 _0895_ _0896_ VPWR VGND sg13g2_a21o_1
X_3583_ _1174_ _1175_ _1184_ _1185_ VPWR VGND sg13g2_nor3_1
X_5322_ _2740_ net1212 VPWR VGND sg13g2_inv_2
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_5253_ _2683_ VPWR _2684_ VGND net1467 net625 sg13g2_o21ai_1
X_5184_ _2621_ net1031 _2622_ _2623_ VPWR VGND sg13g2_a21o_1
X_4204_ net1116 net1154 _1739_ VPWR VGND sg13g2_nor2b_1
X_4135_ net1128 net505 _1674_ VPWR VGND sg13g2_and2_1
X_4066_ s0.data_out\[10\]\[6\] s0.data_out\[9\]\[6\] net1134 _1613_ VPWR VGND sg13g2_mux2_1
XFILLER_19_1007 VPWR VGND sg13g2_decap_8
X_6766__36 VPWR VGND net36 sg13g2_tiehi
X_4968_ _2394_ _2412_ _2420_ _2430_ _2431_ VPWR VGND sg13g2_or4_1
XFILLER_12_629 VPWR VGND sg13g2_fill_1
X_4899_ net1360 _2357_ _0249_ VPWR VGND sg13g2_nor2_1
X_6707_ net125 VGND VPWR net502 s0.data_out\[6\]\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3919_ _1484_ VPWR _1485_ VGND _1475_ _1476_ sg13g2_o21ai_1
XFILLER_20_684 VPWR VGND sg13g2_fill_2
XFILLER_22_35 VPWR VGND sg13g2_fill_1
X_6638_ net199 VGND VPWR _0148_ s0.shift_out\[11\][0] clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_4_817 VPWR VGND sg13g2_decap_8
XFILLER_22_79 VPWR VGND sg13g2_fill_1
X_6569_ net274 VGND VPWR _0079_ s0.data_out\[17\]\[2\] clknet_leaf_34_clk sg13g2_dfrbpq_2
Xfanout1117 s0.shift_out\[8\][0] net1117 VPWR VGND sg13g2_buf_8
Xfanout1128 net1129 net1128 VPWR VGND sg13g2_buf_2
Xfanout1106 net1109 net1106 VPWR VGND sg13g2_buf_1
Xfanout1139 net1141 net1139 VPWR VGND sg13g2_buf_1
XFILLER_47_43 VPWR VGND sg13g2_decap_8
XFILLER_47_32 VPWR VGND sg13g2_fill_2
XFILLER_19_239 VPWR VGND sg13g2_fill_2
XFILLER_28_751 VPWR VGND sg13g2_decap_4
X_6641__196 VPWR VGND net196 sg13g2_tiehi
XFILLER_43_798 VPWR VGND sg13g2_fill_2
XFILLER_7_600 VPWR VGND sg13g2_decap_4
XFILLER_7_611 VPWR VGND sg13g2_decap_4
XFILLER_3_894 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_fill_1
XFILLER_19_751 VPWR VGND sg13g2_fill_2
X_5940_ _0512_ VPWR _0513_ VGND net1281 _2786_ sg13g2_o21ai_1
XFILLER_18_250 VPWR VGND sg13g2_decap_8
XFILLER_18_272 VPWR VGND sg13g2_fill_2
XFILLER_19_795 VPWR VGND sg13g2_fill_1
X_5871_ _0446_ VPWR _0447_ VGND net1287 _0327_ sg13g2_o21ai_1
XFILLER_22_905 VPWR VGND sg13g2_fill_2
XFILLER_33_242 VPWR VGND sg13g2_decap_8
X_4822_ _2297_ _2296_ net1410 _2289_ net1401 VPWR VGND sg13g2_a22oi_1
XFILLER_33_275 VPWR VGND sg13g2_fill_2
X_4753_ _2233_ VPWR _2234_ VGND net1475 net568 sg13g2_o21ai_1
XFILLER_21_448 VPWR VGND sg13g2_fill_2
X_3704_ net1432 _1289_ _1294_ VPWR VGND sg13g2_nor2_1
XFILLER_30_982 VPWR VGND sg13g2_decap_8
X_4684_ net1065 net1148 _2171_ VPWR VGND sg13g2_nor2b_1
X_6423_ _0946_ net1223 _0947_ _0948_ VPWR VGND sg13g2_a21o_1
X_3635_ net1382 _1220_ _0122_ VPWR VGND sg13g2_nor2_1
X_6354_ net1365 _0818_ _0883_ VPWR VGND sg13g2_nor2_1
X_3566_ net1205 net1154 _1168_ VPWR VGND sg13g2_nor2b_1
X_5305_ net1466 net395 _2726_ VPWR VGND sg13g2_nor2_1
X_6285_ net1237 net1149 _0822_ VPWR VGND sg13g2_nor2b_1
X_3497_ net1017 _2819_ _1103_ VPWR VGND sg13g2_nor2_1
X_6588__253 VPWR VGND net253 sg13g2_tiehi
X_5236_ VGND VPWR net1005 _2629_ _2670_ net1347 sg13g2_a21oi_1
XFILLER_25_1022 VPWR VGND sg13g2_decap_8
X_5167_ net1020 net1161 _2606_ VPWR VGND sg13g2_nor2b_1
X_4118_ net1137 VPWR _1661_ VGND _1594_ _1660_ sg13g2_o21ai_1
X_5098_ _2547_ VPWR _2548_ VGND net1009 _2546_ sg13g2_o21ai_1
XFILLER_29_559 VPWR VGND sg13g2_fill_2
XFILLER_44_507 VPWR VGND sg13g2_fill_2
X_4049_ _1596_ s0.data_out\[9\]\[3\] net1177 VPWR VGND sg13g2_nand2b_1
XFILLER_17_24 VPWR VGND sg13g2_fill_2
X_6595__246 VPWR VGND net246 sg13g2_tiehi
XFILLER_21_971 VPWR VGND sg13g2_decap_8
XFILLER_33_78 VPWR VGND sg13g2_fill_1
XFILLER_33_89 VPWR VGND sg13g2_fill_1
XFILLER_20_470 VPWR VGND sg13g2_decap_8
X_6712__120 VPWR VGND net120 sg13g2_tiehi
XFILLER_4_614 VPWR VGND sg13g2_fill_1
XFILLER_4_669 VPWR VGND sg13g2_decap_8
XFILLER_0_831 VPWR VGND sg13g2_decap_8
XFILLER_48_802 VPWR VGND sg13g2_decap_8
Xhold8 s0.genblk1\[14\].modules.bubble VPWR VGND net328 sg13g2_dlygate4sd3_1
XFILLER_48_879 VPWR VGND sg13g2_decap_8
XFILLER_43_584 VPWR VGND sg13g2_fill_1
XFILLER_15_286 VPWR VGND sg13g2_fill_2
XFILLER_12_982 VPWR VGND sg13g2_decap_8
XFILLER_8_975 VPWR VGND sg13g2_decap_8
XFILLER_7_452 VPWR VGND sg13g2_decap_4
X_3420_ _1034_ _1033_ net1440 _1010_ net1445 VPWR VGND sg13g2_a22oi_1
XFILLER_3_691 VPWR VGND sg13g2_decap_8
X_6520__31 VPWR VGND net31 sg13g2_tiehi
X_6070_ _0628_ _0630_ _0631_ VPWR VGND sg13g2_nor2_1
XFILLER_38_312 VPWR VGND sg13g2_fill_1
X_5021_ _2472_ net1033 net494 VPWR VGND sg13g2_nand2_1
Xfanout1481 net1482 net1481 VPWR VGND sg13g2_buf_8
XFILLER_39_868 VPWR VGND sg13g2_fill_1
XFILLER_39_857 VPWR VGND sg13g2_fill_1
XFILLER_38_334 VPWR VGND sg13g2_fill_2
Xfanout1492 net1493 net1492 VPWR VGND sg13g2_buf_8
Xfanout1470 net1472 net1470 VPWR VGND sg13g2_buf_8
XFILLER_0_1013 VPWR VGND sg13g2_decap_8
X_5923_ _0494_ net1273 _0495_ _0496_ VPWR VGND sg13g2_a21o_1
X_5854_ VPWR _0033_ _0433_ VGND sg13g2_inv_1
XFILLER_34_573 VPWR VGND sg13g2_fill_2
XFILLER_34_595 VPWR VGND sg13g2_fill_1
X_4805_ VGND VPWR net1063 _2277_ _2280_ _2279_ sg13g2_a21oi_1
XFILLER_9_80 VPWR VGND sg13g2_decap_8
X_5785_ _0369_ VPWR _0370_ VGND _0357_ _0366_ sg13g2_o21ai_1
X_4736_ net995 _2872_ _2220_ VPWR VGND sg13g2_nor2_1
X_4667_ _2154_ _2153_ net1072 VPWR VGND sg13g2_nand2b_1
X_6406_ VGND VPWR net1240 _0928_ _0931_ _0930_ sg13g2_a21oi_1
X_3618_ net1381 _1160_ _1213_ VPWR VGND sg13g2_nor2_1
X_4598_ VGND VPWR _2097_ net1331 net339 sg13g2_or2_1
X_6337_ _0080_ _0868_ _0869_ _2805_ net1366 VPWR VGND sg13g2_a22oi_1
XFILLER_1_639 VPWR VGND sg13g2_decap_8
X_3549_ _1149_ net1206 _1150_ _1151_ VPWR VGND sg13g2_a21o_1
X_6268_ _0804_ VPWR _0805_ VGND net1246 _2805_ sg13g2_o21ai_1
X_6199_ net1252 s0.data_out\[17\]\[0\] _0747_ VPWR VGND sg13g2_and2_1
X_5219_ _2656_ VPWR _2657_ VGND net1465 net652 sg13g2_o21ai_1
XFILLER_29_301 VPWR VGND sg13g2_fill_1
XFILLER_29_345 VPWR VGND sg13g2_fill_2
XFILLER_38_890 VPWR VGND sg13g2_fill_2
XFILLER_12_212 VPWR VGND sg13g2_fill_1
XFILLER_40_532 VPWR VGND sg13g2_decap_8
XFILLER_8_238 VPWR VGND sg13g2_fill_1
XFILLER_5_934 VPWR VGND sg13g2_decap_8
XFILLER_4_433 VPWR VGND sg13g2_fill_2
XFILLER_4_466 VPWR VGND sg13g2_fill_2
XFILLER_4_488 VPWR VGND sg13g2_fill_2
XFILLER_48_676 VPWR VGND sg13g2_decap_8
XFILLER_29_890 VPWR VGND sg13g2_fill_1
X_5570_ net1416 _2973_ _2976_ VPWR VGND sg13g2_nor2_1
XFILLER_31_598 VPWR VGND sg13g2_decap_4
X_4521_ _2020_ net1080 net656 VPWR VGND sg13g2_nand2_1
X_4452_ _1963_ s0.data_out\[6\]\[5\] net1107 VPWR VGND sg13g2_nand2b_1
Xhold216 s0.data_out\[10\]\[7\] VPWR VGND net536 sg13g2_dlygate4sd3_1
Xhold205 s0.data_out\[16\]\[4\] VPWR VGND net525 sg13g2_dlygate4sd3_1
XFILLER_7_271 VPWR VGND sg13g2_fill_2
Xhold249 s0.data_out\[4\]\[4\] VPWR VGND net569 sg13g2_dlygate4sd3_1
X_3403_ VGND VPWR _0901_ _1016_ _1017_ net1225 sg13g2_a21oi_1
Xhold238 _0030_ VPWR VGND net558 sg13g2_dlygate4sd3_1
Xhold227 s0.data_out\[0\]\[0\] VPWR VGND net547 sg13g2_dlygate4sd3_1
X_4383_ net1103 net555 _1898_ VPWR VGND sg13g2_and2_1
X_6122_ net1478 net322 _0063_ VPWR VGND sg13g2_and2_1
X_6769__293 VPWR VGND net293 sg13g2_tiehi
X_6053_ s0.data_out\[19\]\[4\] s0.data_out\[18\]\[4\] net1270 _0614_ VPWR VGND sg13g2_mux2_1
X_5004_ VPWR _0258_ _2459_ VGND sg13g2_inv_1
X_5906_ net1276 net993 _0479_ VPWR VGND sg13g2_nor2_1
XFILLER_34_392 VPWR VGND sg13g2_fill_1
XFILLER_10_727 VPWR VGND sg13g2_fill_1
X_5837_ net1290 s0.data_out\[20\]\[1\] _0420_ VPWR VGND sg13g2_and2_1
XFILLER_10_738 VPWR VGND sg13g2_decap_4
X_5768_ VGND VPWR net1291 _0352_ _0353_ _0350_ sg13g2_a21oi_1
X_6592__249 VPWR VGND net249 sg13g2_tiehi
X_4719_ _2186_ _2203_ _2204_ _2205_ _2206_ VPWR VGND sg13g2_nor4_1
X_5699_ _3011_ VPWR _0296_ VGND _3066_ _3068_ sg13g2_o21ai_1
XFILLER_2_959 VPWR VGND sg13g2_decap_8
XFILLER_45_635 VPWR VGND sg13g2_fill_2
XFILLER_44_112 VPWR VGND sg13g2_decap_4
XFILLER_44_156 VPWR VGND sg13g2_decap_4
XFILLER_41_885 VPWR VGND sg13g2_fill_1
XFILLER_40_373 VPWR VGND sg13g2_fill_1
XFILLER_9_558 VPWR VGND sg13g2_fill_1
XFILLER_36_602 VPWR VGND sg13g2_fill_2
XFILLER_49_996 VPWR VGND sg13g2_decap_8
XFILLER_48_495 VPWR VGND sg13g2_fill_2
X_6740_ net89 VGND VPWR _0250_ s0.genblk1\[2\].modules.bubble clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_17_893 VPWR VGND sg13g2_fill_1
XFILLER_35_178 VPWR VGND sg13g2_decap_8
X_3952_ _1518_ net1432 _1516_ VPWR VGND sg13g2_nand2_1
X_6671_ net164 VGND VPWR net573 s0.data_out\[9\]\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3883_ _1451_ _1452_ _1453_ VPWR VGND sg13g2_nor2_1
X_5622_ net1462 net332 _0015_ VPWR VGND sg13g2_and2_1
X_5553_ _2958_ _2956_ _2959_ VPWR VGND _2957_ sg13g2_nand3b_1
X_4504_ _2007_ VPWR _2008_ VGND net1480 net627 sg13g2_o21ai_1
X_5484_ net1466 net333 _0000_ VPWR VGND sg13g2_and2_1
X_4435_ _1946_ net578 net1107 VPWR VGND sg13g2_nand2b_1
X_4366_ net1099 net632 _1885_ VPWR VGND sg13g2_and2_1
X_6105_ VPWR _0059_ net623 VGND sg13g2_inv_1
X_4297_ s0.data_out\[7\]\[0\] s0.data_out\[8\]\[0\] net1118 _1820_ VPWR VGND sg13g2_mux2_1
XFILLER_39_462 VPWR VGND sg13g2_fill_1
X_6036_ _0595_ net1261 _0596_ _0597_ VPWR VGND sg13g2_a21o_1
XFILLER_26_156 VPWR VGND sg13g2_fill_2
XFILLER_25_79 VPWR VGND sg13g2_fill_1
XFILLER_6_517 VPWR VGND sg13g2_decap_8
XFILLER_2_756 VPWR VGND sg13g2_decap_8
XFILLER_49_204 VPWR VGND sg13g2_fill_1
XFILLER_46_911 VPWR VGND sg13g2_decap_8
XFILLER_18_635 VPWR VGND sg13g2_fill_1
XFILLER_17_123 VPWR VGND sg13g2_fill_1
XFILLER_46_988 VPWR VGND sg13g2_decap_8
XFILLER_45_476 VPWR VGND sg13g2_fill_2
XFILLER_26_690 VPWR VGND sg13g2_fill_2
XFILLER_9_366 VPWR VGND sg13g2_decap_4
XFILLER_12_1024 VPWR VGND sg13g2_decap_4
X_4220_ _1744_ VPWR _1755_ VGND net1442 _1716_ sg13g2_o21ai_1
X_4151_ net1482 net324 _0178_ VPWR VGND sg13g2_and2_1
X_4082_ _1629_ net1013 _1628_ VPWR VGND sg13g2_nand2_1
XFILLER_49_793 VPWR VGND sg13g2_decap_8
XFILLER_37_966 VPWR VGND sg13g2_decap_8
XFILLER_36_432 VPWR VGND sg13g2_fill_1
X_4984_ net1036 s0.data_out\[2\]\[2\] _2444_ VPWR VGND sg13g2_and2_1
X_6723_ net108 VGND VPWR _0233_ s0.data_out\[5\]\[5\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_3935_ net1414 _1499_ _1501_ VPWR VGND sg13g2_nor2_1
XFILLER_20_822 VPWR VGND sg13g2_fill_1
X_6654_ net182 VGND VPWR _0164_ s0.data_new_delayed\[5\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_5605_ net1324 VPWR _3004_ VGND _2953_ _3003_ sg13g2_o21ai_1
X_3866_ VPWR _0141_ net617 VGND sg13g2_inv_1
X_6585_ net257 VGND VPWR _0095_ s0.data_out\[16\]\[6\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3797_ net1182 net1144 _1376_ VPWR VGND sg13g2_nor2b_1
X_5536_ net1323 _2940_ _2941_ _2942_ VPWR VGND sg13g2_nor3_1
X_5467_ s0.was_valid_out\[23\][0] net1326 _2885_ VPWR VGND sg13g2_nor2_1
X_4418_ _1815_ VPWR _1929_ VGND net1105 _2864_ sg13g2_o21ai_1
X_5398_ VPWR _2816_ net553 VGND sg13g2_inv_1
X_4349_ _1860_ VPWR _1872_ VGND _1867_ _1868_ sg13g2_o21ai_1
X_6019_ _0580_ net1278 _0579_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_955 VPWR VGND sg13g2_decap_8
XFILLER_43_914 VPWR VGND sg13g2_decap_8
XFILLER_15_627 VPWR VGND sg13g2_fill_2
XFILLER_14_126 VPWR VGND sg13g2_fill_1
X_6778__156 VPWR VGND net156 sg13g2_tiehi
XFILLER_27_498 VPWR VGND sg13g2_fill_2
XFILLER_35_1002 VPWR VGND sg13g2_decap_8
XFILLER_11_833 VPWR VGND sg13g2_decap_4
XFILLER_23_671 VPWR VGND sg13g2_decap_8
XFILLER_10_321 VPWR VGND sg13g2_decap_8
XFILLER_6_303 VPWR VGND sg13g2_fill_1
XFILLER_6_369 VPWR VGND sg13g2_fill_2
XFILLER_42_1006 VPWR VGND sg13g2_decap_8
XFILLER_19_911 VPWR VGND sg13g2_decap_8
XFILLER_46_785 VPWR VGND sg13g2_decap_8
XFILLER_18_487 VPWR VGND sg13g2_decap_8
XFILLER_33_435 VPWR VGND sg13g2_decap_4
X_3720_ net1378 _1239_ _1308_ VPWR VGND sg13g2_nor2_1
XFILLER_20_107 VPWR VGND sg13g2_fill_2
X_3651_ s0.data_out\[13\]\[0\] s0.data_out\[12\]\[0\] net1197 _1241_ VPWR VGND sg13g2_mux2_1
XFILLER_9_196 VPWR VGND sg13g2_fill_2
X_6370_ net1225 net1164 _0895_ VPWR VGND sg13g2_nor2b_1
X_3582_ _1184_ _2768_ _1182_ VPWR VGND sg13g2_xnor2_1
X_5321_ VPWR _2739_ net392 VGND sg13g2_inv_1
X_5252_ _2682_ VPWR _2683_ VGND net1006 _2681_ sg13g2_o21ai_1
X_5183_ net1031 _2618_ _2622_ VPWR VGND sg13g2_nor2_1
X_4203_ s0.data_out\[9\]\[5\] s0.data_out\[8\]\[5\] net1121 _1738_ VPWR VGND sg13g2_mux2_1
X_4134_ _0174_ _1672_ _1673_ _2842_ net1386 VPWR VGND sg13g2_a22oi_1
XFILLER_49_590 VPWR VGND sg13g2_decap_8
X_4065_ _1612_ net1132 net509 VPWR VGND sg13g2_nand2_1
XFILLER_37_774 VPWR VGND sg13g2_fill_2
XFILLER_24_402 VPWR VGND sg13g2_fill_1
XFILLER_25_914 VPWR VGND sg13g2_fill_1
XFILLER_24_468 VPWR VGND sg13g2_fill_1
XFILLER_40_939 VPWR VGND sg13g2_decap_8
X_4967_ _2429_ VPWR _2430_ VGND net1428 _2427_ sg13g2_o21ai_1
X_4898_ VGND VPWR _2359_ _2362_ _0248_ _2363_ sg13g2_a21oi_1
Xclkbuf_leaf_31_clk clknet_3_5__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
XFILLER_20_652 VPWR VGND sg13g2_decap_8
X_6706_ net126 VGND VPWR _0216_ s0.data_out\[6\]\[0\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3918_ _1484_ _1483_ net1441 _1460_ net1445 VPWR VGND sg13g2_a22oi_1
X_6637_ net200 VGND VPWR _0147_ s0.genblk1\[10\].modules.bubble clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_3849_ VGND VPWR net1016 _1356_ _1425_ net1385 sg13g2_a21oi_1
X_6568_ net275 VGND VPWR _0078_ s0.data_out\[17\]\[1\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_5519_ net1315 net1170 _2925_ VPWR VGND sg13g2_nor2b_1
X_6499_ net54 VGND VPWR net417 s0.data_out\[23\]\[4\] clknet_leaf_0_clk sg13g2_dfrbpq_1
Xfanout1107 net1109 net1107 VPWR VGND sg13g2_buf_8
Xfanout1129 net1130 net1129 VPWR VGND sg13g2_buf_1
Xfanout1118 net1119 net1118 VPWR VGND sg13g2_buf_8
XFILLER_47_11 VPWR VGND sg13g2_decap_8
XFILLER_43_711 VPWR VGND sg13g2_fill_2
XFILLER_27_295 VPWR VGND sg13g2_decap_4
XFILLER_24_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_22_clk clknet_3_7__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_3_873 VPWR VGND sg13g2_decap_8
XFILLER_38_538 VPWR VGND sg13g2_decap_8
XFILLER_38_549 VPWR VGND sg13g2_fill_2
X_5870_ _0446_ _0445_ _0444_ VPWR VGND sg13g2_nand2b_1
X_4821_ VGND VPWR net1064 _2293_ _2296_ _2295_ sg13g2_a21oi_1
XFILLER_34_799 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_13_clk clknet_3_3__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_4752_ _2201_ _2232_ net1475 _2233_ VPWR VGND sg13g2_nand3_1
X_4683_ s0.data_out\[5\]\[6\] s0.data_out\[4\]\[6\] net1070 _2170_ VPWR VGND sg13g2_mux2_1
X_3703_ VGND VPWR _1279_ _1281_ _1293_ net1423 sg13g2_a21oi_1
XFILLER_30_961 VPWR VGND sg13g2_decap_8
X_6422_ net1223 net1158 _0947_ VPWR VGND sg13g2_nor2b_1
X_3634_ VGND VPWR _1222_ _1225_ _0121_ _1226_ sg13g2_a21oi_1
X_6353_ net1250 VPWR _0882_ VGND _0815_ _0881_ sg13g2_o21ai_1
X_3565_ s0.data_out\[14\]\[5\] s0.data_out\[13\]\[5\] net1211 _1167_ VPWR VGND sg13g2_mux2_1
X_3496_ VPWR _0107_ net694 VGND sg13g2_inv_1
X_6284_ s0.data_out\[17\]\[6\] s0.data_out\[16\]\[6\] net1245 _0821_ VPWR VGND sg13g2_mux2_1
X_5304_ VGND VPWR net1465 _2705_ _0292_ _2725_ sg13g2_a21oi_1
XFILLER_25_1001 VPWR VGND sg13g2_decap_8
X_5235_ VGND VPWR net1021 net385 _2669_ _2634_ sg13g2_a21oi_1
X_5166_ s0.data_out\[1\]\[3\] s0.data_out\[0\]\[3\] net1024 _2605_ VPWR VGND sg13g2_mux2_1
X_5097_ VGND VPWR net1009 _2479_ _2547_ net1348 sg13g2_a21oi_1
X_4117_ net1127 s0.data_out\[9\]\[3\] _1660_ VPWR VGND sg13g2_and2_1
X_4048_ _1593_ net1130 _1594_ _1595_ VPWR VGND sg13g2_a21o_1
XFILLER_13_917 VPWR VGND sg13g2_decap_4
X_5999_ net1470 _0556_ _0050_ VPWR VGND sg13g2_and2_1
XFILLER_32_1027 VPWR VGND sg13g2_fill_2
XFILLER_4_626 VPWR VGND sg13g2_decap_8
XFILLER_0_810 VPWR VGND sg13g2_decap_8
Xhold9 s0.genblk1\[10\].modules.bubble VPWR VGND net329 sg13g2_dlygate4sd3_1
XFILLER_0_887 VPWR VGND sg13g2_decap_8
XFILLER_48_858 VPWR VGND sg13g2_decap_8
XFILLER_28_571 VPWR VGND sg13g2_fill_2
XFILLER_43_552 VPWR VGND sg13g2_fill_2
XFILLER_43_541 VPWR VGND sg13g2_fill_2
XFILLER_31_725 VPWR VGND sg13g2_fill_1
XFILLER_31_758 VPWR VGND sg13g2_decap_4
X_6738__92 VPWR VGND net92 sg13g2_tiehi
XFILLER_12_961 VPWR VGND sg13g2_decap_8
XFILLER_8_954 VPWR VGND sg13g2_decap_8
XFILLER_7_431 VPWR VGND sg13g2_fill_1
XFILLER_11_471 VPWR VGND sg13g2_fill_1
XFILLER_48_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_670 VPWR VGND sg13g2_decap_8
X_5020_ net1463 net335 _0262_ VPWR VGND sg13g2_and2_1
XFILLER_39_836 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_2_clk clknet_3_0__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
Xfanout1471 net1472 net1471 VPWR VGND sg13g2_buf_1
Xfanout1460 net1461 net1460 VPWR VGND sg13g2_buf_8
Xfanout1482 net1483 net1482 VPWR VGND sg13g2_buf_8
Xfanout1493 rst_n net1493 VPWR VGND sg13g2_buf_8
XFILLER_38_379 VPWR VGND sg13g2_fill_2
X_5922_ net1273 net1148 _0495_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_72 VPWR VGND sg13g2_decap_8
XFILLER_34_530 VPWR VGND sg13g2_fill_2
X_5853_ _0432_ VPWR _0433_ VGND net1462 net609 sg13g2_o21ai_1
XFILLER_22_736 VPWR VGND sg13g2_fill_2
X_5784_ _0369_ net1437 _0365_ VPWR VGND sg13g2_nand2_1
X_4804_ VGND VPWR _2156_ _2278_ _2279_ net1060 sg13g2_a21oi_1
X_4735_ _0229_ _2218_ _2219_ _2865_ net1363 VPWR VGND sg13g2_a22oi_1
X_4666_ _2043_ VPWR _2153_ VGND net1080 _2872_ sg13g2_o21ai_1
X_4597_ _2095_ _2094_ _2096_ VPWR VGND sg13g2_nor2b_1
X_6405_ VGND VPWR _0820_ _0929_ _0930_ net1240 sg13g2_a21oi_1
X_3617_ net1218 VPWR _1212_ VGND _1157_ _1211_ sg13g2_o21ai_1
X_3548_ net1206 net1145 _1150_ VPWR VGND sg13g2_nor2b_1
X_6336_ net1365 _0809_ _0869_ VPWR VGND sg13g2_nor2_1
XFILLER_1_618 VPWR VGND sg13g2_decap_8
X_6267_ _0804_ net1246 net482 VPWR VGND sg13g2_nand2_1
X_3479_ net1018 _2822_ _1089_ VPWR VGND sg13g2_nor2_1
X_6198_ VGND VPWR _0742_ _0745_ _0064_ _0746_ sg13g2_a21oi_1
X_5218_ _2655_ VPWR _2656_ VGND net1004 _2654_ sg13g2_o21ai_1
XFILLER_28_46 VPWR VGND sg13g2_fill_2
X_5149_ VGND VPWR net1004 _2583_ _2588_ _2587_ sg13g2_a21oi_1
XFILLER_44_338 VPWR VGND sg13g2_fill_2
XFILLER_37_390 VPWR VGND sg13g2_fill_2
XFILLER_13_769 VPWR VGND sg13g2_fill_1
X_6735__95 VPWR VGND net95 sg13g2_tiehi
XFILLER_5_913 VPWR VGND sg13g2_decap_8
XFILLER_48_611 VPWR VGND sg13g2_decap_8
XFILLER_0_684 VPWR VGND sg13g2_decap_8
XFILLER_48_655 VPWR VGND sg13g2_decap_8
XFILLER_35_338 VPWR VGND sg13g2_decap_4
XFILLER_43_382 VPWR VGND sg13g2_fill_1
X_6578__264 VPWR VGND net264 sg13g2_tiehi
X_4520_ net1474 net331 _0214_ VPWR VGND sg13g2_and2_1
XFILLER_11_290 VPWR VGND sg13g2_fill_2
X_4451_ _1960_ net1090 _1961_ _1962_ VPWR VGND sg13g2_a21o_1
Xhold206 _0093_ VPWR VGND net526 sg13g2_dlygate4sd3_1
Xhold217 s0.data_out\[8\]\[0\] VPWR VGND net537 sg13g2_dlygate4sd3_1
Xhold239 s0.was_valid_out\[23\][0] VPWR VGND net559 sg13g2_dlygate4sd3_1
Xhold228 s0.data_out\[14\]\[2\] VPWR VGND net548 sg13g2_dlygate4sd3_1
X_3402_ _1016_ s0.data_out\[14\]\[1\] net1235 VPWR VGND sg13g2_nand2b_1
X_4382_ VPWR _0198_ net655 VGND sg13g2_inv_1
X_6121_ net1356 _0665_ _0062_ VPWR VGND sg13g2_nor2_1
X_6052_ _0613_ net1271 net440 VPWR VGND sg13g2_nand2_1
X_5003_ _2458_ VPWR _2459_ VGND net1475 net678 sg13g2_o21ai_1
X_6585__257 VPWR VGND net257 sg13g2_tiehi
XFILLER_22_1015 VPWR VGND sg13g2_decap_8
Xfanout1290 net1292 net1290 VPWR VGND sg13g2_buf_2
XFILLER_26_338 VPWR VGND sg13g2_fill_2
X_6702__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_35_850 VPWR VGND sg13g2_fill_2
XFILLER_35_872 VPWR VGND sg13g2_fill_2
X_5905_ _0477_ VPWR _0478_ VGND net1283 _2788_ sg13g2_o21ai_1
XFILLER_34_360 VPWR VGND sg13g2_fill_1
X_5836_ VPWR _0029_ _0419_ VGND sg13g2_inv_1
X_5767_ s0.data_out\[21\]\[2\] s0.data_out\[20\]\[2\] net1297 _0352_ VPWR VGND sg13g2_mux2_1
X_4718_ VGND VPWR _2199_ _2201_ _2205_ net1418 sg13g2_a21oi_1
X_5698_ _3092_ _3091_ _3069_ VPWR VGND sg13g2_nand2b_1
X_4649_ net1061 net1167 _2136_ VPWR VGND sg13g2_nor2b_1
X_6732__98 VPWR VGND net98 sg13g2_tiehi
XFILLER_30_58 VPWR VGND sg13g2_fill_1
XFILLER_2_938 VPWR VGND sg13g2_decap_8
X_6319_ VPWR VGND _0831_ _0855_ _0854_ _0812_ _0856_ _0853_ sg13g2_a221oi_1
XFILLER_7_1009 VPWR VGND sg13g2_decap_8
XFILLER_29_110 VPWR VGND sg13g2_fill_1
XFILLER_29_165 VPWR VGND sg13g2_decap_8
XFILLER_44_124 VPWR VGND sg13g2_fill_1
XFILLER_40_385 VPWR VGND sg13g2_decap_8
XFILLER_5_721 VPWR VGND sg13g2_fill_2
XFILLER_45_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_91 VPWR VGND sg13g2_fill_1
XFILLER_0_481 VPWR VGND sg13g2_decap_8
XFILLER_1_982 VPWR VGND sg13g2_decap_8
XFILLER_49_975 VPWR VGND sg13g2_decap_8
XFILLER_35_113 VPWR VGND sg13g2_fill_1
XFILLER_24_809 VPWR VGND sg13g2_decap_8
XFILLER_17_861 VPWR VGND sg13g2_fill_1
X_3951_ net1432 _1516_ _1517_ VPWR VGND sg13g2_nor2_1
XFILLER_44_680 VPWR VGND sg13g2_fill_1
X_6670_ net165 VGND VPWR _0180_ s0.data_out\[9\]\[0\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3882_ VGND VPWR _2733_ _2745_ _1452_ net1185 sg13g2_a21oi_1
X_5621_ net1463 _3011_ _0014_ VPWR VGND sg13g2_and2_1
X_5552_ VGND VPWR _2958_ _2955_ net1407 sg13g2_or2_1
X_4503_ _2006_ net1480 _2007_ VPWR VGND _1947_ sg13g2_nand3b_1
X_6591__250 VPWR VGND net250 sg13g2_tiehi
X_5483_ _2893_ VPWR net9 VGND _2764_ net991 sg13g2_o21ai_1
X_4434_ _1943_ net1089 _1944_ _1945_ VPWR VGND sg13g2_a21o_1
X_4365_ _0194_ _1883_ _1884_ _2852_ net1374 VPWR VGND sg13g2_a22oi_1
X_6104_ _0657_ VPWR _0658_ VGND net1470 net622 sg13g2_o21ai_1
X_6035_ net1261 net1143 _0596_ VPWR VGND sg13g2_nor2b_1
X_4296_ _1819_ net1110 _1818_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_496 VPWR VGND sg13g2_decap_4
XFILLER_26_135 VPWR VGND sg13g2_decap_8
XFILLER_26_146 VPWR VGND sg13g2_fill_2
XFILLER_42_617 VPWR VGND sg13g2_decap_4
XFILLER_26_168 VPWR VGND sg13g2_decap_4
XFILLER_41_138 VPWR VGND sg13g2_decap_8
X_5819_ _0404_ net1008 _0403_ VPWR VGND sg13g2_nand2_1
XFILLER_10_525 VPWR VGND sg13g2_fill_2
XFILLER_22_363 VPWR VGND sg13g2_decap_8
XFILLER_23_897 VPWR VGND sg13g2_fill_1
XFILLER_2_735 VPWR VGND sg13g2_decap_8
XFILLER_46_967 VPWR VGND sg13g2_decap_8
XFILLER_14_831 VPWR VGND sg13g2_fill_2
XFILLER_33_639 VPWR VGND sg13g2_decap_4
XFILLER_13_352 VPWR VGND sg13g2_fill_1
XFILLER_14_875 VPWR VGND sg13g2_decap_4
XFILLER_9_323 VPWR VGND sg13g2_fill_1
XFILLER_9_334 VPWR VGND sg13g2_decap_8
XFILLER_12_1003 VPWR VGND sg13g2_decap_8
XFILLER_31_90 VPWR VGND sg13g2_fill_1
X_4150_ net1384 _1680_ _0177_ VPWR VGND sg13g2_nor2_1
X_4081_ s0.data_out\[9\]\[4\] s0.data_out\[10\]\[4\] net1175 _1628_ VPWR VGND sg13g2_mux2_1
XFILLER_49_772 VPWR VGND sg13g2_decap_8
XFILLER_37_934 VPWR VGND sg13g2_fill_2
XFILLER_37_945 VPWR VGND sg13g2_decap_8
XFILLER_23_116 VPWR VGND sg13g2_decap_4
X_4983_ _0253_ _2442_ _2443_ _2879_ net1358 VPWR VGND sg13g2_a22oi_1
X_3934_ _1500_ _1499_ net1414 _1492_ net1405 VPWR VGND sg13g2_a22oi_1
X_6722_ net109 VGND VPWR _0232_ s0.data_out\[5\]\[4\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_6653_ net183 VGND VPWR _0163_ s0.data_new_delayed\[4\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3865_ _1437_ VPWR _1438_ VGND net1490 net616 sg13g2_o21ai_1
X_5604_ net1012 _2765_ _3003_ VPWR VGND sg13g2_nor2_1
X_6584_ net258 VGND VPWR net476 s0.data_out\[16\]\[5\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_3796_ s0.data_out\[12\]\[7\] s0.data_out\[11\]\[7\] net1188 _1375_ VPWR VGND sg13g2_mux2_1
X_5535_ net1327 net377 _2941_ VPWR VGND sg13g2_nor2_1
X_5466_ VPWR _2884_ net494 VGND sg13g2_inv_1
X_4417_ _1928_ net1096 _1927_ VPWR VGND sg13g2_nand2b_1
X_5397_ VPWR _2815_ net430 VGND sg13g2_inv_1
X_4348_ _1852_ _1868_ _1869_ _1870_ _1871_ VPWR VGND sg13g2_nor4_1
X_4279_ net1098 net1164 _1802_ VPWR VGND sg13g2_nor2b_1
X_6018_ VGND VPWR net1265 _0577_ _0579_ _0578_ sg13g2_a21oi_1
XFILLER_36_35 VPWR VGND sg13g2_fill_1
XFILLER_15_606 VPWR VGND sg13g2_decap_8
XFILLER_10_377 VPWR VGND sg13g2_fill_1
XFILLER_10_366 VPWR VGND sg13g2_decap_8
XFILLER_46_764 VPWR VGND sg13g2_decap_8
XFILLER_42_992 VPWR VGND sg13g2_decap_8
X_3650_ VGND VPWR net1202 _1237_ _1240_ _1239_ sg13g2_a21oi_1
X_3581_ VGND VPWR _1183_ _1182_ _2768_ sg13g2_or2_1
X_5320_ VPWR _2738_ net366 VGND sg13g2_inv_1
X_5251_ VGND VPWR _2754_ _2612_ _2682_ net1347 sg13g2_a21oi_1
XFILLER_6_893 VPWR VGND sg13g2_decap_8
X_4202_ _1737_ net1120 net687 VPWR VGND sg13g2_nand2_1
X_5182_ VGND VPWR net1022 _2619_ _2621_ _2620_ sg13g2_a21oi_1
X_4133_ net1386 _1617_ _1673_ VPWR VGND sg13g2_nor2_1
X_4064_ VGND VPWR net1139 _1608_ _1611_ _1610_ sg13g2_a21oi_1
XFILLER_37_731 VPWR VGND sg13g2_fill_2
XFILLER_25_959 VPWR VGND sg13g2_decap_8
XFILLER_12_609 VPWR VGND sg13g2_decap_8
X_6705_ net127 VGND VPWR _0215_ s0.shift_out\[6\][0] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_4966_ _2421_ _2428_ _2429_ VPWR VGND sg13g2_nor2b_1
X_4897_ net1473 VPWR _2363_ VGND net524 _2357_ sg13g2_o21ai_1
X_3917_ VGND VPWR net1181 _1480_ _1483_ _1482_ sg13g2_a21oi_1
X_3848_ VGND VPWR net1180 net422 _1424_ _1354_ sg13g2_a21oi_1
X_6636_ net201 VGND VPWR _0146_ s0.genblk1\[11\].modules.bubble clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
XFILLER_20_686 VPWR VGND sg13g2_fill_1
X_6567_ net276 VGND VPWR _0077_ s0.data_out\[17\]\[0\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3779_ _1357_ VPWR _1358_ VGND net1016 _1355_ sg13g2_o21ai_1
X_5518_ _2923_ VPWR _2924_ VGND net1320 _2778_ sg13g2_o21ai_1
X_6498_ net55 VGND VPWR _0008_ s0.data_out\[23\]\[3\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5449_ VPWR _2867_ net488 VGND sg13g2_inv_1
Xfanout1119 s0.valid_out\[8\][0] net1119 VPWR VGND sg13g2_buf_8
Xfanout1108 net1109 net1108 VPWR VGND sg13g2_buf_2
XFILLER_47_34 VPWR VGND sg13g2_fill_1
XFILLER_47_67 VPWR VGND sg13g2_fill_2
XFILLER_28_731 VPWR VGND sg13g2_fill_2
XFILLER_28_775 VPWR VGND sg13g2_fill_2
XFILLER_16_959 VPWR VGND sg13g2_decap_8
XFILLER_42_233 VPWR VGND sg13g2_decap_8
XFILLER_42_288 VPWR VGND sg13g2_fill_1
XFILLER_24_970 VPWR VGND sg13g2_decap_8
XFILLER_31_929 VPWR VGND sg13g2_fill_1
XFILLER_6_101 VPWR VGND sg13g2_fill_2
XFILLER_3_852 VPWR VGND sg13g2_decap_8
XFILLER_19_753 VPWR VGND sg13g2_fill_1
XFILLER_18_274 VPWR VGND sg13g2_fill_1
X_4820_ VGND VPWR _2169_ _2294_ _2295_ net1064 sg13g2_a21oi_1
XFILLER_22_929 VPWR VGND sg13g2_fill_2
X_4751_ net1077 VPWR _2232_ VGND _2197_ _2231_ sg13g2_o21ai_1
XFILLER_15_992 VPWR VGND sg13g2_decap_8
XFILLER_30_940 VPWR VGND sg13g2_decap_8
X_4682_ _2169_ net1069 net507 VPWR VGND sg13g2_nand2_1
X_3702_ net1440 _1255_ _1292_ VPWR VGND sg13g2_nor2_1
X_6421_ _0945_ VPWR _0946_ VGND net1233 _2810_ sg13g2_o21ai_1
X_3633_ net1486 VPWR _1226_ VGND net566 _1220_ sg13g2_o21ai_1
XFILLER_6_690 VPWR VGND sg13g2_fill_1
X_6352_ net1236 net503 _0881_ VPWR VGND sg13g2_and2_1
X_3564_ _1166_ _1162_ _1164_ _1165_ VPWR VGND sg13g2_and3_1
X_3495_ _1101_ VPWR _1102_ VGND net1485 net693 sg13g2_o21ai_1
X_6283_ _0820_ net1247 net599 VPWR VGND sg13g2_nand2_1
X_5303_ net1464 net385 _2725_ VPWR VGND sg13g2_nor2_1
X_5234_ VPWR _0279_ net542 VGND sg13g2_inv_1
X_5165_ s0.data_out\[0\]\[3\] s0.data_out\[1\]\[3\] net1033 _2604_ VPWR VGND sg13g2_mux2_1
X_4116_ VPWR _0170_ _1659_ VGND sg13g2_inv_1
X_5096_ VGND VPWR net1027 net652 _2546_ _2481_ sg13g2_a21oi_1
XFILLER_17_26 VPWR VGND sg13g2_fill_1
X_4047_ net1130 s0.data_new_delayed\[3\] _1594_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_211 VPWR VGND sg13g2_decap_8
XFILLER_24_244 VPWR VGND sg13g2_fill_1
XFILLER_25_745 VPWR VGND sg13g2_decap_8
X_5998_ VGND VPWR _2738_ _0556_ _0049_ _0561_ sg13g2_a21oi_1
XFILLER_40_748 VPWR VGND sg13g2_fill_2
X_4949_ _2411_ _2409_ _2412_ VPWR VGND _2410_ sg13g2_nand3b_1
X_6636__201 VPWR VGND net201 sg13g2_tiehi
X_6747__82 VPWR VGND net82 sg13g2_tiehi
XFILLER_32_1006 VPWR VGND sg13g2_decap_8
X_6619_ net220 VGND VPWR _0129_ s0.data_out\[13\]\[4\] clknet_leaf_28_clk sg13g2_dfrbpq_2
XFILLER_0_866 VPWR VGND sg13g2_decap_8
XFILLER_48_837 VPWR VGND sg13g2_decap_8
XFILLER_16_712 VPWR VGND sg13g2_fill_2
XFILLER_15_255 VPWR VGND sg13g2_decap_4
XFILLER_15_288 VPWR VGND sg13g2_fill_1
XFILLER_30_269 VPWR VGND sg13g2_fill_1
XFILLER_8_933 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_decap_8
Xfanout1450 net1451 net1450 VPWR VGND sg13g2_buf_1
Xfanout1472 net1476 net1472 VPWR VGND sg13g2_buf_8
Xfanout1461 ui_in[0] net1461 VPWR VGND sg13g2_buf_8
Xfanout1483 net1493 net1483 VPWR VGND sg13g2_buf_8
XFILLER_47_892 VPWR VGND sg13g2_decap_8
X_5921_ s0.data_out\[20\]\[6\] s0.data_out\[19\]\[6\] net1281 _0494_ VPWR VGND sg13g2_mux2_1
XFILLER_0_51 VPWR VGND sg13g2_decap_4
X_5852_ _0431_ VPWR _0432_ VGND _2752_ _0430_ sg13g2_o21ai_1
XFILLER_34_575 VPWR VGND sg13g2_fill_1
X_5783_ _0349_ _0358_ _0366_ _0367_ _0368_ VPWR VGND sg13g2_nor4_1
X_4803_ _2278_ s0.data_out\[3\]\[3\] net1067 VPWR VGND sg13g2_nand2b_1
XFILLER_21_269 VPWR VGND sg13g2_fill_1
X_4734_ net1363 _2139_ _2219_ VPWR VGND sg13g2_nor2_1
X_6744__85 VPWR VGND net85 sg13g2_tiehi
X_4665_ _2152_ net1072 _2151_ VPWR VGND sg13g2_nand2b_1
X_4596_ _2014_ VPWR _2095_ VGND _2070_ _2072_ sg13g2_o21ai_1
X_6404_ _0929_ s0.data_out\[15\]\[6\] net1247 VPWR VGND sg13g2_nand2b_1
X_3616_ net1206 s0.data_out\[13\]\[6\] _1211_ VPWR VGND sg13g2_and2_1
X_3547_ _1148_ VPWR _1149_ VGND net1211 _2819_ sg13g2_o21ai_1
X_6335_ net1254 VPWR _0868_ VGND _0806_ _0867_ sg13g2_o21ai_1
X_3478_ _0103_ _1087_ _1088_ _2817_ net1368 VPWR VGND sg13g2_a22oi_1
X_6266_ VPWR VGND _0801_ net1460 _0799_ net1453 _0803_ _0795_ sg13g2_a221oi_1
X_6197_ VGND VPWR _0746_ net1330 net337 sg13g2_or2_1
X_5217_ VGND VPWR net1004 _2595_ _2655_ net1346 sg13g2_a21oi_1
X_5148_ net1004 _2586_ _2587_ VPWR VGND sg13g2_nor2_1
XFILLER_45_807 VPWR VGND sg13g2_decap_4
X_5079_ net1030 net1151 _2530_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_347 VPWR VGND sg13g2_fill_1
XFILLER_44_328 VPWR VGND sg13g2_fill_1
XFILLER_44_46 VPWR VGND sg13g2_fill_2
XFILLER_13_704 VPWR VGND sg13g2_decap_4
XFILLER_8_229 VPWR VGND sg13g2_decap_8
XFILLER_20_280 VPWR VGND sg13g2_fill_1
XFILLER_5_969 VPWR VGND sg13g2_decap_8
XFILLER_0_663 VPWR VGND sg13g2_decap_8
XFILLER_48_634 VPWR VGND sg13g2_decap_8
XFILLER_16_564 VPWR VGND sg13g2_decap_4
XFILLER_8_752 VPWR VGND sg13g2_fill_1
X_4450_ net1090 net1153 _1961_ VPWR VGND sg13g2_nor2b_1
XFILLER_7_262 VPWR VGND sg13g2_decap_4
Xhold207 s0.data_out\[21\]\[7\] VPWR VGND net527 sg13g2_dlygate4sd3_1
X_4381_ _1896_ VPWR _1897_ VGND net1481 net654 sg13g2_o21ai_1
X_6741__88 VPWR VGND net88 sg13g2_tiehi
X_3401_ _1014_ net1213 _1012_ _1015_ VPWR VGND sg13g2_a21o_1
Xhold218 _1878_ VPWR VGND net538 sg13g2_dlygate4sd3_1
Xhold229 s0.data_out\[5\]\[3\] VPWR VGND net549 sg13g2_dlygate4sd3_1
X_6120_ VGND VPWR _0667_ _0670_ _0061_ _0671_ sg13g2_a21oi_1
X_6051_ _0612_ _0608_ _0609_ _0610_ VPWR VGND sg13g2_and3_1
X_5002_ _2457_ net1475 _2458_ VPWR VGND _2407_ sg13g2_nand3b_1
XFILLER_39_634 VPWR VGND sg13g2_fill_2
XFILLER_15_0 VPWR VGND sg13g2_fill_1
Xfanout1291 net1292 net1291 VPWR VGND sg13g2_buf_1
Xfanout1280 s0.shift_out\[19\][0] net1280 VPWR VGND sg13g2_buf_2
XFILLER_27_807 VPWR VGND sg13g2_fill_2
XFILLER_38_166 VPWR VGND sg13g2_fill_2
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
X_5904_ _0477_ net1284 net690 VPWR VGND sg13g2_nand2_1
X_5835_ _0418_ VPWR _0419_ VGND net1463 net648 sg13g2_o21ai_1
XFILLER_34_383 VPWR VGND sg13g2_decap_8
XFILLER_22_545 VPWR VGND sg13g2_fill_1
X_5766_ _0351_ net1298 net424 VPWR VGND sg13g2_nand2_1
X_4717_ VGND VPWR _2191_ _2193_ _2204_ net1427 sg13g2_a21oi_1
X_5697_ _3085_ VPWR _3091_ VGND _3077_ _3088_ sg13g2_o21ai_1
X_4648_ _2134_ VPWR _2135_ VGND net1068 _2865_ sg13g2_o21ai_1
XFILLER_2_917 VPWR VGND sg13g2_decap_8
X_4579_ s0.data_out\[5\]\[4\] s0.data_out\[6\]\[4\] net1093 _2078_ VPWR VGND sg13g2_mux2_1
X_6318_ _0775_ VPWR _0855_ VGND _0827_ _0830_ sg13g2_o21ai_1
X_6249_ VGND VPWR _0672_ _0785_ _0786_ net1254 sg13g2_a21oi_1
XFILLER_29_122 VPWR VGND sg13g2_fill_1
XFILLER_45_615 VPWR VGND sg13g2_decap_4
XFILLER_17_317 VPWR VGND sg13g2_fill_2
XFILLER_38_1012 VPWR VGND sg13g2_decap_8
XFILLER_13_501 VPWR VGND sg13g2_decap_4
XFILLER_41_854 VPWR VGND sg13g2_fill_2
XFILLER_45_1005 VPWR VGND sg13g2_decap_8
XFILLER_1_961 VPWR VGND sg13g2_decap_8
XFILLER_49_954 VPWR VGND sg13g2_decap_8
XFILLER_36_615 VPWR VGND sg13g2_decap_4
Xhold90 s0.data_out\[18\]\[3\] VPWR VGND net410 sg13g2_dlygate4sd3_1
XFILLER_23_309 VPWR VGND sg13g2_fill_2
X_3950_ VGND VPWR net1185 _1513_ _1516_ _1515_ sg13g2_a21oi_1
XFILLER_16_372 VPWR VGND sg13g2_fill_1
XFILLER_32_876 VPWR VGND sg13g2_decap_8
X_3881_ net1140 _1445_ _1451_ VPWR VGND sg13g2_nor2_1
X_5620_ VGND VPWR _2739_ _3011_ _0013_ _3016_ sg13g2_a21oi_1
XFILLER_31_375 VPWR VGND sg13g2_decap_4
X_5551_ net1398 _2947_ _2957_ VPWR VGND sg13g2_nor2_1
X_4502_ net1100 VPWR _2006_ VGND _1944_ _2005_ sg13g2_o21ai_1
XFILLER_6_50 VPWR VGND sg13g2_fill_1
X_5482_ _2893_ net1398 net992 VPWR VGND sg13g2_nand2_1
X_4433_ net1089 net1149 _1944_ VPWR VGND sg13g2_nor2b_1
X_4364_ net1374 _1805_ _1884_ VPWR VGND sg13g2_nor2_1
X_6103_ _0656_ net1470 _0657_ VPWR VGND _0606_ sg13g2_nand3b_1
X_4295_ VGND VPWR net1098 _1816_ _1818_ _1817_ sg13g2_a21oi_1
X_6034_ s0.data_out\[19\]\[7\] s0.data_out\[18\]\[7\] net1269 _0595_ VPWR VGND sg13g2_mux2_1
XFILLER_39_475 VPWR VGND sg13g2_decap_8
XFILLER_22_320 VPWR VGND sg13g2_fill_1
XFILLER_34_191 VPWR VGND sg13g2_fill_2
X_5818_ _3078_ VPWR _0403_ VGND net1308 _2786_ sg13g2_o21ai_1
XFILLER_41_36 VPWR VGND sg13g2_decap_4
X_5749_ net1344 _0328_ _0329_ _0026_ VPWR VGND sg13g2_nor3_1
XFILLER_2_714 VPWR VGND sg13g2_decap_8
XFILLER_1_246 VPWR VGND sg13g2_decap_8
X_6568__275 VPWR VGND net275 sg13g2_tiehi
XFILLER_18_604 VPWR VGND sg13g2_decap_4
XFILLER_46_946 VPWR VGND sg13g2_decap_8
XFILLER_45_478 VPWR VGND sg13g2_fill_1
XFILLER_17_158 VPWR VGND sg13g2_decap_8
XFILLER_26_692 VPWR VGND sg13g2_fill_1
XFILLER_32_128 VPWR VGND sg13g2_fill_2
XFILLER_40_194 VPWR VGND sg13g2_fill_1
X_6575__268 VPWR VGND net268 sg13g2_tiehi
Xoutput1 net1 uio_out[2] VPWR VGND sg13g2_buf_1
XFILLER_49_751 VPWR VGND sg13g2_decap_8
X_4080_ _1627_ net1141 _1626_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_489 VPWR VGND sg13g2_decap_4
X_4982_ net1358 _2376_ _2443_ VPWR VGND sg13g2_nor2_1
X_3933_ VGND VPWR net1184 _1496_ _1499_ _1498_ sg13g2_a21oi_1
X_6721_ net110 VGND VPWR _0231_ s0.data_out\[5\]\[3\] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_6652_ net184 VGND VPWR _0162_ s0.data_new_delayed\[3\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_3864_ _1436_ VPWR _1437_ VGND _2744_ _1435_ sg13g2_o21ai_1
X_5603_ _0010_ _3001_ _3002_ _2767_ net1339 VPWR VGND sg13g2_a22oi_1
X_6583_ net259 VGND VPWR net526 s0.data_out\[16\]\[4\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3795_ _1374_ net1188 net451 VPWR VGND sg13g2_nand2_1
X_5534_ net438 net1327 _2940_ VPWR VGND sg13g2_nor2b_1
XFILLER_11_28 VPWR VGND sg13g2_fill_1
XFILLER_11_39 VPWR VGND sg13g2_fill_2
X_5465_ VPWR _2883_ net514 VGND sg13g2_inv_1
X_4416_ VGND VPWR net1086 _1925_ _1927_ _1926_ sg13g2_a21oi_1
X_5396_ VPWR _2814_ net561 VGND sg13g2_inv_1
XFILLER_28_1011 VPWR VGND sg13g2_decap_8
X_4347_ _1867_ VPWR _1870_ VGND net1441 _1830_ sg13g2_o21ai_1
X_4278_ s0.data_out\[8\]\[2\] s0.data_out\[7\]\[2\] net1105 _1801_ VPWR VGND sg13g2_mux2_1
XFILLER_39_261 VPWR VGND sg13g2_fill_2
XFILLER_39_250 VPWR VGND sg13g2_decap_8
X_6017_ net1265 net1173 _0578_ VPWR VGND sg13g2_nor2b_1
XFILLER_43_949 VPWR VGND sg13g2_decap_8
XFILLER_15_629 VPWR VGND sg13g2_fill_1
XFILLER_10_301 VPWR VGND sg13g2_fill_1
XFILLER_11_879 VPWR VGND sg13g2_decap_4
XFILLER_10_389 VPWR VGND sg13g2_fill_1
Xhold390 s0.shift_out\[1\][0] VPWR VGND net710 sg13g2_dlygate4sd3_1
XFILLER_2_588 VPWR VGND sg13g2_fill_1
XFILLER_2_577 VPWR VGND sg13g2_decap_8
XFILLER_46_721 VPWR VGND sg13g2_fill_1
XFILLER_18_412 VPWR VGND sg13g2_decap_8
X_6581__261 VPWR VGND net261 sg13g2_tiehi
XFILLER_19_979 VPWR VGND sg13g2_decap_8
XFILLER_34_949 VPWR VGND sg13g2_decap_8
XFILLER_42_971 VPWR VGND sg13g2_decap_8
XFILLER_14_684 VPWR VGND sg13g2_fill_1
XFILLER_42_90 VPWR VGND sg13g2_decap_4
X_3580_ _1181_ VPWR _1182_ VGND net1017 _1179_ sg13g2_o21ai_1
X_5250_ VGND VPWR net1022 net361 _2681_ _2614_ sg13g2_a21oi_1
X_4201_ _1734_ _1735_ _1736_ VPWR VGND sg13g2_nor2_1
X_5181_ net1022 net1147 _2620_ VPWR VGND sg13g2_nor2b_1
X_4132_ net1139 VPWR _1672_ VGND _1614_ _1671_ sg13g2_o21ai_1
X_4063_ VGND VPWR _1486_ _1609_ _1610_ net1138 sg13g2_a21oi_1
XFILLER_37_721 VPWR VGND sg13g2_fill_2
XFILLER_3_1013 VPWR VGND sg13g2_decap_8
XFILLER_40_919 VPWR VGND sg13g2_decap_4
XFILLER_40_908 VPWR VGND sg13g2_decap_8
X_4965_ _2428_ net1428 _2427_ VPWR VGND sg13g2_nand2_1
X_6704_ net128 VGND VPWR _0214_ s0.genblk1\[5\].modules.bubble clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_3916_ VGND VPWR _1362_ _1481_ _1482_ net1181 sg13g2_a21oi_1
XFILLER_33_993 VPWR VGND sg13g2_decap_8
X_4896_ _2360_ _2361_ _2362_ VPWR VGND sg13g2_nor2_1
XFILLER_20_610 VPWR VGND sg13g2_decap_8
XFILLER_32_481 VPWR VGND sg13g2_fill_1
X_3847_ _0137_ _1422_ _1423_ _2833_ net1378 VPWR VGND sg13g2_a22oi_1
X_6635_ net202 VGND VPWR _0145_ s0.valid_out\[11\][0] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_6566_ net277 VGND VPWR _0076_ s0.shift_out\[17\][0] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3778_ _1357_ net1016 _1356_ VPWR VGND sg13g2_nand2_1
X_5517_ _2923_ net1321 net603 VPWR VGND sg13g2_nand2_1
XFILLER_3_319 VPWR VGND sg13g2_fill_2
X_6497_ net56 VGND VPWR net413 s0.data_out\[23\]\[2\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5448_ VPWR _2866_ net549 VGND sg13g2_inv_1
Xfanout1109 s0.valid_out\[7\][0] net1109 VPWR VGND sg13g2_buf_2
X_5379_ VPWR _2797_ net499 VGND sg13g2_inv_1
XFILLER_47_57 VPWR VGND sg13g2_fill_2
X_6565__278 VPWR VGND net278 sg13g2_tiehi
XFILLER_28_710 VPWR VGND sg13g2_decap_8
XFILLER_30_407 VPWR VGND sg13g2_decap_4
XFILLER_30_418 VPWR VGND sg13g2_fill_1
XFILLER_11_676 VPWR VGND sg13g2_fill_1
XFILLER_12_60 VPWR VGND sg13g2_fill_1
XFILLER_3_831 VPWR VGND sg13g2_decap_8
XFILLER_19_765 VPWR VGND sg13g2_fill_2
XFILLER_33_201 VPWR VGND sg13g2_fill_1
XFILLER_34_735 VPWR VGND sg13g2_fill_2
XFILLER_15_971 VPWR VGND sg13g2_decap_8
X_4750_ net1065 s0.data_out\[4\]\[5\] _2231_ VPWR VGND sg13g2_and2_1
X_6756__72 VPWR VGND net72 sg13g2_tiehi
X_3701_ _1291_ _1282_ _1290_ VPWR VGND sg13g2_nand2_1
X_4681_ _2167_ VPWR _2168_ VGND _2163_ _2164_ sg13g2_o21ai_1
X_6420_ _0945_ net1233 s0.data_out\[15\]\[4\] VPWR VGND sg13g2_nand2_1
X_3632_ _1223_ _1224_ _1225_ VPWR VGND sg13g2_nor2_1
XFILLER_30_996 VPWR VGND sg13g2_decap_8
X_6351_ VPWR _0083_ net665 VGND sg13g2_inv_1
XFILLER_6_680 VPWR VGND sg13g2_fill_2
X_3563_ VGND VPWR _1165_ _1154_ net1404 sg13g2_or2_1
X_5302_ VGND VPWR net1464 _2702_ _0291_ _2724_ sg13g2_a21oi_1
XFILLER_45_0 VPWR VGND sg13g2_fill_1
X_3494_ _1100_ net1485 _1101_ VPWR VGND _1048_ sg13g2_nand3b_1
X_6282_ VGND VPWR net1250 _0816_ _0819_ _0818_ sg13g2_a21oi_1
X_5233_ _2667_ VPWR _2668_ VGND net1465 net541 sg13g2_o21ai_1
X_5164_ _2601_ VPWR _2603_ VGND net1443 _2588_ sg13g2_o21ai_1
X_4115_ _1658_ VPWR _1659_ VGND net1488 net674 sg13g2_o21ai_1
X_5095_ VGND VPWR _2540_ _2544_ _0263_ _2545_ sg13g2_a21oi_1
X_4046_ s0.data_out\[10\]\[3\] s0.data_out\[9\]\[3\] net1133 _1593_ VPWR VGND sg13g2_mux2_1
X_5997_ net1470 VPWR _0561_ VGND _0558_ _0560_ sg13g2_o21ai_1
XFILLER_40_738 VPWR VGND sg13g2_decap_4
X_4948_ VGND VPWR _2411_ _2401_ net1400 sg13g2_or2_1
X_4879_ VPWR _0245_ _2347_ VGND sg13g2_inv_1
XFILLER_20_440 VPWR VGND sg13g2_decap_4
X_6618_ net221 VGND VPWR net533 s0.data_out\[13\]\[3\] clknet_leaf_28_clk sg13g2_dfrbpq_2
XFILLER_21_985 VPWR VGND sg13g2_decap_8
X_6549_ net296 VGND VPWR _0059_ s0.data_out\[19\]\[6\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_0_845 VPWR VGND sg13g2_decap_8
XFILLER_48_816 VPWR VGND sg13g2_decap_8
XFILLER_15_201 VPWR VGND sg13g2_decap_4
XFILLER_43_543 VPWR VGND sg13g2_fill_1
XFILLER_43_554 VPWR VGND sg13g2_fill_1
XFILLER_30_215 VPWR VGND sg13g2_fill_1
XFILLER_30_226 VPWR VGND sg13g2_decap_4
XFILLER_8_912 VPWR VGND sg13g2_decap_8
XFILLER_30_248 VPWR VGND sg13g2_decap_8
XFILLER_12_996 VPWR VGND sg13g2_decap_8
X_6753__75 VPWR VGND net75 sg13g2_tiehi
XFILLER_8_989 VPWR VGND sg13g2_decap_8
XFILLER_11_495 VPWR VGND sg13g2_fill_2
XFILLER_39_816 VPWR VGND sg13g2_fill_1
Xfanout1440 net1441 net1440 VPWR VGND sg13g2_buf_8
Xfanout1473 net1475 net1473 VPWR VGND sg13g2_buf_8
Xfanout1462 net1463 net1462 VPWR VGND sg13g2_buf_8
Xfanout1484 net1487 net1484 VPWR VGND sg13g2_buf_8
Xfanout1451 net1457 net1451 VPWR VGND sg13g2_buf_8
XFILLER_47_871 VPWR VGND sg13g2_decap_8
X_5920_ _0493_ net1282 net622 VPWR VGND sg13g2_nand2_1
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
XFILLER_19_584 VPWR VGND sg13g2_fill_2
XFILLER_34_532 VPWR VGND sg13g2_fill_1
X_5851_ VGND VPWR net1008 _0395_ _0431_ net1344 sg13g2_a21oi_1
XFILLER_15_790 VPWR VGND sg13g2_fill_2
X_5782_ net1451 _0342_ _0367_ VPWR VGND sg13g2_nor2_1
X_4802_ _2275_ net1050 _2276_ _2277_ VPWR VGND sg13g2_a21o_1
X_4733_ net1072 VPWR _2218_ VGND _2136_ _2217_ sg13g2_o21ai_1
XFILLER_30_793 VPWR VGND sg13g2_fill_1
X_6403_ _0926_ net1223 _0927_ _0928_ VPWR VGND sg13g2_a21o_1
X_4664_ VGND VPWR net1061 _2149_ _2151_ _2150_ sg13g2_a21oi_1
X_4595_ _2094_ _2093_ _2073_ VPWR VGND sg13g2_nand2b_1
X_3615_ VPWR _0118_ net685 VGND sg13g2_inv_1
X_3546_ _1148_ net1211 net406 VPWR VGND sg13g2_nand2_1
X_6334_ net1239 net482 _0867_ VPWR VGND sg13g2_and2_1
X_6265_ _0788_ VPWR _0802_ VGND net1453 _0795_ sg13g2_o21ai_1
X_3477_ net1367 _1009_ _1088_ VPWR VGND sg13g2_nor2_1
X_5216_ VGND VPWR net1020 net547 _2654_ _2598_ sg13g2_a21oi_1
X_6196_ _0665_ _0743_ _0744_ _0745_ VPWR VGND sg13g2_nor3_1
X_5147_ VGND VPWR net1020 _2584_ _2586_ _2585_ sg13g2_a21oi_1
XFILLER_28_15 VPWR VGND sg13g2_fill_1
X_5078_ s0.data_out\[2\]\[5\] s0.data_out\[1\]\[5\] net1035 _2529_ VPWR VGND sg13g2_mux2_1
X_4029_ _1576_ net1014 _1575_ VPWR VGND sg13g2_nand2_1
XFILLER_40_513 VPWR VGND sg13g2_fill_2
XFILLER_40_579 VPWR VGND sg13g2_fill_2
XFILLER_5_948 VPWR VGND sg13g2_decap_8
XFILLER_0_642 VPWR VGND sg13g2_decap_8
XFILLER_44_863 VPWR VGND sg13g2_decap_4
XFILLER_43_362 VPWR VGND sg13g2_fill_2
XFILLER_15_1013 VPWR VGND sg13g2_decap_8
XFILLER_7_230 VPWR VGND sg13g2_fill_2
XFILLER_11_292 VPWR VGND sg13g2_fill_1
XFILLER_12_793 VPWR VGND sg13g2_fill_1
Xhold208 _0324_ VPWR VGND net528 sg13g2_dlygate4sd3_1
X_4380_ _1895_ net1481 _1896_ VPWR VGND _1838_ sg13g2_nand3b_1
Xhold219 s0.valid_out\[21\][0] VPWR VGND net539 sg13g2_dlygate4sd3_1
X_3400_ _1013_ VPWR _1014_ VGND net1220 _2818_ sg13g2_o21ai_1
XFILLER_4_992 VPWR VGND sg13g2_decap_8
X_6050_ VPWR _0611_ _0610_ VGND sg13g2_inv_1
X_5001_ net1052 VPWR _2457_ VGND _2404_ _2456_ sg13g2_o21ai_1
X_6626__212 VPWR VGND net212 sg13g2_tiehi
XFILLER_39_657 VPWR VGND sg13g2_decap_8
XFILLER_39_646 VPWR VGND sg13g2_fill_1
Xfanout1281 net1285 net1281 VPWR VGND sg13g2_buf_8
Xfanout1292 s0.shift_out\[20\][0] net1292 VPWR VGND sg13g2_buf_1
Xfanout1270 net1272 net1270 VPWR VGND sg13g2_buf_8
XFILLER_26_329 VPWR VGND sg13g2_decap_4
X_5903_ _0461_ VPWR _0476_ VGND net1451 _0468_ sg13g2_o21ai_1
X_5834_ _0344_ _0417_ net1462 _0418_ VPWR VGND sg13g2_nand3_1
XFILLER_10_708 VPWR VGND sg13g2_fill_2
XFILLER_10_719 VPWR VGND sg13g2_fill_1
X_5765_ net1291 net1163 _0350_ VPWR VGND sg13g2_nor2b_1
X_4716_ _2203_ _2194_ _2202_ VPWR VGND sg13g2_nand2_1
X_5696_ _3051_ _3069_ _3086_ _3089_ _3090_ VPWR VGND sg13g2_or4_1
X_6633__205 VPWR VGND net205 sg13g2_tiehi
XFILLER_30_27 VPWR VGND sg13g2_fill_2
X_4647_ _2134_ net1067 net642 VPWR VGND sg13g2_nand2_1
X_4578_ _2077_ net1090 _2076_ VPWR VGND sg13g2_nand2b_1
X_6317_ _0840_ VPWR _0854_ VGND _0848_ _0850_ sg13g2_o21ai_1
XFILLER_39_14 VPWR VGND sg13g2_decap_8
X_3529_ s0.data_out\[14\]\[0\] s0.data_out\[13\]\[0\] net1210 _1131_ VPWR VGND sg13g2_mux2_1
X_6248_ _0785_ net426 net1259 VPWR VGND sg13g2_nand2b_1
XFILLER_39_58 VPWR VGND sg13g2_fill_2
X_6179_ VGND VPWR net1268 _0725_ _0728_ _0727_ sg13g2_a21oi_1
XFILLER_5_734 VPWR VGND sg13g2_fill_2
XFILLER_4_244 VPWR VGND sg13g2_fill_2
XFILLER_20_82 VPWR VGND sg13g2_decap_8
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_940 VPWR VGND sg13g2_decap_8
XFILLER_49_933 VPWR VGND sg13g2_decap_8
Xhold91 _0068_ VPWR VGND net411 sg13g2_dlygate4sd3_1
Xhold80 s0.data_out\[3\]\[1\] VPWR VGND net400 sg13g2_dlygate4sd3_1
XFILLER_43_181 VPWR VGND sg13g2_fill_2
XFILLER_16_395 VPWR VGND sg13g2_fill_1
X_3880_ VGND VPWR _1450_ _1449_ _1447_ sg13g2_or2_1
X_5550_ _2956_ _2955_ net1407 _2947_ net1398 VPWR VGND sg13g2_a22oi_1
X_4501_ net998 _2861_ _2005_ VPWR VGND sg13g2_nor2_1
X_5481_ _2892_ VPWR net8 VGND _2766_ net991 sg13g2_o21ai_1
X_4432_ s0.data_out\[7\]\[6\] s0.data_out\[6\]\[6\] net1094 _1943_ VPWR VGND sg13g2_mux2_1
XFILLER_6_73 VPWR VGND sg13g2_decap_4
XFILLER_6_62 VPWR VGND sg13g2_decap_8
X_4363_ net1110 VPWR _1883_ VGND _1802_ _1882_ sg13g2_o21ai_1
X_6102_ net1274 VPWR _0656_ VGND _0603_ _0655_ sg13g2_o21ai_1
X_4294_ net1098 net1171 _1817_ VPWR VGND sg13g2_nor2b_1
X_6033_ _0594_ net1269 net499 VPWR VGND sg13g2_nand2_1
XFILLER_39_421 VPWR VGND sg13g2_fill_2
XFILLER_35_693 VPWR VGND sg13g2_fill_2
XFILLER_22_310 VPWR VGND sg13g2_decap_4
XFILLER_23_811 VPWR VGND sg13g2_decap_8
XFILLER_23_833 VPWR VGND sg13g2_decap_4
X_5817_ _0402_ net1302 _0401_ VPWR VGND sg13g2_nand2b_1
X_5748_ _0025_ net1462 _0331_ _0335_ VPWR VGND sg13g2_and3_1
X_5679_ VGND VPWR net1304 _3072_ _3073_ _3070_ sg13g2_a21oi_1
XFILLER_46_925 VPWR VGND sg13g2_decap_8
XFILLER_14_811 VPWR VGND sg13g2_fill_1
XFILLER_41_685 VPWR VGND sg13g2_fill_1
XFILLER_14_888 VPWR VGND sg13g2_fill_2
XFILLER_15_71 VPWR VGND sg13g2_decap_4
XFILLER_13_387 VPWR VGND sg13g2_fill_2
XFILLER_31_81 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
Xoutput2 net2 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_49_730 VPWR VGND sg13g2_decap_8
XFILLER_36_468 VPWR VGND sg13g2_fill_1
XFILLER_36_457 VPWR VGND sg13g2_decap_8
XFILLER_45_991 VPWR VGND sg13g2_decap_8
XFILLER_17_671 VPWR VGND sg13g2_fill_1
X_4981_ net1047 VPWR _2442_ VGND _2373_ _2441_ sg13g2_o21ai_1
X_3932_ VGND VPWR _1381_ _1497_ _1498_ net1184 sg13g2_a21oi_1
X_6720_ net111 VGND VPWR _0230_ s0.data_out\[5\]\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_6651_ net185 VGND VPWR _0161_ s0.data_new_delayed\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_3863_ VGND VPWR _2744_ _1404_ _1436_ net1386 sg13g2_a21oi_1
X_5602_ net1339 _2969_ _3002_ VPWR VGND sg13g2_nor2_1
X_6582_ net260 VGND VPWR net483 s0.data_out\[16\]\[3\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_20_836 VPWR VGND sg13g2_fill_2
X_5533_ VPWR _2939_ _2938_ VGND sg13g2_inv_1
XFILLER_20_869 VPWR VGND sg13g2_decap_4
X_3794_ _1370_ _1372_ _1373_ VPWR VGND sg13g2_nor2_1
X_6630__208 VPWR VGND net208 sg13g2_tiehi
X_5464_ VPWR _2882_ net463 VGND sg13g2_inv_1
X_5395_ VPWR _2813_ net479 VGND sg13g2_inv_1
X_4415_ net1086 net1172 _1926_ VPWR VGND sg13g2_nor2b_1
X_4346_ _1860_ VPWR _1869_ VGND net1431 _1866_ sg13g2_o21ai_1
X_4277_ _1800_ net1105 net453 VPWR VGND sg13g2_nand2_1
X_6016_ s0.data_out\[19\]\[0\] s0.data_out\[18\]\[0\] net1270 _0577_ VPWR VGND sg13g2_mux2_1
XFILLER_28_969 VPWR VGND sg13g2_decap_8
XFILLER_43_928 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_34_clk clknet_3_4__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_35_1016 VPWR VGND sg13g2_decap_8
XFILLER_22_151 VPWR VGND sg13g2_fill_2
XFILLER_23_663 VPWR VGND sg13g2_fill_1
XFILLER_23_685 VPWR VGND sg13g2_fill_1
XFILLER_10_335 VPWR VGND sg13g2_fill_1
XFILLER_11_869 VPWR VGND sg13g2_decap_4
Xhold380 s0.data_new_delayed\[2\] VPWR VGND net700 sg13g2_dlygate4sd3_1
Xhold391 s0.valid_out\[5\][0] VPWR VGND net711 sg13g2_dlygate4sd3_1
XFILLER_19_925 VPWR VGND sg13g2_fill_2
XFILLER_45_210 VPWR VGND sg13g2_decap_8
XFILLER_18_457 VPWR VGND sg13g2_fill_1
XFILLER_46_799 VPWR VGND sg13g2_decap_8
XFILLER_34_928 VPWR VGND sg13g2_decap_4
XFILLER_42_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_25_clk clknet_3_4__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_9_111 VPWR VGND sg13g2_decap_4
X_6768__306 VPWR VGND net306 sg13g2_tiehi
X_4200_ net1405 _1732_ _1735_ VPWR VGND sg13g2_nor2_1
X_5180_ s0.data_out\[1\]\[6\] s0.data_out\[0\]\[6\] net1025 _2619_ VPWR VGND sg13g2_mux2_1
X_4131_ net1128 net509 _1671_ VPWR VGND sg13g2_and2_1
X_4062_ _1609_ net505 net1175 VPWR VGND sg13g2_nand2b_1
XFILLER_37_711 VPWR VGND sg13g2_fill_1
XFILLER_18_980 VPWR VGND sg13g2_decap_8
X_4964_ VGND VPWR net1051 _2424_ _2427_ _2426_ sg13g2_a21oi_1
XFILLER_24_438 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_16_clk clknet_3_6__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_6703_ net129 VGND VPWR _0213_ s0.valid_out\[6\][0] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_3915_ _1481_ s0.data_out\[10\]\[3\] net1190 VPWR VGND sg13g2_nand2b_1
XFILLER_33_972 VPWR VGND sg13g2_decap_8
X_4895_ VGND VPWR _2729_ _2748_ _2361_ net1051 sg13g2_a21oi_1
X_6558__286 VPWR VGND net286 sg13g2_tiehi
X_3846_ net1379 _1343_ _1423_ VPWR VGND sg13g2_nor2_1
XFILLER_22_17 VPWR VGND sg13g2_fill_1
X_6634_ net204 VGND VPWR net645 s0.was_valid_out\[11\][0] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_6565_ net278 VGND VPWR _0075_ s0.genblk1\[16\].modules.bubble clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_3777_ s0.data_out\[11\]\[2\] s0.data_out\[12\]\[2\] net1200 _1356_ VPWR VGND sg13g2_mux2_1
X_6496_ net57 VGND VPWR net382 s0.data_out\[23\]\[1\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5516_ VGND VPWR net1328 _2778_ _2922_ _2921_ sg13g2_a21oi_1
X_5447_ VPWR _2865_ net656 VGND sg13g2_inv_1
X_5378_ VPWR _2796_ net695 VGND sg13g2_inv_1
X_4329_ _1848_ _1849_ _1847_ _1852_ VPWR VGND sg13g2_nand3_1
XFILLER_47_25 VPWR VGND sg13g2_decap_8
XFILLER_27_210 VPWR VGND sg13g2_fill_1
XFILLER_28_755 VPWR VGND sg13g2_fill_2
XFILLER_11_611 VPWR VGND sg13g2_decap_8
XFILLER_7_604 VPWR VGND sg13g2_fill_2
XFILLER_10_143 VPWR VGND sg13g2_decap_8
XFILLER_7_626 VPWR VGND sg13g2_fill_1
XFILLER_6_103 VPWR VGND sg13g2_fill_1
XFILLER_12_72 VPWR VGND sg13g2_fill_2
XFILLER_3_810 VPWR VGND sg13g2_decap_8
XFILLER_3_887 VPWR VGND sg13g2_decap_8
XFILLER_18_243 VPWR VGND sg13g2_decap_8
XFILLER_19_744 VPWR VGND sg13g2_decap_8
XFILLER_19_788 VPWR VGND sg13g2_fill_2
XFILLER_33_235 VPWR VGND sg13g2_decap_8
XFILLER_18_1022 VPWR VGND sg13g2_decap_8
X_3700_ _1290_ net1432 _1289_ VPWR VGND sg13g2_nand2_1
XFILLER_30_975 VPWR VGND sg13g2_decap_8
X_4680_ _2167_ net1439 _2162_ VPWR VGND sg13g2_nand2_1
X_3631_ VGND VPWR _2734_ _2740_ _1224_ net1208 sg13g2_a21oi_1
X_6350_ _0879_ VPWR _0880_ VGND net1478 net664 sg13g2_o21ai_1
X_3562_ VGND VPWR _1164_ _1161_ net1413 sg13g2_or2_1
X_5301_ net1464 net402 _2724_ VPWR VGND sg13g2_nor2_1
X_6281_ VGND VPWR _0704_ _0817_ _0818_ net1250 sg13g2_a21oi_1
X_3493_ net1229 VPWR _1100_ VGND _1045_ _1099_ sg13g2_o21ai_1
Xclkbuf_leaf_5_clk clknet_3_4__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_5232_ _2666_ VPWR _2667_ VGND net1005 _2665_ sg13g2_o21ai_1
XFILLER_38_0 VPWR VGND sg13g2_fill_2
XFILLER_25_1015 VPWR VGND sg13g2_decap_8
X_5163_ VPWR VGND _2600_ net1458 _2596_ net1449 _2602_ _2594_ sg13g2_a221oi_1
XFILLER_29_508 VPWR VGND sg13g2_fill_1
X_4114_ _1657_ VPWR _1658_ VGND net1014 _1656_ sg13g2_o21ai_1
X_5094_ VGND VPWR _2545_ net1329 net334 sg13g2_or2_1
X_4045_ _1592_ net1131 net589 VPWR VGND sg13g2_nand2_1
XFILLER_40_706 VPWR VGND sg13g2_decap_4
X_5996_ _0560_ _0557_ _0559_ VPWR VGND sg13g2_nand2_1
X_4947_ net1409 _2408_ _2410_ VPWR VGND sg13g2_nor2_1
X_4878_ _2346_ VPWR _2347_ VGND net1473 net681 sg13g2_o21ai_1
XFILLER_21_964 VPWR VGND sg13g2_decap_8
X_6617_ net222 VGND VPWR net458 s0.data_out\[13\]\[2\] clknet_leaf_28_clk sg13g2_dfrbpq_2
XFILLER_20_463 VPWR VGND sg13g2_decap_8
XFILLER_20_485 VPWR VGND sg13g2_fill_2
X_3829_ VGND VPWR _1396_ _1398_ _1408_ net1432 sg13g2_a21oi_1
X_6548_ net297 VGND VPWR _0058_ s0.data_out\[19\]\[5\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_6571__272 VPWR VGND net272 sg13g2_tiehi
X_6479_ net1395 net1221 _0995_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_824 VPWR VGND sg13g2_decap_8
XFILLER_47_316 VPWR VGND sg13g2_fill_1
XFILLER_16_714 VPWR VGND sg13g2_fill_1
XFILLER_15_235 VPWR VGND sg13g2_fill_2
XFILLER_16_758 VPWR VGND sg13g2_decap_8
XFILLER_12_920 VPWR VGND sg13g2_fill_2
XFILLER_11_463 VPWR VGND sg13g2_fill_2
XFILLER_12_975 VPWR VGND sg13g2_decap_8
XFILLER_23_82 VPWR VGND sg13g2_decap_8
XFILLER_8_968 VPWR VGND sg13g2_decap_8
XFILLER_48_1026 VPWR VGND sg13g2_fill_2
XFILLER_3_684 VPWR VGND sg13g2_decap_8
Xfanout1441 net1442 net1441 VPWR VGND sg13g2_buf_8
Xfanout1430 net1434 net1430 VPWR VGND sg13g2_buf_8
XFILLER_2_194 VPWR VGND sg13g2_fill_2
Xfanout1474 net1475 net1474 VPWR VGND sg13g2_buf_8
XFILLER_38_305 VPWR VGND sg13g2_decap_8
Xfanout1463 net1476 net1463 VPWR VGND sg13g2_buf_8
Xfanout1452 net1457 net1452 VPWR VGND sg13g2_buf_8
XFILLER_47_850 VPWR VGND sg13g2_decap_8
XFILLER_48_90 VPWR VGND sg13g2_decap_4
XFILLER_19_541 VPWR VGND sg13g2_fill_1
Xfanout1485 net1487 net1485 VPWR VGND sg13g2_buf_8
XFILLER_0_1006 VPWR VGND sg13g2_decap_8
X_5850_ VGND VPWR net1292 net496 _0430_ _0390_ sg13g2_a21oi_1
XFILLER_15_780 VPWR VGND sg13g2_fill_2
X_5781_ net1437 _0365_ _0366_ VPWR VGND sg13g2_nor2_1
XFILLER_21_205 VPWR VGND sg13g2_decap_4
X_4801_ net1050 net1161 _2276_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_588 VPWR VGND sg13g2_fill_1
X_4732_ net995 _2873_ _2217_ VPWR VGND sg13g2_nor2_1
XFILLER_9_73 VPWR VGND sg13g2_fill_2
X_4663_ net1061 net1163 _2150_ VPWR VGND sg13g2_nor2b_1
X_3614_ _1209_ VPWR _1210_ VGND net1485 net684 sg13g2_o21ai_1
X_6402_ net1223 net1149 _0927_ VPWR VGND sg13g2_nor2b_1
X_4594_ _2087_ VPWR _2093_ VGND _2080_ _2090_ sg13g2_o21ai_1
X_6555__289 VPWR VGND net289 sg13g2_tiehi
X_6333_ _0079_ _0865_ _0866_ _2806_ net1366 VPWR VGND sg13g2_a22oi_1
X_3545_ _1146_ VPWR _1147_ VGND _1137_ _1138_ sg13g2_o21ai_1
X_3476_ net1227 VPWR _1087_ VGND _1006_ _1086_ sg13g2_o21ai_1
X_6264_ _0801_ _2757_ _0800_ VPWR VGND sg13g2_nand2_1
X_5215_ net325 net1329 _2653_ _0275_ VPWR VGND sg13g2_nor3_1
X_6195_ _0718_ _0720_ _0744_ VPWR VGND sg13g2_nor2b_1
X_5146_ net1019 net1162 _2585_ VPWR VGND sg13g2_nor2b_1
X_5077_ _2525_ _2527_ net1426 _2528_ VPWR VGND sg13g2_nand3_1
XFILLER_38_883 VPWR VGND sg13g2_fill_2
X_4028_ s0.data_out\[9\]\[0\] s0.data_out\[10\]\[0\] net1174 _1575_ VPWR VGND sg13g2_mux2_1
XFILLER_40_503 VPWR VGND sg13g2_decap_4
X_5979_ net1352 net353 _0546_ VPWR VGND sg13g2_nor2_1
XFILLER_21_794 VPWR VGND sg13g2_decap_8
XFILLER_5_927 VPWR VGND sg13g2_decap_8
X_6750__79 VPWR VGND net79 sg13g2_tiehi
XFILLER_0_621 VPWR VGND sg13g2_decap_8
XFILLER_0_698 VPWR VGND sg13g2_decap_8
XFILLER_48_669 VPWR VGND sg13g2_decap_8
XFILLER_44_897 VPWR VGND sg13g2_decap_8
XFILLER_43_374 VPWR VGND sg13g2_fill_2
XFILLER_16_599 VPWR VGND sg13g2_decap_8
X_6619__220 VPWR VGND net220 sg13g2_tiehi
Xhold209 s0.data_out\[17\]\[1\] VPWR VGND net529 sg13g2_dlygate4sd3_1
XFILLER_4_971 VPWR VGND sg13g2_decap_8
X_5000_ net1010 _2881_ _2456_ VPWR VGND sg13g2_nor2_1
XFILLER_39_636 VPWR VGND sg13g2_fill_1
XFILLER_39_614 VPWR VGND sg13g2_fill_1
Xfanout1282 net1285 net1282 VPWR VGND sg13g2_buf_1
Xfanout1271 net1272 net1271 VPWR VGND sg13g2_buf_1
Xfanout1260 s0.valid_out\[17\][0] net1260 VPWR VGND sg13g2_buf_1
XFILLER_38_168 VPWR VGND sg13g2_fill_1
XFILLER_38_157 VPWR VGND sg13g2_decap_4
Xfanout1293 net1295 net1293 VPWR VGND sg13g2_buf_8
XFILLER_19_393 VPWR VGND sg13g2_fill_1
X_5902_ VPWR VGND _0474_ net1461 _0472_ net1451 _0475_ _0468_ sg13g2_a221oi_1
X_5833_ net1305 VPWR _0417_ VGND _0345_ _0416_ sg13g2_o21ai_1
X_5764_ VPWR VGND _0348_ net1461 _0344_ net1451 _0349_ _0342_ sg13g2_a221oi_1
X_4715_ _2199_ _2201_ net1418 _2202_ VPWR VGND sg13g2_nand3_1
X_5695_ VGND VPWR _3089_ _3088_ _3087_ sg13g2_or2_1
X_4646_ net1475 net321 _0226_ VPWR VGND sg13g2_and2_1
X_4577_ VGND VPWR net1075 _2075_ _2076_ _2074_ sg13g2_a21oi_1
X_6316_ _0832_ _0850_ _0851_ _0852_ _0853_ VPWR VGND sg13g2_nor4_1
X_3528_ VGND VPWR net1214 _1127_ _1130_ _1129_ sg13g2_a21oi_1
X_3459_ _1071_ VPWR _1073_ VGND net1440 _1033_ sg13g2_o21ai_1
X_6247_ _0782_ net1238 _0783_ _0784_ VPWR VGND sg13g2_a21o_1
X_6178_ VGND VPWR _0613_ _0726_ _0727_ net1268 sg13g2_a21oi_1
X_5129_ net1041 VPWR _2572_ VGND _2507_ _2571_ sg13g2_o21ai_1
XFILLER_17_319 VPWR VGND sg13g2_fill_1
XFILLER_44_116 VPWR VGND sg13g2_fill_2
XFILLER_44_105 VPWR VGND sg13g2_decap_8
XFILLER_41_856 VPWR VGND sg13g2_fill_1
XFILLER_40_399 VPWR VGND sg13g2_fill_2
XFILLER_20_50 VPWR VGND sg13g2_decap_4
XFILLER_49_912 VPWR VGND sg13g2_decap_8
XFILLER_1_996 VPWR VGND sg13g2_decap_8
XFILLER_0_495 VPWR VGND sg13g2_decap_8
XFILLER_49_989 VPWR VGND sg13g2_decap_8
XFILLER_48_466 VPWR VGND sg13g2_fill_1
Xhold92 s0.data_out\[23\]\[2\] VPWR VGND net412 sg13g2_dlygate4sd3_1
Xhold81 _0253_ VPWR VGND net401 sg13g2_dlygate4sd3_1
Xhold70 _1939_ VPWR VGND net390 sg13g2_dlygate4sd3_1
XFILLER_35_127 VPWR VGND sg13g2_fill_2
XFILLER_16_330 VPWR VGND sg13g2_decap_4
XFILLER_32_856 VPWR VGND sg13g2_fill_1
X_4500_ _0209_ _2003_ _2004_ _2856_ net1372 VPWR VGND sg13g2_a22oi_1
X_5480_ _2892_ net1407 net991 VPWR VGND sg13g2_nand2_1
X_4431_ _1942_ net1094 net578 VPWR VGND sg13g2_nand2_1
X_4362_ net1098 net453 _1882_ VPWR VGND sg13g2_and2_1
XFILLER_4_790 VPWR VGND sg13g2_fill_2
X_6101_ net1261 s0.data_out\[18\]\[6\] _0655_ VPWR VGND sg13g2_and2_1
X_4293_ _1815_ VPWR _1816_ VGND net1106 _2854_ sg13g2_o21ai_1
XFILLER_6_1012 VPWR VGND sg13g2_decap_8
X_6032_ _0592_ VPWR _0593_ VGND _0583_ _0584_ sg13g2_o21ai_1
Xfanout1090 net1091 net1090 VPWR VGND sg13g2_buf_8
XFILLER_41_108 VPWR VGND sg13g2_decap_4
X_5816_ VGND VPWR net1289 _0399_ _0401_ _0400_ sg13g2_a21oi_1
XFILLER_22_355 VPWR VGND sg13g2_decap_4
X_5747_ _0333_ _0334_ _0332_ _0335_ VPWR VGND sg13g2_nand3_1
X_5678_ s0.data_out\[22\]\[4\] s0.data_out\[21\]\[4\] net1307 _3072_ VPWR VGND sg13g2_mux2_1
X_4629_ net1372 _2068_ _2121_ VPWR VGND sg13g2_nor2_1
XFILLER_2_749 VPWR VGND sg13g2_decap_8
XFILLER_49_208 VPWR VGND sg13g2_fill_2
XFILLER_46_904 VPWR VGND sg13g2_decap_8
XFILLER_45_414 VPWR VGND sg13g2_fill_1
XFILLER_45_469 VPWR VGND sg13g2_decap_8
XFILLER_32_108 VPWR VGND sg13g2_fill_2
XFILLER_12_1017 VPWR VGND sg13g2_decap_8
X_6616__223 VPWR VGND net223 sg13g2_tiehi
XFILLER_5_510 VPWR VGND sg13g2_fill_2
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
Xoutput3 net3 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_793 VPWR VGND sg13g2_decap_8
XFILLER_49_786 VPWR VGND sg13g2_decap_8
XFILLER_37_915 VPWR VGND sg13g2_fill_2
XFILLER_37_959 VPWR VGND sg13g2_decap_8
X_6623__216 VPWR VGND net216 sg13g2_tiehi
XFILLER_45_970 VPWR VGND sg13g2_decap_8
X_4980_ net1009 _2883_ _2441_ VPWR VGND sg13g2_nor2_1
X_3931_ _1497_ net636 net1189 VPWR VGND sg13g2_nand2b_1
XFILLER_20_815 VPWR VGND sg13g2_decap_8
X_6650_ net186 VGND VPWR _0160_ s0.data_new_delayed\[1\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_3862_ VGND VPWR net1182 s0.data_out\[11\]\[5\] _1435_ _1401_ sg13g2_a21oi_1
XFILLER_31_141 VPWR VGND sg13g2_fill_1
XFILLER_31_152 VPWR VGND sg13g2_fill_1
X_5601_ net1323 VPWR _3001_ VGND _2971_ _3000_ sg13g2_o21ai_1
X_6581_ net261 VGND VPWR _0091_ s0.data_out\[16\]\[2\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_20_848 VPWR VGND sg13g2_fill_1
XFILLER_32_686 VPWR VGND sg13g2_fill_1
X_5532_ _2938_ _2937_ net1435 _2911_ net1443 VPWR VGND sg13g2_a22oi_1
X_3793_ _1371_ VPWR _1372_ VGND _1359_ _1369_ sg13g2_o21ai_1
X_5463_ VPWR _2881_ net580 VGND sg13g2_inv_1
X_5394_ VPWR _2812_ net426 VGND sg13g2_inv_1
X_4414_ s0.data_out\[7\]\[0\] s0.data_out\[6\]\[0\] net1092 _1925_ VPWR VGND sg13g2_mux2_1
X_4345_ net1422 _1859_ _1868_ VPWR VGND sg13g2_nor2_1
X_4276_ net1480 net344 _0190_ VPWR VGND sg13g2_and2_1
X_6015_ VGND VPWR net1278 _0573_ _0576_ _0575_ sg13g2_a21oi_1
XFILLER_39_285 VPWR VGND sg13g2_decap_4
XFILLER_43_907 VPWR VGND sg13g2_decap_8
XFILLER_11_837 VPWR VGND sg13g2_fill_2
X_6779_ net143 VGND VPWR net376 s0.data_out\[0\]\[1\] clknet_leaf_8_clk sg13g2_dfrbpq_2
XFILLER_7_4 VPWR VGND sg13g2_fill_1
Xhold381 s0.valid_out\[15\][0] VPWR VGND net701 sg13g2_dlygate4sd3_1
Xhold370 s0.data_out\[19\]\[3\] VPWR VGND net690 sg13g2_dlygate4sd3_1
Xhold392 s0.data_new_delayed\[3\] VPWR VGND net712 sg13g2_dlygate4sd3_1
XFILLER_46_778 VPWR VGND sg13g2_decap_8
XFILLER_18_469 VPWR VGND sg13g2_fill_1
XFILLER_33_428 VPWR VGND sg13g2_decap_8
XFILLER_45_299 VPWR VGND sg13g2_fill_2
XFILLER_27_992 VPWR VGND sg13g2_decap_8
XFILLER_13_141 VPWR VGND sg13g2_fill_2
XFILLER_9_134 VPWR VGND sg13g2_fill_1
XFILLER_14_697 VPWR VGND sg13g2_fill_2
XFILLER_5_384 VPWR VGND sg13g2_fill_1
X_4130_ VPWR _0173_ net614 VGND sg13g2_inv_1
X_4061_ _1606_ net1128 _1607_ _1608_ VPWR VGND sg13g2_a21o_1
XFILLER_49_583 VPWR VGND sg13g2_decap_8
XFILLER_36_299 VPWR VGND sg13g2_decap_4
X_4963_ VGND VPWR _2303_ _2425_ _2426_ net1048 sg13g2_a21oi_1
X_6697__136 VPWR VGND net136 sg13g2_tiehi
X_6702_ net131 VGND VPWR _0212_ s0.was_valid_out\[6\][0] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3914_ _1478_ net1137 _1479_ _1480_ VPWR VGND sg13g2_a21o_1
XFILLER_33_951 VPWR VGND sg13g2_decap_8
X_4894_ net1040 _2354_ _2360_ VPWR VGND sg13g2_nor2_1
X_6633_ net205 VGND VPWR _0143_ s0.data_out\[12\]\[7\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_3845_ net1191 VPWR _1422_ VGND _1340_ _1421_ sg13g2_o21ai_1
X_6564_ net279 VGND VPWR _0074_ s0.valid_out\[17\][0] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3776_ VGND VPWR net1180 _1353_ _1355_ _1354_ sg13g2_a21oi_1
X_5515_ _2777_ _2750_ net1325 _2921_ VPWR VGND sg13g2_a21o_1
X_6495_ net58 VGND VPWR net380 s0.data_out\[23\]\[0\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5446_ VPWR _2864_ net692 VGND sg13g2_inv_1
X_5377_ VPWR _2795_ net657 VGND sg13g2_inv_1
X_4328_ _1851_ _1847_ _1848_ _1849_ VPWR VGND sg13g2_and3_1
XFILLER_47_509 VPWR VGND sg13g2_decap_4
X_4259_ net1384 _1724_ _1787_ VPWR VGND sg13g2_nor2_1
XFILLER_24_984 VPWR VGND sg13g2_decap_8
XFILLER_7_638 VPWR VGND sg13g2_fill_2
XFILLER_6_159 VPWR VGND sg13g2_decap_4
X_6613__226 VPWR VGND net226 sg13g2_tiehi
XFILLER_3_866 VPWR VGND sg13g2_decap_8
XFILLER_19_9 VPWR VGND sg13g2_fill_2
XFILLER_46_586 VPWR VGND sg13g2_decap_4
XFILLER_46_597 VPWR VGND sg13g2_fill_2
X_6620__219 VPWR VGND net219 sg13g2_tiehi
XFILLER_18_1001 VPWR VGND sg13g2_decap_8
XFILLER_42_781 VPWR VGND sg13g2_decap_8
XFILLER_30_954 VPWR VGND sg13g2_decap_8
X_3630_ net1196 _1217_ _1223_ VPWR VGND sg13g2_nor2_1
X_3561_ VPWR _1163_ _1162_ VGND sg13g2_inv_1
X_5300_ VGND VPWR net1464 _2696_ _0290_ _2723_ sg13g2_a21oi_1
X_6280_ _0817_ net503 net1257 VPWR VGND sg13g2_nand2b_1
X_3492_ net1017 _2820_ _1099_ VPWR VGND sg13g2_nor2_1
X_5231_ VGND VPWR net1005 _2604_ _2666_ net1346 sg13g2_a21oi_1
X_5162_ VGND VPWR _2601_ _2594_ net1450 sg13g2_or2_1
X_5093_ _2542_ _2543_ _2544_ VPWR VGND sg13g2_nor2_1
X_4113_ VGND VPWR net1014 _1587_ _1657_ net1385 sg13g2_a21oi_1
X_4044_ _1591_ net1335 _1589_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_225 VPWR VGND sg13g2_decap_4
X_5995_ net1003 VPWR _0559_ VGND s0.was_valid_out\[18\][0] net1281 sg13g2_o21ai_1
XFILLER_24_258 VPWR VGND sg13g2_decap_4
X_4946_ _2409_ _2408_ net1409 _2401_ net1400 VPWR VGND sg13g2_a22oi_1
X_4877_ _2345_ VPWR _2346_ VGND net996 _2344_ sg13g2_o21ai_1
X_6616_ net223 VGND VPWR _0126_ s0.data_out\[13\]\[1\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3828_ _1407_ _1399_ _1406_ VPWR VGND sg13g2_nand2_1
X_6762__66 VPWR VGND net66 sg13g2_tiehi
X_6547_ net298 VGND VPWR net487 s0.data_out\[19\]\[4\] clknet_leaf_35_clk sg13g2_dfrbpq_1
XFILLER_4_619 VPWR VGND sg13g2_decap_8
X_3759_ _1338_ net1187 net588 VPWR VGND sg13g2_nand2_1
X_6478_ net1229 VPWR _0994_ VGND net1217 net1395 sg13g2_o21ai_1
X_5429_ VPWR _2847_ net509 VGND sg13g2_inv_1
XFILLER_0_803 VPWR VGND sg13g2_decap_8
XFILLER_28_564 VPWR VGND sg13g2_decap_8
XFILLER_43_512 VPWR VGND sg13g2_fill_1
XFILLER_12_954 VPWR VGND sg13g2_decap_8
XFILLER_30_239 VPWR VGND sg13g2_fill_2
XFILLER_8_947 VPWR VGND sg13g2_decap_8
XFILLER_48_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_641 VPWR VGND sg13g2_fill_1
Xfanout1431 net1434 net1431 VPWR VGND sg13g2_buf_1
Xfanout1420 ui_in[5] net1420 VPWR VGND sg13g2_buf_8
Xfanout1475 net1476 net1475 VPWR VGND sg13g2_buf_8
Xfanout1453 net1457 net1453 VPWR VGND sg13g2_buf_1
Xfanout1464 net1465 net1464 VPWR VGND sg13g2_buf_8
Xfanout1442 ui_in[3] net1442 VPWR VGND sg13g2_buf_8
X_6548__297 VPWR VGND net297 sg13g2_tiehi
Xfanout1486 net1487 net1486 VPWR VGND sg13g2_buf_8
XFILLER_0_43 VPWR VGND sg13g2_fill_1
XFILLER_0_65 VPWR VGND sg13g2_decap_8
XFILLER_22_718 VPWR VGND sg13g2_fill_2
X_4800_ s0.data_out\[4\]\[3\] s0.data_out\[3\]\[3\] net1057 _2275_ VPWR VGND sg13g2_mux2_1
X_5780_ VGND VPWR net1305 _0362_ _0365_ _0364_ sg13g2_a21oi_1
X_6694__139 VPWR VGND net139 sg13g2_tiehi
X_4731_ VPWR _0228_ _2216_ VGND sg13g2_inv_1
X_4662_ s0.data_out\[5\]\[2\] s0.data_out\[4\]\[2\] net1068 _2149_ VPWR VGND sg13g2_mux2_1
X_6401_ s0.data_out\[16\]\[6\] s0.data_out\[15\]\[6\] net1233 _0926_ VPWR VGND sg13g2_mux2_1
X_3613_ _1208_ VPWR _1209_ VGND net1017 _1207_ sg13g2_o21ai_1
XFILLER_31_1020 VPWR VGND sg13g2_decap_8
X_4593_ _2055_ _2073_ _2088_ _2091_ _2092_ VPWR VGND sg13g2_or4_1
X_6332_ net1366 _0786_ _0866_ VPWR VGND sg13g2_nor2_1
X_3544_ _1146_ _1145_ net1441 _1122_ net1445 VPWR VGND sg13g2_a22oi_1
X_3475_ net1018 _2823_ _1086_ VPWR VGND sg13g2_nor2_1
X_6263_ s0.data_out\[16\]\[0\] s0.data_out\[17\]\[0\] net1260 _0800_ VPWR VGND sg13g2_mux2_1
X_5214_ VPWR VGND _2627_ _2652_ _2650_ _2611_ _2653_ _2649_ sg13g2_a221oi_1
XFILLER_9_1010 VPWR VGND sg13g2_decap_8
X_6194_ _0721_ _0736_ _0738_ _0743_ VPWR VGND sg13g2_nor3_1
X_5145_ s0.data_out\[1\]\[2\] s0.data_out\[0\]\[2\] net1024 _2584_ VPWR VGND sg13g2_mux2_1
XFILLER_29_328 VPWR VGND sg13g2_fill_2
X_5076_ _2527_ _2751_ _2526_ VPWR VGND sg13g2_nand2_1
X_4027_ VGND VPWR net1136 _1571_ _1574_ _1573_ sg13g2_a21oi_1
X_5978_ net1288 VPWR _0545_ VGND _0514_ _0544_ sg13g2_o21ai_1
XFILLER_25_589 VPWR VGND sg13g2_decap_8
X_4929_ VGND VPWR _2274_ _2391_ _2392_ net1048 sg13g2_a21oi_1
XFILLER_21_773 VPWR VGND sg13g2_decap_4
XFILLER_5_906 VPWR VGND sg13g2_decap_8
XFILLER_20_261 VPWR VGND sg13g2_fill_1
X_6499__54 VPWR VGND net54 sg13g2_tiehi
XFILLER_0_600 VPWR VGND sg13g2_decap_8
XFILLER_48_604 VPWR VGND sg13g2_decap_8
XFILLER_0_677 VPWR VGND sg13g2_decap_8
XFILLER_48_648 VPWR VGND sg13g2_decap_8
XFILLER_29_862 VPWR VGND sg13g2_fill_2
XFILLER_28_361 VPWR VGND sg13g2_fill_1
XFILLER_7_232 VPWR VGND sg13g2_fill_1
XFILLER_8_788 VPWR VGND sg13g2_fill_2
XFILLER_8_766 VPWR VGND sg13g2_fill_1
XFILLER_7_287 VPWR VGND sg13g2_fill_1
X_6554__290 VPWR VGND net290 sg13g2_tiehi
XFILLER_4_950 VPWR VGND sg13g2_decap_8
Xfanout1250 net1251 net1250 VPWR VGND sg13g2_buf_8
XFILLER_22_4 VPWR VGND sg13g2_fill_2
Xfanout1261 net1264 net1261 VPWR VGND sg13g2_buf_8
Xfanout1272 s0.valid_out\[18\][0] net1272 VPWR VGND sg13g2_buf_8
Xfanout1283 net1285 net1283 VPWR VGND sg13g2_buf_8
XFILLER_22_1008 VPWR VGND sg13g2_decap_8
Xfanout1294 net1295 net1294 VPWR VGND sg13g2_buf_1
XFILLER_19_350 VPWR VGND sg13g2_fill_2
XFILLER_47_692 VPWR VGND sg13g2_decap_8
X_5901_ _0474_ _0473_ net1293 VPWR VGND sg13g2_nand2b_1
X_6561__283 VPWR VGND net283 sg13g2_tiehi
XFILLER_35_898 VPWR VGND sg13g2_fill_2
X_5832_ net1291 s0.data_out\[20\]\[0\] _0416_ VPWR VGND sg13g2_and2_1
XFILLER_34_353 VPWR VGND sg13g2_fill_2
X_5763_ _0348_ net1305 _0347_ VPWR VGND sg13g2_nand2b_1
X_4714_ _2201_ _2200_ net1077 VPWR VGND sg13g2_nand2b_1
X_5694_ VGND VPWR _3082_ _3084_ _3088_ net1416 sg13g2_a21oi_1
X_4645_ net1363 _2126_ _2127_ _0225_ VPWR VGND sg13g2_nor3_1
XFILLER_30_29 VPWR VGND sg13g2_fill_1
X_4576_ s0.data_out\[6\]\[4\] s0.data_out\[5\]\[4\] net1081 _2075_ VPWR VGND sg13g2_mux2_1
X_6315_ _0840_ VPWR _0852_ VGND net1439 _0810_ sg13g2_o21ai_1
X_3527_ VGND VPWR _1013_ _1128_ _1129_ net1214 sg13g2_a21oi_1
X_3458_ VGND VPWR _1067_ _1069_ _1072_ net1432 sg13g2_a21oi_1
X_6246_ net1238 net1165 _0783_ VPWR VGND sg13g2_nor2b_1
X_6496__57 VPWR VGND net57 sg13g2_tiehi
X_3389_ net328 net1485 _0099_ VPWR VGND sg13g2_and2_1
X_6177_ _0726_ s0.data_out\[17\]\[4\] net1271 VPWR VGND sg13g2_nand2b_1
X_5128_ net1032 s0.data_out\[1\]\[7\] _2571_ VPWR VGND sg13g2_and2_1
XFILLER_29_136 VPWR VGND sg13g2_decap_4
XFILLER_45_629 VPWR VGND sg13g2_fill_1
X_5059_ VGND VPWR _2395_ _2509_ _2510_ net1039 sg13g2_a21oi_1
XFILLER_41_824 VPWR VGND sg13g2_fill_2
XFILLER_40_301 VPWR VGND sg13g2_fill_1
XFILLER_38_1026 VPWR VGND sg13g2_fill_2
XFILLER_9_519 VPWR VGND sg13g2_decap_4
XFILLER_21_581 VPWR VGND sg13g2_fill_2
XFILLER_5_714 VPWR VGND sg13g2_decap_8
XFILLER_5_736 VPWR VGND sg13g2_fill_1
XFILLER_45_1019 VPWR VGND sg13g2_decap_8
XFILLER_1_975 VPWR VGND sg13g2_decap_8
XFILLER_49_968 VPWR VGND sg13g2_decap_8
XFILLER_0_474 VPWR VGND sg13g2_decap_8
Xhold60 _0005_ VPWR VGND net380 sg13g2_dlygate4sd3_1
Xhold71 s0.shift_out\[12\][0] VPWR VGND net391 sg13g2_dlygate4sd3_1
Xhold82 s0.data_out\[0\]\[3\] VPWR VGND net402 sg13g2_dlygate4sd3_1
Xhold93 _0007_ VPWR VGND net413 sg13g2_dlygate4sd3_1
XFILLER_45_70 VPWR VGND sg13g2_fill_1
XFILLER_44_695 VPWR VGND sg13g2_fill_2
XFILLER_16_386 VPWR VGND sg13g2_decap_4
X_4430_ VPWR VGND net1442 _1933_ _1940_ net1447 _1941_ _1916_ sg13g2_a221oi_1
X_6100_ _0058_ net437 _0654_ _2792_ net1353 VPWR VGND sg13g2_a22oi_1
X_4361_ _0193_ _1880_ _1881_ _2853_ net1374 VPWR VGND sg13g2_a22oi_1
X_4292_ _1815_ net1106 s0.data_out\[7\]\[0\] VPWR VGND sg13g2_nand2_1
X_6031_ _0592_ _0591_ net1437 _0568_ net1444 VPWR VGND sg13g2_a22oi_1
Xfanout1091 net446 net1091 VPWR VGND sg13g2_buf_2
XFILLER_13_0 VPWR VGND sg13g2_fill_2
Xfanout1080 net1084 net1080 VPWR VGND sg13g2_buf_8
XFILLER_39_489 VPWR VGND sg13g2_decap_8
XFILLER_35_695 VPWR VGND sg13g2_fill_1
X_5815_ net1289 net1151 _0400_ VPWR VGND sg13g2_nor2b_1
XFILLER_41_17 VPWR VGND sg13g2_fill_1
X_5746_ net1008 VPWR _0334_ VGND net649 net1308 sg13g2_o21ai_1
X_5677_ _3071_ net1309 s0.data_out\[21\]\[4\] VPWR VGND sg13g2_nand2_1
X_4628_ net1088 VPWR _2120_ VGND _2065_ _2119_ sg13g2_o21ai_1
X_4559_ net1078 net1144 _2058_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_728 VPWR VGND sg13g2_decap_8
X_6229_ net1002 _2803_ _0770_ VPWR VGND sg13g2_nor2_1
X_6609__231 VPWR VGND net231 sg13g2_tiehi
XFILLER_17_117 VPWR VGND sg13g2_fill_1
XFILLER_45_437 VPWR VGND sg13g2_fill_2
XFILLER_14_802 VPWR VGND sg13g2_decap_8
XFILLER_25_183 VPWR VGND sg13g2_fill_2
XFILLER_9_316 VPWR VGND sg13g2_decap_4
XFILLER_15_51 VPWR VGND sg13g2_fill_1
XFILLER_13_389 VPWR VGND sg13g2_fill_1
XFILLER_5_522 VPWR VGND sg13g2_decap_8
XFILLER_5_588 VPWR VGND sg13g2_fill_2
Xoutput4 net4 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_772 VPWR VGND sg13g2_decap_8
XFILLER_49_765 VPWR VGND sg13g2_decap_8
XFILLER_0_293 VPWR VGND sg13g2_decap_4
XFILLER_17_640 VPWR VGND sg13g2_fill_2
X_3930_ _1494_ net1138 _1495_ _1496_ VPWR VGND sg13g2_a21o_1
X_3861_ VPWR _0140_ _1434_ VGND sg13g2_inv_1
X_5600_ net1311 s0.data_out\[22\]\[5\] _3000_ VPWR VGND sg13g2_and2_1
X_6580_ net262 VGND VPWR net480 s0.data_out\[16\]\[1\] clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_20_838 VPWR VGND sg13g2_fill_1
X_3792_ _1371_ net1440 _1368_ VPWR VGND sg13g2_nand2_1
XFILLER_31_164 VPWR VGND sg13g2_decap_4
XFILLER_9_872 VPWR VGND sg13g2_decap_4
X_5531_ VGND VPWR net1326 _2936_ _2937_ _2932_ sg13g2_a21oi_1
XFILLER_8_360 VPWR VGND sg13g2_decap_8
X_5462_ VPWR _2880_ net512 VGND sg13g2_inv_1
X_5393_ VPWR _2811_ net482 VGND sg13g2_inv_1
X_4413_ VGND VPWR net1096 _1921_ _1924_ _1923_ sg13g2_a21oi_1
X_4344_ _1867_ net1431 _1866_ VPWR VGND sg13g2_nand2_1
XFILLER_28_1025 VPWR VGND sg13g2_decap_4
X_4275_ net1481 _1794_ _0189_ VPWR VGND sg13g2_and2_1
X_6014_ VGND VPWR _0462_ _0574_ _0575_ net1279 sg13g2_a21oi_1
XFILLER_27_448 VPWR VGND sg13g2_fill_1
XFILLER_36_993 VPWR VGND sg13g2_decap_8
XFILLER_22_153 VPWR VGND sg13g2_fill_1
X_6778_ net156 VGND VPWR _0288_ s0.data_out\[0\]\[0\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_5729_ VPWR _0022_ net565 VGND sg13g2_inv_1
Xhold360 s0.data_out\[9\]\[5\] VPWR VGND net680 sg13g2_dlygate4sd3_1
Xhold371 _0056_ VPWR VGND net691 sg13g2_dlygate4sd3_1
Xhold382 s0.data_new_delayed\[1\] VPWR VGND net702 sg13g2_dlygate4sd3_1
XFILLER_18_426 VPWR VGND sg13g2_fill_2
XFILLER_19_927 VPWR VGND sg13g2_fill_1
XFILLER_46_757 VPWR VGND sg13g2_decap_8
XFILLER_18_437 VPWR VGND sg13g2_fill_1
XFILLER_27_971 VPWR VGND sg13g2_decap_8
XFILLER_13_120 VPWR VGND sg13g2_fill_2
XFILLER_42_985 VPWR VGND sg13g2_decap_8
XFILLER_13_153 VPWR VGND sg13g2_decap_4
XFILLER_42_71 VPWR VGND sg13g2_fill_1
XFILLER_6_886 VPWR VGND sg13g2_decap_8
XFILLER_3_10 VPWR VGND sg13g2_fill_1
X_4060_ net1128 net1144 _1607_ VPWR VGND sg13g2_nor2b_1
XFILLER_3_76 VPWR VGND sg13g2_fill_2
XFILLER_49_562 VPWR VGND sg13g2_decap_8
XFILLER_3_1027 VPWR VGND sg13g2_fill_2
XFILLER_36_245 VPWR VGND sg13g2_decap_8
X_4962_ _2425_ s0.data_out\[2\]\[4\] net1056 VPWR VGND sg13g2_nand2b_1
X_6701_ net132 VGND VPWR _0211_ s0.data_out\[7\]\[7\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_4893_ VGND VPWR _2359_ _2358_ _2356_ sg13g2_or2_1
XFILLER_32_451 VPWR VGND sg13g2_fill_2
X_3913_ net1136 net1161 _1479_ VPWR VGND sg13g2_nor2b_1
X_6632_ net206 VGND VPWR net620 s0.data_out\[12\]\[6\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_3844_ net1178 s0.data_out\[11\]\[1\] _1421_ VPWR VGND sg13g2_and2_1
X_6563_ net281 VGND VPWR _0073_ s0.was_valid_out\[17\][0] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3775_ net1180 net1164 _1354_ VPWR VGND sg13g2_nor2b_1
X_6494_ net59 VGND VPWR _0004_ s0.shift_out\[23\][0] clknet_leaf_1_clk sg13g2_dfrbpq_2
X_5514_ _2920_ net1449 _2919_ VPWR VGND sg13g2_nand2_1
X_5445_ VPWR _2863_ net501 VGND sg13g2_inv_1
X_5376_ VPWR _2794_ net690 VGND sg13g2_inv_1
X_4327_ VPWR _1850_ _1849_ VGND sg13g2_inv_1
X_4258_ net1126 VPWR _1786_ VGND _1721_ _1785_ sg13g2_o21ai_1
XFILLER_41_1022 VPWR VGND sg13g2_decap_8
XFILLER_28_724 VPWR VGND sg13g2_decap_8
X_4189_ VGND VPWR _1612_ _1723_ _1724_ net1126 sg13g2_a21oi_1
X_6606__234 VPWR VGND net234 sg13g2_tiehi
XFILLER_16_919 VPWR VGND sg13g2_fill_2
XFILLER_24_963 VPWR VGND sg13g2_decap_8
XFILLER_6_127 VPWR VGND sg13g2_fill_2
XFILLER_12_74 VPWR VGND sg13g2_fill_1
XFILLER_3_845 VPWR VGND sg13g2_decap_8
Xhold190 _0186_ VPWR VGND net510 sg13g2_dlygate4sd3_1
XFILLER_15_985 VPWR VGND sg13g2_decap_8
XFILLER_30_933 VPWR VGND sg13g2_fill_2
XFILLER_41_292 VPWR VGND sg13g2_decap_4
X_3560_ _1162_ _1161_ net1413 _1154_ net1404 VPWR VGND sg13g2_a22oi_1
X_3491_ _0106_ _1097_ _1098_ _2815_ net1380 VPWR VGND sg13g2_a22oi_1
XFILLER_5_160 VPWR VGND sg13g2_fill_1
X_5230_ VGND VPWR net1021 net402 _2665_ _2606_ sg13g2_a21oi_1
XFILLER_38_2 VPWR VGND sg13g2_fill_1
X_5161_ _2600_ net1029 _2599_ VPWR VGND sg13g2_nand2b_1
X_5092_ _2466_ VPWR _2543_ VGND _2518_ _2520_ sg13g2_o21ai_1
X_4112_ VGND VPWR net1124 net465 _1656_ _1585_ sg13g2_a21oi_1
X_4043_ VGND VPWR _1590_ _1589_ net1335 sg13g2_or2_1
X_5994_ net1261 _0553_ _0558_ VPWR VGND sg13g2_nor2_1
X_4945_ VGND VPWR net1052 _2405_ _2408_ _2407_ sg13g2_a21oi_1
X_4876_ VGND VPWR net996 _2316_ _2345_ net1361 sg13g2_a21oi_1
XFILLER_21_999 VPWR VGND sg13g2_decap_8
X_6615_ net224 VGND VPWR _0125_ s0.data_out\[13\]\[0\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3827_ _1403_ _1405_ net1423 _1406_ VPWR VGND sg13g2_nand3_1
X_6546_ net299 VGND VPWR net691 s0.data_out\[19\]\[3\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3758_ net1485 _1332_ _0134_ VPWR VGND sg13g2_and2_1
XFILLER_3_108 VPWR VGND sg13g2_fill_2
X_6477_ _0096_ _0992_ _0993_ _2808_ net1368 VPWR VGND sg13g2_a22oi_1
X_3689_ _1279_ net1207 _1278_ VPWR VGND sg13g2_nand2b_1
X_5428_ VPWR _2846_ net505 VGND sg13g2_inv_1
X_5359_ VPWR _2777_ net603 VGND sg13g2_inv_1
XFILLER_0_859 VPWR VGND sg13g2_decap_8
XFILLER_16_738 VPWR VGND sg13g2_fill_2
XFILLER_28_598 VPWR VGND sg13g2_decap_4
XFILLER_15_248 VPWR VGND sg13g2_decap_8
XFILLER_31_708 VPWR VGND sg13g2_decap_4
XFILLER_8_926 VPWR VGND sg13g2_decap_8
XFILLER_23_40 VPWR VGND sg13g2_decap_8
XFILLER_7_469 VPWR VGND sg13g2_fill_1
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
X_6687__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_2_130 VPWR VGND sg13g2_fill_2
XFILLER_2_174 VPWR VGND sg13g2_fill_2
XFILLER_39_808 VPWR VGND sg13g2_fill_2
Xfanout1421 net1425 net1421 VPWR VGND sg13g2_buf_8
Xfanout1410 ui_in[6] net1410 VPWR VGND sg13g2_buf_8
Xfanout1432 net1434 net1432 VPWR VGND sg13g2_buf_8
Xfanout1443 net1448 net1443 VPWR VGND sg13g2_buf_8
Xfanout1454 net1456 net1454 VPWR VGND sg13g2_buf_8
Xfanout1465 net1469 net1465 VPWR VGND sg13g2_buf_8
XFILLER_0_11 VPWR VGND sg13g2_decap_8
Xfanout1476 net1493 net1476 VPWR VGND sg13g2_buf_8
Xfanout1487 net1493 net1487 VPWR VGND sg13g2_buf_8
XFILLER_47_885 VPWR VGND sg13g2_decap_8
XFILLER_0_55 VPWR VGND sg13g2_fill_1
XFILLER_0_99 VPWR VGND sg13g2_decap_4
XFILLER_0_88 VPWR VGND sg13g2_decap_8
X_4730_ _2215_ VPWR _2216_ VGND net1474 net571 sg13g2_o21ai_1
XFILLER_9_75 VPWR VGND sg13g2_fill_1
X_4661_ _2148_ net1067 net676 VPWR VGND sg13g2_nand2_1
X_6400_ _0925_ net1234 s0.data_out\[15\]\[6\] VPWR VGND sg13g2_nand2_1
X_3612_ VGND VPWR net1017 _1171_ _1208_ net1381 sg13g2_a21oi_1
X_4592_ VGND VPWR _2091_ _2090_ _2089_ sg13g2_or2_1
X_6331_ net1254 VPWR _0865_ VGND _0783_ _0864_ sg13g2_o21ai_1
XFILLER_7_981 VPWR VGND sg13g2_decap_8
X_3543_ VGND VPWR net1216 _1142_ _1145_ _1144_ sg13g2_a21oi_1
XFILLER_43_0 VPWR VGND sg13g2_fill_1
X_3474_ _0102_ _1084_ _1085_ _2818_ net1369 VPWR VGND sg13g2_a22oi_1
X_6262_ _0799_ net1255 _0798_ VPWR VGND sg13g2_nand2b_1
X_5213_ _2652_ _2651_ _2577_ VPWR VGND sg13g2_nand2b_1
X_6193_ _0703_ _0721_ _0741_ _0742_ VPWR VGND sg13g2_or3_1
X_5144_ s0.data_out\[0\]\[2\] s0.data_out\[1\]\[2\] net1033 _2583_ VPWR VGND sg13g2_mux2_1
X_5075_ s0.data_out\[1\]\[4\] s0.data_out\[2\]\[4\] net1043 _2526_ VPWR VGND sg13g2_mux2_1
X_4026_ VGND VPWR _1462_ _1572_ _1573_ net1135 sg13g2_a21oi_1
XFILLER_37_384 VPWR VGND sg13g2_fill_1
XFILLER_25_502 VPWR VGND sg13g2_fill_2
XFILLER_44_39 VPWR VGND sg13g2_fill_2
X_6603__237 VPWR VGND net237 sg13g2_tiehi
XFILLER_25_535 VPWR VGND sg13g2_decap_4
X_5977_ net1003 _2792_ _0544_ VPWR VGND sg13g2_nor2_1
X_4928_ _2391_ _2748_ net463 VPWR VGND sg13g2_nand2_1
X_4859_ net1060 VPWR _2332_ VGND _2261_ _2331_ sg13g2_o21ai_1
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
X_6529_ net317 VGND VPWR _0039_ s0.genblk1\[1\].modules.bubble clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
XFILLER_0_656 VPWR VGND sg13g2_decap_8
XFILLER_48_627 VPWR VGND sg13g2_decap_8
XFILLER_18_73 VPWR VGND sg13g2_fill_2
XFILLER_16_546 VPWR VGND sg13g2_fill_2
XFILLER_16_557 VPWR VGND sg13g2_decap_8
XFILLER_43_376 VPWR VGND sg13g2_fill_1
X_6693__140 VPWR VGND net140 sg13g2_tiehi
XFILLER_15_1027 VPWR VGND sg13g2_fill_2
XFILLER_11_251 VPWR VGND sg13g2_fill_2
XFILLER_8_778 VPWR VGND sg13g2_fill_1
XFILLER_7_266 VPWR VGND sg13g2_fill_1
XFILLER_7_255 VPWR VGND sg13g2_decap_8
Xfanout1240 net1244 net1240 VPWR VGND sg13g2_buf_8
Xfanout1273 net1275 net1273 VPWR VGND sg13g2_buf_8
Xfanout1262 net1263 net1262 VPWR VGND sg13g2_buf_8
Xfanout1251 net498 net1251 VPWR VGND sg13g2_buf_8
Xfanout1295 s0.shift_out\[20\][0] net1295 VPWR VGND sg13g2_buf_1
Xfanout1284 net1285 net1284 VPWR VGND sg13g2_buf_2
XFILLER_47_671 VPWR VGND sg13g2_decap_8
X_5900_ s0.data_out\[19\]\[0\] s0.data_out\[20\]\[0\] net1298 _0473_ VPWR VGND sg13g2_mux2_1
X_5831_ VGND VPWR _0410_ _0414_ _0028_ _0415_ sg13g2_a21oi_1
X_5762_ VGND VPWR net1290 _0346_ _0347_ _0345_ sg13g2_a21oi_1
XFILLER_22_527 VPWR VGND sg13g2_fill_1
X_4713_ s0.data_out\[4\]\[5\] s0.data_out\[5\]\[5\] net1082 _2200_ VPWR VGND sg13g2_mux2_1
X_5693_ VGND VPWR _3074_ _3076_ _3087_ net1426 sg13g2_a21oi_1
XFILLER_30_571 VPWR VGND sg13g2_fill_2
X_4644_ VGND VPWR _2730_ _2128_ _0224_ _2133_ sg13g2_a21oi_1
X_4575_ net1075 net1158 _2074_ VPWR VGND sg13g2_nor2b_1
X_6314_ _0851_ _0848_ _0849_ VPWR VGND sg13g2_nand2_1
X_3526_ _1128_ net481 net1219 VPWR VGND sg13g2_nand2b_1
X_6245_ s0.data_out\[17\]\[2\] s0.data_out\[16\]\[2\] net1246 _0782_ VPWR VGND sg13g2_mux2_1
XFILLER_39_39 VPWR VGND sg13g2_fill_2
X_3457_ _1071_ net1423 _1061_ VPWR VGND sg13g2_nand2_1
X_6176_ _0723_ net1252 _0724_ _0725_ VPWR VGND sg13g2_a21o_1
X_5127_ _0270_ _2569_ _2570_ _2881_ net1349 VPWR VGND sg13g2_a22oi_1
XFILLER_29_115 VPWR VGND sg13g2_decap_8
X_5058_ _2509_ s0.data_out\[1\]\[7\] net1045 VPWR VGND sg13g2_nand2b_1
X_4009_ net1491 _1559_ _0158_ VPWR VGND sg13g2_and2_1
XFILLER_38_1005 VPWR VGND sg13g2_decap_8
XFILLER_13_527 VPWR VGND sg13g2_decap_4
XFILLER_25_387 VPWR VGND sg13g2_decap_4
XFILLER_40_379 VPWR VGND sg13g2_fill_1
XFILLER_0_431 VPWR VGND sg13g2_decap_8
XFILLER_1_954 VPWR VGND sg13g2_decap_8
XFILLER_0_442 VPWR VGND sg13g2_fill_1
XFILLER_49_947 VPWR VGND sg13g2_decap_8
Xhold50 s0.was_valid_out\[16\][0] VPWR VGND net370 sg13g2_dlygate4sd3_1
XFILLER_36_619 VPWR VGND sg13g2_fill_1
XFILLER_36_608 VPWR VGND sg13g2_decap_8
Xhold72 s0.was_valid_out\[22\][0] VPWR VGND net392 sg13g2_dlygate4sd3_1
Xhold61 s0.data_out\[23\]\[1\] VPWR VGND net381 sg13g2_dlygate4sd3_1
XFILLER_21_1020 VPWR VGND sg13g2_decap_8
XFILLER_29_72 VPWR VGND sg13g2_fill_1
Xhold83 _0291_ VPWR VGND net403 sg13g2_dlygate4sd3_1
Xhold94 s0.data_out\[12\]\[4\] VPWR VGND net414 sg13g2_dlygate4sd3_1
XFILLER_29_660 VPWR VGND sg13g2_decap_8
XFILLER_17_833 VPWR VGND sg13g2_fill_2
XFILLER_28_170 VPWR VGND sg13g2_decap_8
XFILLER_28_181 VPWR VGND sg13g2_fill_2
XFILLER_17_899 VPWR VGND sg13g2_fill_2
XFILLER_43_162 VPWR VGND sg13g2_fill_1
XFILLER_31_346 VPWR VGND sg13g2_fill_1
XFILLER_31_368 VPWR VGND sg13g2_decap_8
XFILLER_12_582 VPWR VGND sg13g2_fill_1
XFILLER_8_553 VPWR VGND sg13g2_fill_1
X_4360_ net1374 _1813_ _1881_ VPWR VGND sg13g2_nor2_1
X_4291_ VGND VPWR net1110 _1811_ _1814_ _1813_ sg13g2_a21oi_1
XFILLER_3_291 VPWR VGND sg13g2_fill_1
X_6030_ VGND VPWR net1279 _0588_ _0591_ _0590_ sg13g2_a21oi_1
Xfanout1070 net1071 net1070 VPWR VGND sg13g2_buf_2
XFILLER_39_468 VPWR VGND sg13g2_decap_8
Xfanout1081 net1084 net1081 VPWR VGND sg13g2_buf_8
Xfanout1092 s0.valid_out\[6\][0] net1092 VPWR VGND sg13g2_buf_8
XFILLER_48_991 VPWR VGND sg13g2_decap_8
XFILLER_27_619 VPWR VGND sg13g2_fill_2
X_5814_ s0.data_out\[21\]\[5\] s0.data_out\[20\]\[5\] net1296 _0399_ VPWR VGND sg13g2_mux2_1
X_5745_ VGND VPWR _0333_ _0326_ net1286 sg13g2_or2_1
XFILLER_31_880 VPWR VGND sg13g2_fill_2
X_5676_ net1304 net1156 _3070_ VPWR VGND sg13g2_nor2b_1
X_4627_ net1079 net449 _2119_ VPWR VGND sg13g2_and2_1
X_4558_ s0.data_out\[6\]\[7\] s0.data_out\[5\]\[7\] net1083 _2057_ VPWR VGND sg13g2_mux2_1
XFILLER_2_707 VPWR VGND sg13g2_decap_8
X_4489_ net1097 VPWR _1996_ VGND _1936_ _1995_ sg13g2_o21ai_1
XFILLER_1_239 VPWR VGND sg13g2_decap_8
X_3509_ VGND VPWR _1108_ _1111_ _1114_ _1113_ sg13g2_a21oi_1
X_6228_ VPWR _0071_ net535 VGND sg13g2_inv_1
X_6159_ _0708_ s0.data_out\[17\]\[7\] net1269 VPWR VGND sg13g2_nand2b_1
X_6492__61 VPWR VGND net61 sg13g2_tiehi
XFILLER_18_608 VPWR VGND sg13g2_fill_2
XFILLER_46_939 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_37_clk clknet_3_1__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_25_140 VPWR VGND sg13g2_decap_8
XFILLER_25_151 VPWR VGND sg13g2_fill_1
XFILLER_25_162 VPWR VGND sg13g2_decap_8
XFILLER_25_173 VPWR VGND sg13g2_fill_1
XFILLER_40_143 VPWR VGND sg13g2_fill_1
XFILLER_9_306 VPWR VGND sg13g2_decap_4
Xoutput5 net5 uo_out[3] VPWR VGND sg13g2_buf_1
X_6551__294 VPWR VGND net294 sg13g2_tiehi
XFILLER_1_751 VPWR VGND sg13g2_decap_8
XFILLER_49_744 VPWR VGND sg13g2_decap_8
XFILLER_37_917 VPWR VGND sg13g2_fill_1
XFILLER_36_416 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_28_clk clknet_3_5__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_44_482 VPWR VGND sg13g2_decap_4
X_3860_ _1433_ VPWR _1434_ VGND net1486 net414 sg13g2_o21ai_1
X_3791_ _1351_ _1360_ _1361_ _1369_ _1370_ VPWR VGND sg13g2_nor4_1
X_5530_ _2934_ net1315 _2935_ _2936_ VPWR VGND sg13g2_a21o_1
X_5461_ VPWR _2879_ net400 VGND sg13g2_inv_1
X_4412_ VGND VPWR _1808_ _1922_ _1923_ net1096 sg13g2_a21oi_1
X_5392_ _2810_ net525 VPWR VGND sg13g2_inv_2
X_4343_ VGND VPWR net1114 _1863_ _1866_ _1865_ sg13g2_a21oi_1
XFILLER_28_1004 VPWR VGND sg13g2_decap_8
X_4274_ VGND VPWR _2732_ _1794_ _0188_ _1799_ sg13g2_a21oi_1
X_6013_ _0574_ net418 net1283 VPWR VGND sg13g2_nand2b_1
XFILLER_39_243 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_19_clk clknet_3_7__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_36_972 VPWR VGND sg13g2_decap_8
X_6777_ net169 VGND VPWR _0287_ s0.shift_out\[0\][0] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_5728_ _0318_ VPWR _0319_ VGND net1463 net564 sg13g2_o21ai_1
X_3989_ VPWR _0154_ _1548_ VGND sg13g2_inv_1
X_5659_ s0.data_out\[22\]\[7\] s0.data_out\[21\]\[7\] net1307 _3053_ VPWR VGND sg13g2_mux2_1
Xhold361 s0.data_out\[4\]\[5\] VPWR VGND net681 sg13g2_dlygate4sd3_1
Xhold350 s0.data_out\[8\]\[4\] VPWR VGND net670 sg13g2_dlygate4sd3_1
XFILLER_2_526 VPWR VGND sg13g2_decap_8
Xhold383 s0.shift_out\[16\][0] VPWR VGND net703 sg13g2_dlygate4sd3_1
Xhold372 s0.data_out\[6\]\[0\] VPWR VGND net692 sg13g2_dlygate4sd3_1
XFILLER_45_257 VPWR VGND sg13g2_decap_4
XFILLER_33_419 VPWR VGND sg13g2_fill_2
XFILLER_26_73 VPWR VGND sg13g2_fill_1
XFILLER_42_964 VPWR VGND sg13g2_decap_8
XFILLER_14_633 VPWR VGND sg13g2_fill_1
XFILLER_41_474 VPWR VGND sg13g2_decap_4
XFILLER_9_125 VPWR VGND sg13g2_fill_1
XFILLER_14_677 VPWR VGND sg13g2_fill_2
XFILLER_42_83 VPWR VGND sg13g2_decap_8
XFILLER_5_342 VPWR VGND sg13g2_fill_2
XFILLER_49_541 VPWR VGND sg13g2_decap_8
XFILLER_3_1006 VPWR VGND sg13g2_decap_8
XFILLER_36_213 VPWR VGND sg13g2_decap_4
XFILLER_18_994 VPWR VGND sg13g2_decap_8
X_4961_ _2422_ net1037 _2423_ _2424_ VPWR VGND sg13g2_a21o_1
X_6700_ net133 VGND VPWR _0210_ s0.data_out\[7\]\[6\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_4892_ net356 net1045 _2358_ VPWR VGND sg13g2_nor2_1
XFILLER_17_493 VPWR VGND sg13g2_decap_8
XFILLER_32_441 VPWR VGND sg13g2_decap_4
X_3912_ s0.data_out\[11\]\[3\] s0.data_out\[10\]\[3\] net1177 _1478_ VPWR VGND sg13g2_mux2_1
XFILLER_20_603 VPWR VGND sg13g2_decap_8
X_3843_ VPWR _0136_ _1420_ VGND sg13g2_inv_1
X_6631_ net207 VGND VPWR _0141_ s0.data_out\[12\]\[5\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_33_986 VPWR VGND sg13g2_decap_8
X_6562_ net282 VGND VPWR net500 s0.data_out\[18\]\[7\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3774_ s0.data_out\[12\]\[2\] s0.data_out\[11\]\[2\] net1187 _1353_ VPWR VGND sg13g2_mux2_1
X_6493_ net60 VGND VPWR _0003_ s0.genblk1\[22\].modules.bubble clknet_leaf_0_clk sg13g2_dfrbpq_1
X_5513_ VGND VPWR net1325 _2918_ _2919_ _2914_ sg13g2_a21oi_1
Xclkbuf_leaf_8_clk clknet_3_2__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_5444_ VPWR _2862_ net389 VGND sg13g2_inv_1
X_5375_ VPWR _2793_ net486 VGND sg13g2_inv_1
X_4326_ VGND VPWR _1849_ _1846_ net1403 sg13g2_or2_1
X_4257_ net1117 s0.data_out\[8\]\[6\] _1785_ VPWR VGND sg13g2_and2_1
XFILLER_41_1001 VPWR VGND sg13g2_decap_8
X_4188_ _1723_ s0.data_out\[8\]\[6\] net1132 VPWR VGND sg13g2_nand2b_1
XFILLER_27_235 VPWR VGND sg13g2_fill_1
XFILLER_3_824 VPWR VGND sg13g2_decap_8
Xhold180 _0072_ VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold191 s0.data_out\[17\]\[2\] VPWR VGND net511 sg13g2_dlygate4sd3_1
XFILLER_46_533 VPWR VGND sg13g2_decap_4
XFILLER_18_202 VPWR VGND sg13g2_decap_8
XFILLER_19_758 VPWR VGND sg13g2_fill_2
XFILLER_46_566 VPWR VGND sg13g2_fill_2
XFILLER_46_599 VPWR VGND sg13g2_fill_1
XFILLER_15_964 VPWR VGND sg13g2_decap_8
XFILLER_30_989 VPWR VGND sg13g2_decap_8
XFILLER_10_680 VPWR VGND sg13g2_decap_4
X_3490_ net1380 _1060_ _1098_ VPWR VGND sg13g2_nor2_1
X_5160_ VGND VPWR net1020 _2597_ _2599_ _2598_ sg13g2_a21oi_1
X_5091_ _2521_ _2541_ _2542_ VPWR VGND sg13g2_nor2b_1
X_4111_ _0169_ _1654_ _1655_ _2839_ net1385 VPWR VGND sg13g2_a22oi_1
XFILLER_49_360 VPWR VGND sg13g2_decap_8
X_4042_ _1588_ VPWR _1589_ VGND net1014 _1586_ sg13g2_o21ai_1
XFILLER_49_382 VPWR VGND sg13g2_fill_2
XFILLER_37_522 VPWR VGND sg13g2_decap_8
X_5993_ _0555_ VPWR _0557_ VGND s0.was_valid_out\[18\][0] net1269 sg13g2_o21ai_1
XFILLER_24_205 VPWR VGND sg13g2_fill_2
X_4944_ VGND VPWR _2290_ _2406_ _2407_ net1052 sg13g2_a21oi_1
XFILLER_17_290 VPWR VGND sg13g2_fill_2
XFILLER_21_901 VPWR VGND sg13g2_fill_2
X_4875_ VGND VPWR net1053 net601 _2344_ _2313_ sg13g2_a21oi_1
XFILLER_20_422 VPWR VGND sg13g2_fill_2
X_6614_ net225 VGND VPWR _0124_ s0.shift_out\[13\][0] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_21_978 VPWR VGND sg13g2_decap_8
X_3826_ _1405_ net1015 _1404_ VPWR VGND sg13g2_nand2_1
X_6545_ net300 VGND VPWR net658 s0.data_out\[19\]\[2\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3757_ VGND VPWR _2734_ _1332_ _0133_ _1337_ sg13g2_a21oi_1
X_6476_ net1368 _0937_ _0993_ VPWR VGND sg13g2_nor2_1
X_3688_ VGND VPWR net1194 _1276_ _1278_ _1277_ sg13g2_a21oi_1
X_5427_ VPWR _2845_ net465 VGND sg13g2_inv_1
XFILLER_0_838 VPWR VGND sg13g2_decap_8
X_5358_ _2776_ net381 VPWR VGND sg13g2_inv_2
XFILLER_48_809 VPWR VGND sg13g2_decap_8
X_4309_ _1831_ VPWR _1832_ VGND _1822_ _1823_ sg13g2_o21ai_1
X_5289_ _2715_ VPWR _2716_ VGND _2758_ net1142 sg13g2_o21ai_1
XFILLER_12_989 VPWR VGND sg13g2_decap_8
XFILLER_3_698 VPWR VGND sg13g2_decap_8
Xfanout1411 net1415 net1411 VPWR VGND sg13g2_buf_8
Xfanout1422 net1425 net1422 VPWR VGND sg13g2_buf_1
Xfanout1400 net1401 net1400 VPWR VGND sg13g2_buf_8
Xfanout1466 net1467 net1466 VPWR VGND sg13g2_buf_8
Xfanout1433 net1434 net1433 VPWR VGND sg13g2_buf_1
Xfanout1444 net1448 net1444 VPWR VGND sg13g2_buf_8
Xfanout1455 net1456 net1455 VPWR VGND sg13g2_buf_8
Xfanout1488 net1492 net1488 VPWR VGND sg13g2_buf_8
Xfanout1477 net1483 net1477 VPWR VGND sg13g2_buf_8
XFILLER_47_864 VPWR VGND sg13g2_decap_8
XFILLER_46_374 VPWR VGND sg13g2_decap_4
XFILLER_42_580 VPWR VGND sg13g2_fill_2
XFILLER_9_43 VPWR VGND sg13g2_fill_2
XFILLER_14_260 VPWR VGND sg13g2_fill_2
X_4660_ VPWR VGND _2146_ net1460 _2142_ net1452 _2147_ _2140_ sg13g2_a221oi_1
X_3611_ VGND VPWR net1205 s0.data_out\[13\]\[5\] _1207_ _1168_ sg13g2_a21oi_1
XFILLER_30_786 VPWR VGND sg13g2_fill_2
X_4591_ VGND VPWR _2084_ _2086_ _2090_ net1422 sg13g2_a21oi_1
XFILLER_7_960 VPWR VGND sg13g2_decap_8
X_6330_ net1238 net426 _0864_ VPWR VGND sg13g2_and2_1
X_3542_ VGND VPWR _1027_ _1143_ _1144_ net1214 sg13g2_a21oi_1
X_3473_ net1369 _1017_ _1085_ VPWR VGND sg13g2_nor2_1
X_6261_ VGND VPWR net1238 _0796_ _0798_ _0797_ sg13g2_a21oi_1
X_5212_ _2651_ _2626_ _2624_ VPWR VGND sg13g2_nand2b_1
X_6192_ _0741_ _0736_ _0740_ VPWR VGND sg13g2_nand2_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_5143_ net1471 net327 _0274_ VPWR VGND sg13g2_and2_1
XFILLER_38_831 VPWR VGND sg13g2_fill_1
X_5074_ _2525_ net1039 _2524_ VPWR VGND sg13g2_nand2b_1
X_4025_ _1572_ s0.data_out\[9\]\[1\] net1174 VPWR VGND sg13g2_nand2b_1
X_5976_ _0045_ _0542_ _0543_ _2787_ net1352 VPWR VGND sg13g2_a22oi_1
X_4927_ _2388_ net1037 _2389_ _2390_ VPWR VGND sg13g2_a21o_1
X_4858_ net1049 net400 _2331_ VPWR VGND sg13g2_and2_1
X_3809_ _1388_ _1387_ net1413 _1380_ net1404 VPWR VGND sg13g2_a22oi_1
XFILLER_4_407 VPWR VGND sg13g2_fill_1
X_4789_ VGND VPWR _2134_ _2263_ _2264_ net1060 sg13g2_a21oi_1
X_6528_ net318 VGND VPWR _0038_ s0.valid_out\[20\][0] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_6459_ net1369 _0921_ _0980_ VPWR VGND sg13g2_nor2_1
XFILLER_0_635 VPWR VGND sg13g2_decap_8
XFILLER_47_127 VPWR VGND sg13g2_fill_2
XFILLER_29_842 VPWR VGND sg13g2_fill_1
XFILLER_44_801 VPWR VGND sg13g2_decap_8
XFILLER_16_514 VPWR VGND sg13g2_decap_4
XFILLER_29_886 VPWR VGND sg13g2_decap_4
XFILLER_44_867 VPWR VGND sg13g2_fill_2
XFILLER_15_1006 VPWR VGND sg13g2_decap_8
XFILLER_4_985 VPWR VGND sg13g2_decap_8
XFILLER_3_484 VPWR VGND sg13g2_fill_2
Xfanout1230 net1231 net1230 VPWR VGND sg13g2_buf_8
Xfanout1241 net1244 net1241 VPWR VGND sg13g2_buf_2
Xfanout1263 net1264 net1263 VPWR VGND sg13g2_buf_2
Xfanout1274 net1275 net1274 VPWR VGND sg13g2_buf_8
Xfanout1252 net1256 net1252 VPWR VGND sg13g2_buf_8
Xfanout1285 s0.valid_out\[19\][0] net1285 VPWR VGND sg13g2_buf_2
Xfanout1296 net1299 net1296 VPWR VGND sg13g2_buf_8
X_5830_ VGND VPWR _0415_ net1329 net332 sg13g2_or2_1
X_5761_ s0.data_out\[21\]\[0\] s0.data_out\[20\]\[0\] net1297 _0346_ VPWR VGND sg13g2_mux2_1
X_4712_ _2199_ net1077 _2198_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_550 VPWR VGND sg13g2_decap_8
X_5692_ _3086_ _3077_ _3085_ VPWR VGND sg13g2_nand2_1
X_4643_ net1474 VPWR _2133_ VGND _2130_ _2132_ sg13g2_o21ai_1
X_4574_ _2070_ _2071_ _2073_ VPWR VGND _2072_ sg13g2_nand3b_1
X_6313_ net1421 _0839_ _0850_ VPWR VGND sg13g2_nor2_1
X_3525_ _1125_ net1201 _1126_ _1127_ VPWR VGND sg13g2_a21o_1
X_6244_ _0781_ net1248 net426 VPWR VGND sg13g2_nand2_1
X_3456_ _1067_ _1069_ net1432 _1070_ VPWR VGND sg13g2_nand3_1
X_6175_ net1252 net1158 _0724_ VPWR VGND sg13g2_nor2b_1
X_5126_ net1349 _2516_ _2570_ VPWR VGND sg13g2_nor2_1
X_5057_ _2506_ net1030 _2507_ _2508_ VPWR VGND sg13g2_a21o_1
X_4008_ VGND VPWR _2733_ _1559_ _0157_ _1564_ sg13g2_a21oi_1
XFILLER_26_845 VPWR VGND sg13g2_fill_2
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_26_867 VPWR VGND sg13g2_fill_2
X_6677__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_41_826 VPWR VGND sg13g2_fill_1
X_5959_ _0530_ VPWR _0531_ VGND net1472 net672 sg13g2_o21ai_1
XFILLER_21_583 VPWR VGND sg13g2_fill_1
XFILLER_5_727 VPWR VGND sg13g2_decap_8
XFILLER_20_75 VPWR VGND sg13g2_fill_2
XFILLER_1_933 VPWR VGND sg13g2_decap_8
XFILLER_49_926 VPWR VGND sg13g2_decap_8
Xhold40 s0.shift_out\[10\][0] VPWR VGND net360 sg13g2_dlygate4sd3_1
Xhold51 s0.data_out\[8\]\[7\] VPWR VGND net371 sg13g2_dlygate4sd3_1
Xhold73 _0013_ VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold62 _0006_ VPWR VGND net382 sg13g2_dlygate4sd3_1
Xhold84 s0.data_out\[6\]\[7\] VPWR VGND net404 sg13g2_dlygate4sd3_1
Xhold95 _1288_ VPWR VGND net415 sg13g2_dlygate4sd3_1
XFILLER_29_672 VPWR VGND sg13g2_decap_8
XFILLER_40_892 VPWR VGND sg13g2_fill_1
XFILLER_6_77 VPWR VGND sg13g2_fill_1
X_4290_ VGND VPWR _1696_ _1812_ _1813_ net1110 sg13g2_a21oi_1
XFILLER_6_1026 VPWR VGND sg13g2_fill_2
Xfanout1082 net1084 net1082 VPWR VGND sg13g2_buf_8
Xfanout1071 net706 net1071 VPWR VGND sg13g2_buf_8
XFILLER_13_2 VPWR VGND sg13g2_fill_1
Xfanout1060 net1063 net1060 VPWR VGND sg13g2_buf_8
XFILLER_48_970 VPWR VGND sg13g2_decap_8
Xfanout1093 s0.valid_out\[6\][0] net1093 VPWR VGND sg13g2_buf_1
XFILLER_26_108 VPWR VGND sg13g2_decap_8
XFILLER_35_664 VPWR VGND sg13g2_fill_1
X_5813_ _0398_ net1299 s0.data_out\[20\]\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_22_314 VPWR VGND sg13g2_fill_2
XFILLER_23_837 VPWR VGND sg13g2_fill_1
XFILLER_34_185 VPWR VGND sg13g2_fill_1
X_5744_ _0328_ VPWR _0332_ VGND net649 net1296 sg13g2_o21ai_1
X_5675_ _3066_ _3067_ _3069_ VPWR VGND _3068_ sg13g2_nand3b_1
X_4626_ VPWR _0221_ _2118_ VGND sg13g2_inv_1
X_4557_ _2056_ net1082 net488 VPWR VGND sg13g2_nand2_1
X_3508_ _1112_ VPWR _1113_ VGND net1205 _1106_ sg13g2_o21ai_1
X_4488_ net998 _2862_ _1995_ VPWR VGND sg13g2_nor2_1
X_6227_ _0768_ VPWR _0769_ VGND net1470 net534 sg13g2_o21ai_1
X_3439_ VPWR _1053_ _1052_ VGND sg13g2_inv_1
X_6158_ _0705_ net1249 _0706_ _0707_ VPWR VGND sg13g2_a21o_1
XFILLER_46_918 VPWR VGND sg13g2_decap_8
X_5109_ VPWR _0266_ _2556_ VGND sg13g2_inv_1
X_6683__151 VPWR VGND net151 sg13g2_tiehi
X_6089_ net1265 net410 _0646_ VPWR VGND sg13g2_and2_1
XFILLER_17_108 VPWR VGND sg13g2_decap_4
XFILLER_45_439 VPWR VGND sg13g2_fill_1
XFILLER_41_612 VPWR VGND sg13g2_fill_1
XFILLER_13_303 VPWR VGND sg13g2_fill_2
XFILLER_40_111 VPWR VGND sg13g2_fill_2
XFILLER_13_336 VPWR VGND sg13g2_fill_1
XFILLER_15_64 VPWR VGND sg13g2_fill_2
XFILLER_41_678 VPWR VGND sg13g2_decap_8
XFILLER_22_870 VPWR VGND sg13g2_fill_1
X_6690__144 VPWR VGND net144 sg13g2_tiehi
Xoutput6 net6 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_5_557 VPWR VGND sg13g2_fill_1
XFILLER_31_96 VPWR VGND sg13g2_fill_2
XFILLER_1_730 VPWR VGND sg13g2_decap_8
XFILLER_49_723 VPWR VGND sg13g2_decap_8
XFILLER_0_262 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_320 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_17_642 VPWR VGND sg13g2_fill_1
XFILLER_45_984 VPWR VGND sg13g2_decap_8
XFILLER_13_881 VPWR VGND sg13g2_fill_1
X_3790_ net1440 _1368_ _1369_ VPWR VGND sg13g2_nor2_1
XFILLER_32_678 VPWR VGND sg13g2_decap_4
XFILLER_13_892 VPWR VGND sg13g2_decap_8
X_5460_ VPWR _2878_ net434 VGND sg13g2_inv_1
X_4411_ _1922_ s0.data_out\[6\]\[1\] net1105 VPWR VGND sg13g2_nand2b_1
X_5391_ VPWR _2809_ net475 VGND sg13g2_inv_1
X_4342_ VGND VPWR _1746_ _1864_ _1865_ net1114 sg13g2_a21oi_1
X_4273_ net1481 VPWR _1799_ VGND _1796_ _1798_ sg13g2_o21ai_1
X_6667__168 VPWR VGND net168 sg13g2_tiehi
X_6012_ _0571_ net1266 _0572_ _0573_ VPWR VGND sg13g2_a21o_1
.ends

