* NGSPICE file created from heichips25_top_sorter.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

.subckt heichips25_top_sorter VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_277 VPWR VGND sg13g2_fill_2
XFILLER_28_918 VPWR VGND sg13g2_fill_2
X_7963_ net191 VGND VPWR _0097_ s0.valid_out\[0\][0] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_6914_ VGND VPWR _2719_ _2721_ _2724_ net1679 sg13g2_a21oi_1
X_7894_ net115 VGND VPWR _0028_ s0.data_out\[6\]\[0\] clknet_leaf_6_clk sg13g2_dfrbpq_2
XFILLER_22_133 VPWR VGND sg13g2_fill_2
X_6845_ _2654_ VPWR _2655_ VGND net1266 _3523_ sg13g2_o21ai_1
XFILLER_35_494 VPWR VGND sg13g2_decap_4
X_3988_ VPWR _3364_ net416 VGND sg13g2_inv_1
X_6776_ _2598_ net1176 _2597_ VPWR VGND sg13g2_nand2_1
XFILLER_10_306 VPWR VGND sg13g2_decap_8
XFILLER_11_818 VPWR VGND sg13g2_fill_1
XFILLER_11_829 VPWR VGND sg13g2_decap_4
X_5727_ _1652_ net1409 net612 VPWR VGND sg13g2_nand2_1
X_5658_ net1425 VPWR _1594_ VGND _1535_ _1593_ sg13g2_o21ai_1
X_4609_ VGND VPWR net1526 _0639_ _0642_ _0641_ sg13g2_a21oi_1
X_5589_ _1526_ net1419 net702 VPWR VGND sg13g2_nand2_1
Xhold351 s0.data_out\[10\]\[6\] VPWR VGND net720 sg13g2_dlygate4sd3_1
Xhold362 s0.data_out\[9\]\[6\] VPWR VGND net731 sg13g2_dlygate4sd3_1
X_7639__47 VPWR VGND net47 sg13g2_tiehi
Xhold340 s0.data_out\[19\]\[1\] VPWR VGND net709 sg13g2_dlygate4sd3_1
X_7328_ net1239 VPWR _3094_ VGND _3034_ _3093_ sg13g2_o21ai_1
Xhold395 s0.data_out\[23\]\[4\] VPWR VGND net764 sg13g2_dlygate4sd3_1
Xhold384 s0.data_out\[17\]\[6\] VPWR VGND net753 sg13g2_dlygate4sd3_1
Xhold373 s0.data_out\[16\]\[6\] VPWR VGND net742 sg13g2_dlygate4sd3_1
X_7259_ s0.data_out\[3\]\[7\] s0.data_out\[2\]\[7\] net1235 _3033_ VPWR VGND sg13g2_mux2_1
X_7887__123 VPWR VGND net123 sg13g2_tiehi
XFILLER_46_737 VPWR VGND sg13g2_decap_8
XFILLER_26_30 VPWR VGND sg13g2_fill_2
XFILLER_26_63 VPWR VGND sg13g2_decap_8
XFILLER_42_954 VPWR VGND sg13g2_decap_8
XFILLER_13_177 VPWR VGND sg13g2_fill_1
XFILLER_42_73 VPWR VGND sg13g2_fill_2
XFILLER_10_851 VPWR VGND sg13g2_fill_1
XFILLER_3_56 VPWR VGND sg13g2_fill_1
XFILLER_49_542 VPWR VGND sg13g2_decap_8
XFILLER_37_704 VPWR VGND sg13g2_fill_2
X_4960_ _0958_ net1481 net497 VPWR VGND sg13g2_nand2_1
XFILLER_17_450 VPWR VGND sg13g2_fill_2
XFILLER_17_483 VPWR VGND sg13g2_fill_1
XFILLER_18_995 VPWR VGND sg13g2_decap_8
X_4891_ _0900_ _0899_ net1500 VPWR VGND sg13g2_nand2b_1
X_6630_ VGND VPWR _2343_ _2463_ _2464_ net1294 sg13g2_a21oi_1
X_7803__213 VPWR VGND net213 sg13g2_tiehi
X_6561_ _3394_ _3512_ _2404_ VPWR VGND sg13g2_nor2_1
X_5512_ net1426 net1345 _1461_ VPWR VGND sg13g2_nor2b_1
X_6492_ s0.data_out\[8\]\[0\] s0.data_out\[9\]\[0\] net1315 _2338_ VPWR VGND sg13g2_mux2_1
X_5443_ net1429 _1389_ _1395_ VPWR VGND sg13g2_nor2_1
X_5374_ _1334_ _1332_ _1335_ VPWR VGND _1333_ sg13g2_nand3b_1
X_4325_ VGND VPWR _3372_ _0379_ _0121_ _0384_ sg13g2_a21oi_1
X_7113_ VPWR VGND _2897_ _2898_ _2890_ net1571 _2899_ _2883_ sg13g2_a221oi_1
XFILLER_47_18 VPWR VGND sg13g2_fill_1
X_4256_ _3620_ net1554 net491 VPWR VGND sg13g2_nand2_1
X_7044_ VGND VPWR _2842_ net1566 net378 sg13g2_or2_1
X_7810__206 VPWR VGND net206 sg13g2_tiehi
XFILLER_41_1024 VPWR VGND sg13g2_decap_4
X_4187_ VGND VPWR net1633 net1554 _3554_ _3553_ sg13g2_a21oi_1
X_7946_ net59 VGND VPWR net521 s0.data_out\[2\]\[4\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_7877_ net134 VGND VPWR net562 s0.data_out\[8\]\[7\] clknet_leaf_15_clk sg13g2_dfrbpq_2
XFILLER_24_965 VPWR VGND sg13g2_decap_8
X_6828_ VPWR _0022_ _2642_ VGND sg13g2_inv_1
X_6759_ VGND VPWR net1285 _2578_ _2581_ _2580_ sg13g2_a21oi_1
XFILLER_10_169 VPWR VGND sg13g2_fill_1
XFILLER_3_858 VPWR VGND sg13g2_decap_8
Xhold170 _0191_ VPWR VGND net539 sg13g2_dlygate4sd3_1
Xhold192 s0.data_out\[8\]\[7\] VPWR VGND net561 sg13g2_dlygate4sd3_1
Xfanout1604 net1605 net1604 VPWR VGND sg13g2_buf_8
Xfanout1615 net1616 net1615 VPWR VGND sg13g2_buf_8
Xhold181 _0337_ VPWR VGND net550 sg13g2_dlygate4sd3_1
Xfanout1648 net1649 net1648 VPWR VGND sg13g2_buf_8
Xfanout1637 net1638 net1637 VPWR VGND sg13g2_buf_8
Xfanout1626 net1627 net1626 VPWR VGND sg13g2_buf_8
Xfanout1659 net1662 net1659 VPWR VGND sg13g2_buf_8
XFILLER_18_258 VPWR VGND sg13g2_fill_1
XFILLER_26_291 VPWR VGND sg13g2_fill_1
XFILLER_42_762 VPWR VGND sg13g2_fill_2
XFILLER_14_442 VPWR VGND sg13g2_fill_1
XFILLER_14_497 VPWR VGND sg13g2_fill_2
XFILLER_30_979 VPWR VGND sg13g2_decap_8
XFILLER_6_696 VPWR VGND sg13g2_fill_2
XFILLER_38_4 VPWR VGND sg13g2_fill_1
X_5090_ VGND VPWR _1075_ _1074_ net1697 sg13g2_or2_1
X_4110_ VPWR _3486_ net624 VGND sg13g2_inv_1
X_4041_ VPWR _3417_ net559 VGND sg13g2_inv_1
X_7800_ net216 VGND VPWR _0278_ s0.valid_out\[13\][0] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_37_578 VPWR VGND sg13g2_fill_2
X_5992_ _1892_ VPWR _1893_ VGND net1389 _3484_ sg13g2_o21ai_1
X_4943_ net1483 _0825_ _0943_ VPWR VGND sg13g2_nor2_1
XFILLER_17_291 VPWR VGND sg13g2_fill_1
X_7731_ net291 VGND VPWR _0209_ s0.data_out\[19\]\[0\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_7662_ net366 VGND VPWR _0140_ s0.data_out\[25\]\[3\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_4874_ net1663 _0880_ _0883_ VPWR VGND sg13g2_nor2_1
X_6613_ _2447_ s0.data_out\[7\]\[1\] net1301 VPWR VGND sg13g2_nand2b_1
X_7593_ _3393_ net570 net1214 _3331_ VPWR VGND sg13g2_nand3_1
X_6544_ _2387_ _2388_ _2389_ _2390_ VPWR VGND sg13g2_or3_1
X_7955__308 VPWR VGND net308 sg13g2_tiehi
X_6475_ net1295 net1351 _2321_ VPWR VGND sg13g2_nor2b_1
X_5426_ net1624 _1348_ _1381_ VPWR VGND sg13g2_nor2_1
X_7738__284 VPWR VGND net284 sg13g2_tiehi
XFILLER_0_817 VPWR VGND sg13g2_decap_8
X_5357_ _1318_ net1444 s0.data_out\[17\]\[6\] VPWR VGND sg13g2_nand2_1
X_4308_ net1558 VPWR _0370_ VGND _3610_ _0369_ sg13g2_o21ai_1
X_5288_ net1203 _3461_ _1258_ VPWR VGND sg13g2_nor2_1
X_4239_ _3601_ net1544 _3602_ _3603_ VPWR VGND sg13g2_a21o_1
X_7027_ VGND VPWR net1259 _2822_ _2825_ _2824_ sg13g2_a21oi_1
XFILLER_28_501 VPWR VGND sg13g2_fill_1
X_7884__126 VPWR VGND net126 sg13g2_tiehi
X_7929_ net77 VGND VPWR _0063_ s0.shift_out\[3\][0] clknet_leaf_8_clk sg13g2_dfrbpq_2
XFILLER_11_456 VPWR VGND sg13g2_fill_1
XFILLER_7_449 VPWR VGND sg13g2_fill_1
XFILLER_23_97 VPWR VGND sg13g2_fill_2
XFILLER_48_1019 VPWR VGND sg13g2_decap_8
Xfanout1423 net1424 net1423 VPWR VGND sg13g2_buf_2
Xfanout1412 net1413 net1412 VPWR VGND sg13g2_buf_8
Xfanout1401 net1402 net1401 VPWR VGND sg13g2_buf_8
Xfanout1456 net820 net1456 VPWR VGND sg13g2_buf_8
Xfanout1445 net1446 net1445 VPWR VGND sg13g2_buf_8
Xfanout1434 net1435 net1434 VPWR VGND sg13g2_buf_1
Xfanout1467 s0.valid_out\[19\][0] net1467 VPWR VGND sg13g2_buf_8
Xfanout1489 net1490 net1489 VPWR VGND sg13g2_buf_8
Xfanout1478 net1481 net1478 VPWR VGND sg13g2_buf_8
XFILLER_47_843 VPWR VGND sg13g2_decap_8
X_7800__216 VPWR VGND net216 sg13g2_tiehi
XFILLER_9_99 VPWR VGND sg13g2_fill_1
X_4590_ _0621_ net1510 _0622_ _0623_ VPWR VGND sg13g2_a21o_1
XFILLER_30_776 VPWR VGND sg13g2_fill_2
XFILLER_7_983 VPWR VGND sg13g2_decap_8
X_6260_ _2136_ _2133_ _2137_ VPWR VGND _2135_ sg13g2_nand3b_1
X_6191_ _2072_ VPWR _2073_ VGND net1740 net723 sg13g2_o21ai_1
XFILLER_9_1002 VPWR VGND sg13g2_decap_8
X_5211_ VGND VPWR _1184_ _1183_ net1697 sg13g2_or2_1
X_5142_ net1457 net1340 _1127_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_0 VPWR VGND sg13g2_fill_1
X_5073_ _1060_ VPWR _1061_ VGND net1473 _0941_ sg13g2_o21ai_1
X_4024_ VPWR _3400_ net472 VGND sg13g2_inv_1
X_5975_ s0.data_out\[12\]\[0\] s0.data_out\[13\]\[0\] net1397 _1876_ VPWR VGND sg13g2_mux2_1
X_7714_ net310 VGND VPWR _0192_ s0.genblk1\[20\].modules.bubble clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_4926_ VPWR _0177_ _0929_ VGND sg13g2_inv_1
X_7645_ net40 VGND VPWR _0123_ s0.genblk1\[25\].modules.bubble clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_4857_ _0865_ VPWR _0866_ VGND _0856_ _0857_ sg13g2_o21ai_1
X_7576_ net1720 VPWR _3317_ VGND net1214 net1209 sg13g2_o21ai_1
X_6527_ _2373_ net1309 _2372_ VPWR VGND sg13g2_nand2b_1
XFILLER_5_909 VPWR VGND sg13g2_decap_8
X_4788_ _0805_ VPWR _0806_ VGND net1728 net619 sg13g2_o21ai_1
X_6458_ _0331_ _2306_ _2307_ _3501_ net1610 VPWR VGND sg13g2_a22oi_1
X_6389_ _2245_ net1311 _2246_ _2247_ VPWR VGND sg13g2_a21o_1
XFILLER_0_603 VPWR VGND sg13g2_decap_8
X_5409_ _1367_ VPWR _1368_ VGND net1743 net808 sg13g2_o21ai_1
X_7751__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_29_821 VPWR VGND sg13g2_fill_1
XFILLER_28_375 VPWR VGND sg13g2_fill_1
XFILLER_44_835 VPWR VGND sg13g2_fill_1
XFILLER_16_559 VPWR VGND sg13g2_fill_2
XFILLER_12_743 VPWR VGND sg13g2_decap_4
XFILLER_34_85 VPWR VGND sg13g2_fill_2
XFILLER_4_920 VPWR VGND sg13g2_decap_8
XFILLER_4_997 VPWR VGND sg13g2_decap_8
Xfanout1220 net529 net1220 VPWR VGND sg13g2_buf_8
Xfanout1231 s0.shift_out\[2\][0] net1231 VPWR VGND sg13g2_buf_2
Xfanout1264 net1265 net1264 VPWR VGND sg13g2_buf_1
Xfanout1253 net1257 net1253 VPWR VGND sg13g2_buf_8
Xfanout1242 net1243 net1242 VPWR VGND sg13g2_buf_8
Xfanout1297 net1299 net1297 VPWR VGND sg13g2_buf_2
Xfanout1286 net1288 net1286 VPWR VGND sg13g2_buf_8
Xfanout1275 net1277 net1275 VPWR VGND sg13g2_buf_2
XFILLER_22_518 VPWR VGND sg13g2_fill_2
X_5760_ VGND VPWR net1404 _1683_ _1685_ _1684_ sg13g2_a21oi_1
X_7728__294 VPWR VGND net294 sg13g2_tiehi
X_4711_ _0732_ net1503 s0.data_out\[22\]\[2\] VPWR VGND sg13g2_nand2_1
X_5691_ net1417 VPWR _1619_ VGND net1645 net1405 sg13g2_o21ai_1
X_7430_ VPWR _0078_ _3188_ VGND sg13g2_inv_1
X_4642_ net1688 _0642_ _0675_ VPWR VGND sg13g2_nor2_1
X_4573_ net1509 _0603_ _0609_ VPWR VGND sg13g2_nor2_1
X_7361_ s0.data_out\[1\]\[0\] s0.data_out\[2\]\[0\] net1236 _3123_ VPWR VGND sg13g2_mux2_1
X_6312_ _2181_ net1739 _2182_ VPWR VGND _2124_ sg13g2_nand3b_1
X_7292_ VGND VPWR _3051_ _3064_ _3066_ _3065_ sg13g2_a21oi_1
X_6243_ s0.data_out\[11\]\[6\] s0.data_out\[10\]\[6\] net1363 _2120_ VPWR VGND sg13g2_mux2_1
X_6174_ _0295_ _2058_ _2059_ _3490_ net1611 VPWR VGND sg13g2_a22oi_1
X_5125_ _1108_ net1457 _1109_ _1110_ VPWR VGND sg13g2_a21o_1
X_7735__287 VPWR VGND net287 sg13g2_tiehi
XFILLER_29_106 VPWR VGND sg13g2_fill_1
X_5056_ net1468 net509 _1048_ VPWR VGND sg13g2_and2_1
X_4007_ net1366 _3383_ VPWR VGND sg13g2_inv_4
X_7881__129 VPWR VGND net129 sg13g2_tiehi
XFILLER_38_1007 VPWR VGND sg13g2_decap_8
X_5958_ _1858_ VPWR _1859_ VGND net1386 _3486_ sg13g2_o21ai_1
X_4909_ net1487 s0.data_out\[21\]\[1\] _0916_ VPWR VGND sg13g2_and2_1
X_5889_ _1802_ _3381_ _1801_ VPWR VGND sg13g2_nand2_1
X_7628_ net1721 net447 _3358_ VPWR VGND sg13g2_nor2_1
X_7559_ VPWR _0092_ _3303_ VGND sg13g2_inv_1
XFILLER_5_728 VPWR VGND sg13g2_fill_1
XFILLER_1_901 VPWR VGND sg13g2_decap_8
XFILLER_20_87 VPWR VGND sg13g2_decap_4
XFILLER_1_978 VPWR VGND sg13g2_decap_8
XFILLER_49_927 VPWR VGND sg13g2_decap_8
Xhold30 _0024_ VPWR VGND net399 sg13g2_dlygate4sd3_1
Xhold41 _0157_ VPWR VGND net410 sg13g2_dlygate4sd3_1
Xhold63 _0436_ VPWR VGND net432 sg13g2_dlygate4sd3_1
Xhold52 s0.was_valid_out\[2\][0] VPWR VGND net421 sg13g2_dlygate4sd3_1
Xhold74 s0.data_out\[10\]\[3\] VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold96 _0127_ VPWR VGND net465 sg13g2_dlygate4sd3_1
XFILLER_17_813 VPWR VGND sg13g2_fill_2
Xhold85 s0.shift_out\[4\][0] VPWR VGND net454 sg13g2_dlygate4sd3_1
XFILLER_44_632 VPWR VGND sg13g2_decap_4
XFILLER_44_654 VPWR VGND sg13g2_fill_1
XFILLER_43_131 VPWR VGND sg13g2_fill_1
XFILLER_16_367 VPWR VGND sg13g2_fill_1
XFILLER_44_687 VPWR VGND sg13g2_fill_2
XFILLER_31_315 VPWR VGND sg13g2_fill_2
XFILLER_31_348 VPWR VGND sg13g2_fill_2
XFILLER_6_45 VPWR VGND sg13g2_fill_2
XFILLER_39_448 VPWR VGND sg13g2_fill_2
X_7689__337 VPWR VGND net337 sg13g2_tiehi
X_6930_ net1270 VPWR _2738_ VGND _2656_ _2737_ sg13g2_o21ai_1
X_6861_ VGND VPWR net1261 _2669_ _2671_ _2670_ sg13g2_a21oi_1
X_6792_ _2608_ VPWR _2614_ VGND _2600_ _2610_ sg13g2_o21ai_1
XFILLER_23_838 VPWR VGND sg13g2_fill_1
X_5812_ net1404 s0.data_out\[14\]\[6\] _1730_ VPWR VGND sg13g2_and2_1
X_5743_ VGND VPWR _1550_ _1667_ _1668_ net1417 sg13g2_a21oi_1
X_5674_ net1415 net777 _1606_ VPWR VGND sg13g2_and2_1
X_4625_ _0658_ _0657_ net1660 _0650_ net1650 VPWR VGND sg13g2_a22oi_1
X_7741__280 VPWR VGND net280 sg13g2_tiehi
X_7413_ _3100_ VPWR _3175_ VGND _3151_ _3153_ sg13g2_o21ai_1
X_7344_ s0.data_out\[2\]\[2\] s0.data_out\[1\]\[2\] net1226 _3106_ VPWR VGND sg13g2_mux2_1
X_4556_ _0594_ VPWR _0595_ VGND net1725 net774 sg13g2_o21ai_1
X_4487_ net1520 net1328 _0532_ VPWR VGND sg13g2_nor2b_1
X_7275_ net1668 _3048_ _3049_ VPWR VGND sg13g2_nor2_1
X_6226_ net1321 net1358 _2103_ VPWR VGND sg13g2_nor2b_1
X_6157_ _2023_ _2045_ _2046_ VPWR VGND sg13g2_nor2b_1
X_5108_ net1459 net1168 _1093_ VPWR VGND sg13g2_nor2_1
XFILLER_39_971 VPWR VGND sg13g2_decap_8
X_6088_ _1975_ net1367 _1976_ _1977_ VPWR VGND sg13g2_a21o_1
XFILLER_38_492 VPWR VGND sg13g2_fill_1
XFILLER_38_470 VPWR VGND sg13g2_fill_2
X_5039_ _1034_ VPWR _1035_ VGND net1178 _1033_ sg13g2_o21ai_1
XFILLER_25_120 VPWR VGND sg13g2_fill_2
XFILLER_15_87 VPWR VGND sg13g2_fill_1
XFILLER_31_53 VPWR VGND sg13g2_fill_1
Xoutput7 net7 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_49_724 VPWR VGND sg13g2_decap_8
XFILLER_0_252 VPWR VGND sg13g2_decap_4
XFILLER_1_775 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_fill_2
XFILLER_45_963 VPWR VGND sg13g2_decap_8
XFILLER_16_120 VPWR VGND sg13g2_fill_1
X_4410_ net1581 _0398_ _0465_ VPWR VGND sg13g2_nor2_1
X_5390_ net1674 _1349_ _1351_ VPWR VGND sg13g2_nor2_1
X_7695__330 VPWR VGND net330 sg13g2_tiehi
X_4341_ VGND VPWR _3572_ _0397_ _0398_ net1552 sg13g2_a21oi_1
X_7648__37 VPWR VGND net37 sg13g2_tiehi
XFILLER_28_1006 VPWR VGND sg13g2_decap_8
X_4272_ _3635_ VPWR _3636_ VGND net1677 _3633_ sg13g2_o21ai_1
X_7060_ net1259 VPWR _2854_ VGND _2795_ _2853_ sg13g2_o21ai_1
X_6011_ s0.data_out\[13\]\[6\] s0.data_out\[12\]\[6\] net1389 _1912_ VPWR VGND sg13g2_mux2_1
X_7962_ net217 VGND VPWR net508 s0.was_valid_out\[0\][0] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_6913_ _2723_ _2714_ _2722_ VPWR VGND sg13g2_nand2_1
X_7893_ net116 VGND VPWR _0027_ s0.shift_out\[6\][0] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_35_451 VPWR VGND sg13g2_fill_1
XFILLER_35_484 VPWR VGND sg13g2_fill_1
X_6844_ _2654_ net1266 net752 VPWR VGND sg13g2_nand2_1
X_3987_ VPWR _3363_ net398 VGND sg13g2_inv_1
X_6775_ s0.data_out\[6\]\[4\] s0.data_out\[7\]\[4\] net1291 _2597_ VPWR VGND sg13g2_mux2_1
X_5726_ net1707 _1634_ _1651_ VPWR VGND sg13g2_nor2_1
X_5657_ net1412 s0.data_out\[15\]\[0\] _1593_ VPWR VGND sg13g2_and2_1
X_4608_ VGND VPWR _0519_ _0640_ _0641_ net1526 sg13g2_a21oi_1
X_5588_ net1697 _1524_ _1525_ VPWR VGND sg13g2_nor2_1
Xhold330 _0153_ VPWR VGND net699 sg13g2_dlygate4sd3_1
X_4539_ net1522 s0.data_out\[24\]\[2\] _0581_ VPWR VGND sg13g2_and2_1
Xhold341 _0210_ VPWR VGND net710 sg13g2_dlygate4sd3_1
Xhold352 s0.data_out\[2\]\[0\] VPWR VGND net721 sg13g2_dlygate4sd3_1
X_7327_ net1189 _3538_ _3093_ VPWR VGND sg13g2_nor2_1
Xhold385 _1504_ VPWR VGND net754 sg13g2_dlygate4sd3_1
Xhold374 _1615_ VPWR VGND net743 sg13g2_dlygate4sd3_1
Xhold363 s0.data_out\[13\]\[0\] VPWR VGND net732 sg13g2_dlygate4sd3_1
Xhold396 s0.data_out\[15\]\[3\] VPWR VGND net765 sg13g2_dlygate4sd3_1
X_7258_ _3032_ net1236 net568 VPWR VGND sg13g2_nand2_1
X_6209_ net388 net1739 _0303_ VPWR VGND sg13g2_and2_1
X_7189_ VGND VPWR net1173 _2924_ _2970_ net1586 sg13g2_a21oi_1
XFILLER_46_716 VPWR VGND sg13g2_decap_8
XFILLER_26_20 VPWR VGND sg13g2_fill_1
XFILLER_27_985 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_42_933 VPWR VGND sg13g2_decap_8
XFILLER_5_344 VPWR VGND sg13g2_fill_2
XFILLER_1_550 VPWR VGND sg13g2_fill_1
XFILLER_49_521 VPWR VGND sg13g2_decap_8
XFILLER_49_598 VPWR VGND sg13g2_decap_8
XFILLER_3_1019 VPWR VGND sg13g2_decap_8
XFILLER_36_259 VPWR VGND sg13g2_fill_2
XFILLER_45_771 VPWR VGND sg13g2_decap_8
XFILLER_18_974 VPWR VGND sg13g2_decap_8
X_4890_ s0.data_out\[21\]\[4\] s0.data_out\[22\]\[4\] net1506 _0899_ VPWR VGND sg13g2_mux2_1
XFILLER_33_988 VPWR VGND sg13g2_decap_8
X_6560_ _0337_ _2402_ _2403_ _3506_ net1608 VPWR VGND sg13g2_a22oi_1
XFILLER_32_498 VPWR VGND sg13g2_fill_2
X_5511_ _1457_ _1459_ net1674 _1460_ VPWR VGND sg13g2_nand3_1
X_6491_ _2337_ net1305 _2336_ VPWR VGND sg13g2_nand2b_1
X_5442_ _1391_ VPWR _1394_ VGND s0.was_valid_out\[16\][0] net1434 sg13g2_o21ai_1
X_5373_ VGND VPWR _1334_ _1331_ net1656 sg13g2_or2_1
X_4324_ net1714 VPWR _0384_ VGND _0381_ _0383_ sg13g2_o21ai_1
X_7112_ VGND VPWR _2887_ _2889_ _2898_ net1701 sg13g2_a21oi_1
X_7043_ _2839_ _2840_ _2841_ VPWR VGND sg13g2_nor2_1
XFILLER_41_1003 VPWR VGND sg13g2_decap_8
X_4255_ net1558 _3617_ _3618_ _3619_ VPWR VGND sg13g2_nor3_1
X_4186_ net1559 VPWR _3553_ VGND net1639 net1544 sg13g2_o21ai_1
X_7945_ net60 VGND VPWR net736 s0.data_out\[2\]\[3\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_36_771 VPWR VGND sg13g2_fill_2
X_7876_ net135 VGND VPWR net609 s0.data_out\[8\]\[6\] clknet_leaf_15_clk sg13g2_dfrbpq_2
XFILLER_36_793 VPWR VGND sg13g2_fill_1
X_6827_ _2641_ VPWR _2642_ VGND net1729 net801 sg13g2_o21ai_1
X_6758_ VGND VPWR _2474_ _2579_ _2580_ net1285 sg13g2_a21oi_1
X_5709_ VGND VPWR net1414 _1631_ _1634_ _1633_ sg13g2_a21oi_1
X_6689_ net1294 VPWR _2519_ VGND _2461_ _2518_ sg13g2_o21ai_1
XFILLER_3_826 VPWR VGND sg13g2_decap_8
Xhold160 s0.shift_out\[1\][0] VPWR VGND net529 sg13g2_dlygate4sd3_1
Xhold171 s0.data_out\[12\]\[7\] VPWR VGND net540 sg13g2_dlygate4sd3_1
Xhold193 _0011_ VPWR VGND net562 sg13g2_dlygate4sd3_1
Xfanout1605 net1616 net1605 VPWR VGND sg13g2_buf_8
Xhold182 s0.data_out\[11\]\[2\] VPWR VGND net551 sg13g2_dlygate4sd3_1
Xfanout1638 net1 net1638 VPWR VGND sg13g2_buf_8
Xfanout1649 net1652 net1649 VPWR VGND sg13g2_buf_8
Xfanout1616 net1632 net1616 VPWR VGND sg13g2_buf_8
Xfanout1627 net1628 net1627 VPWR VGND sg13g2_buf_8
X_7635__51 VPWR VGND net51 sg13g2_tiehi
XFILLER_46_502 VPWR VGND sg13g2_fill_1
XFILLER_46_546 VPWR VGND sg13g2_fill_1
XFILLER_26_270 VPWR VGND sg13g2_fill_1
XFILLER_18_1016 VPWR VGND sg13g2_decap_8
XFILLER_18_1027 VPWR VGND sg13g2_fill_2
XFILLER_6_642 VPWR VGND sg13g2_fill_1
XFILLER_5_130 VPWR VGND sg13g2_decap_8
X_7692__333 VPWR VGND net333 sg13g2_tiehi
XFILLER_25_1009 VPWR VGND sg13g2_decap_8
X_4040_ VPWR _3416_ net621 VGND sg13g2_inv_1
XFILLER_25_719 VPWR VGND sg13g2_decap_4
X_5991_ _1892_ net1387 s0.data_out\[12\]\[4\] VPWR VGND sg13g2_nand2_1
X_4942_ _0940_ _0941_ _0942_ VPWR VGND sg13g2_nor2_2
X_7730_ net292 VGND VPWR _0208_ s0.shift_out\[19\][0] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_7661_ net367 VGND VPWR _0139_ s0.data_out\[25\]\[2\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_4873_ VPWR _0882_ _0881_ VGND sg13g2_inv_1
XFILLER_21_925 VPWR VGND sg13g2_fill_2
X_6612_ _2444_ net1282 _2445_ _2446_ VPWR VGND sg13g2_a21o_1
X_7592_ _3330_ net1208 net1356 VPWR VGND sg13g2_nand2_1
XFILLER_20_457 VPWR VGND sg13g2_fill_1
X_7877__134 VPWR VGND net134 sg13g2_tiehi
X_6543_ net1691 _2349_ _2389_ VPWR VGND sg13g2_nor2_1
X_6474_ s0.data_out\[9\]\[2\] s0.data_out\[8\]\[2\] net1301 _2320_ VPWR VGND sg13g2_mux2_1
X_5425_ net1450 VPWR _1380_ VGND _1345_ _1379_ sg13g2_o21ai_1
X_5356_ _1316_ VPWR _1317_ VGND net1573 _1291_ sg13g2_o21ai_1
X_4307_ net1544 s0.data_out\[26\]\[6\] _0369_ VPWR VGND sg13g2_and2_1
X_5287_ _0210_ _1256_ _1257_ _3456_ net1619 VPWR VGND sg13g2_a22oi_1
X_4238_ net1544 net1328 _3602_ VPWR VGND sg13g2_nor2b_1
X_7026_ VGND VPWR _2716_ _2823_ _2824_ net1263 sg13g2_a21oi_1
XFILLER_28_513 VPWR VGND sg13g2_fill_1
X_7632__54 VPWR VGND net54 sg13g2_tiehi
X_4169_ s0.data_out\[27\]\[0\] net1166 _3545_ VPWR VGND sg13g2_nor2_1
X_7928_ net78 VGND VPWR _0062_ s0.genblk1\[2\].modules.bubble clknet_leaf_8_clk sg13g2_dfrbpq_1
X_7859_ net153 VGND VPWR net550 s0.data_out\[9\]\[1\] clknet_leaf_38_clk sg13g2_dfrbpq_2
XFILLER_23_76 VPWR VGND sg13g2_fill_2
XFILLER_20_991 VPWR VGND sg13g2_decap_8
XFILLER_3_601 VPWR VGND sg13g2_fill_2
Xfanout1413 net1414 net1413 VPWR VGND sg13g2_buf_2
Xfanout1402 net1403 net1402 VPWR VGND sg13g2_buf_8
Xfanout1457 net1460 net1457 VPWR VGND sg13g2_buf_8
Xfanout1446 net823 net1446 VPWR VGND sg13g2_buf_8
Xfanout1435 s0.valid_out\[16\][0] net1435 VPWR VGND sg13g2_buf_8
Xfanout1424 net1425 net1424 VPWR VGND sg13g2_buf_8
XFILLER_47_822 VPWR VGND sg13g2_decap_8
Xfanout1468 net1477 net1468 VPWR VGND sg13g2_buf_8
Xfanout1479 net1481 net1479 VPWR VGND sg13g2_buf_1
XFILLER_47_899 VPWR VGND sg13g2_decap_8
XFILLER_14_240 VPWR VGND sg13g2_fill_2
XFILLER_9_67 VPWR VGND sg13g2_fill_1
XFILLER_30_733 VPWR VGND sg13g2_decap_4
XFILLER_31_1013 VPWR VGND sg13g2_decap_8
XFILLER_7_962 VPWR VGND sg13g2_decap_8
XFILLER_11_991 VPWR VGND sg13g2_decap_8
X_5210_ VGND VPWR net1463 _1180_ _1183_ _1182_ sg13g2_a21oi_1
X_6190_ _2071_ net1741 _2072_ VPWR VGND _2011_ sg13g2_nand3b_1
X_5141_ s0.data_out\[20\]\[5\] s0.data_out\[19\]\[5\] net1464 _1126_ VPWR VGND sg13g2_mux2_1
X_5072_ _1060_ _1059_ _1058_ VPWR VGND sg13g2_nand2b_1
X_4023_ VPWR _3399_ net515 VGND sg13g2_inv_1
XFILLER_49_192 VPWR VGND sg13g2_fill_2
XFILLER_49_181 VPWR VGND sg13g2_fill_2
X_7713_ net311 VGND VPWR net539 s0.data_out\[21\]\[7\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_5974_ VGND VPWR net1378 _1873_ _1875_ _1874_ sg13g2_a21oi_1
X_4925_ _0928_ VPWR _0929_ VGND net1734 net411 sg13g2_o21ai_1
X_7644_ net41 VGND VPWR _0122_ s0.valid_out\[26\][0] clknet_leaf_1_clk sg13g2_dfrbpq_2
X_4856_ _0865_ _0864_ net1690 _0841_ net1699 VPWR VGND sg13g2_a22oi_1
XFILLER_20_221 VPWR VGND sg13g2_fill_2
X_7575_ VGND VPWR net507 _3393_ _3316_ net1640 sg13g2_a21oi_1
XFILLER_21_788 VPWR VGND sg13g2_fill_2
XFILLER_21_799 VPWR VGND sg13g2_fill_1
X_6526_ VGND VPWR net1298 _2370_ _2372_ _2371_ sg13g2_a21oi_1
X_4787_ _0804_ VPWR _0805_ VGND net1182 _0803_ sg13g2_o21ai_1
X_7890__120 VPWR VGND net120 sg13g2_tiehi
X_6457_ net1610 _2242_ _2307_ VPWR VGND sg13g2_nor2_1
X_6388_ net1312 net1335 _2246_ VPWR VGND sg13g2_nor2b_1
X_5408_ _1366_ VPWR _1367_ VGND net1203 _1365_ sg13g2_o21ai_1
X_5339_ s0.data_out\[18\]\[0\] s0.data_out\[17\]\[0\] net1443 _1300_ VPWR VGND sg13g2_mux2_1
XFILLER_0_659 VPWR VGND sg13g2_fill_1
X_7009_ VGND VPWR _2696_ _2806_ _2807_ net1258 sg13g2_a21oi_1
XFILLER_44_869 VPWR VGND sg13g2_decap_8
XFILLER_11_221 VPWR VGND sg13g2_fill_2
XFILLER_11_232 VPWR VGND sg13g2_fill_1
XFILLER_34_97 VPWR VGND sg13g2_fill_1
XFILLER_4_976 VPWR VGND sg13g2_decap_8
Xfanout1210 net1213 net1210 VPWR VGND sg13g2_buf_8
Xfanout1221 net1222 net1221 VPWR VGND sg13g2_buf_2
Xfanout1232 net1233 net1232 VPWR VGND sg13g2_buf_8
Xfanout1254 net1257 net1254 VPWR VGND sg13g2_buf_1
Xfanout1243 net1244 net1243 VPWR VGND sg13g2_buf_8
Xfanout1265 net480 net1265 VPWR VGND sg13g2_buf_8
Xfanout1298 net1299 net1298 VPWR VGND sg13g2_buf_8
Xfanout1287 net1288 net1287 VPWR VGND sg13g2_buf_1
Xfanout1276 net1277 net1276 VPWR VGND sg13g2_buf_8
X_7867__144 VPWR VGND net144 sg13g2_tiehi
XFILLER_47_696 VPWR VGND sg13g2_decap_8
XFILLER_34_302 VPWR VGND sg13g2_fill_2
XFILLER_43_891 VPWR VGND sg13g2_decap_8
X_4710_ VPWR VGND _0730_ net1711 _0726_ net1705 _0731_ _0724_ sg13g2_a221oi_1
X_5690_ _0252_ _1617_ _1618_ _3466_ net1630 VPWR VGND sg13g2_a22oi_1
X_4641_ _0674_ _0673_ net1671 _0667_ net1679 VPWR VGND sg13g2_a22oi_1
XFILLER_30_574 VPWR VGND sg13g2_decap_4
X_4572_ VGND VPWR _0608_ _0607_ _0605_ sg13g2_or2_1
X_7360_ VGND VPWR net1217 _3120_ _3122_ _3121_ sg13g2_a21oi_1
X_6311_ net1369 VPWR _2181_ VGND _2121_ _2180_ sg13g2_o21ai_1
X_7874__137 VPWR VGND net137 sg13g2_tiehi
X_7291_ _2986_ VPWR _3065_ VGND _3039_ _3040_ sg13g2_o21ai_1
X_6242_ _2119_ net1362 net720 VPWR VGND sg13g2_nand2_1
XFILLER_6_291 VPWR VGND sg13g2_fill_1
XFILLER_41_0 VPWR VGND sg13g2_fill_2
X_6173_ net1611 _1979_ _2059_ VPWR VGND sg13g2_nor2_1
X_5124_ net1460 net1331 _1109_ VPWR VGND sg13g2_nor2b_1
X_5055_ VPWR _0188_ _1047_ VGND sg13g2_inv_1
X_4006_ VPWR _3382_ net1395 VGND sg13g2_inv_1
XFILLER_25_357 VPWR VGND sg13g2_fill_2
X_5957_ _1858_ net1386 net789 VPWR VGND sg13g2_nand2_1
XFILLER_40_349 VPWR VGND sg13g2_fill_1
X_4908_ VPWR _0173_ _0915_ VGND sg13g2_inv_1
X_7627_ net404 _3319_ net1721 _0106_ VPWR VGND sg13g2_mux2_1
X_5888_ _1691_ VPWR _1801_ VGND net1409 _3484_ sg13g2_o21ai_1
X_4839_ VGND VPWR _0718_ _0847_ _0848_ net1502 sg13g2_a21oi_1
X_7558_ _3302_ VPWR _3303_ VGND net1722 net714 sg13g2_o21ai_1
X_7489_ VGND VPWR net1211 _3237_ _3239_ _3238_ sg13g2_a21oi_1
X_6509_ _2355_ s0.data_out\[8\]\[7\] net1316 VPWR VGND sg13g2_nand2b_1
XFILLER_49_906 VPWR VGND sg13g2_decap_8
XFILLER_1_957 VPWR VGND sg13g2_decap_8
Xhold20 s0.genblk1\[21\].modules.bubble VPWR VGND net389 sg13g2_dlygate4sd3_1
Xhold31 s0.was_valid_out\[4\][0] VPWR VGND net400 sg13g2_dlygate4sd3_1
Xhold64 s0.data_out\[0\]\[3\] VPWR VGND net433 sg13g2_dlygate4sd3_1
Xhold42 s0.data_out\[22\]\[4\] VPWR VGND net411 sg13g2_dlygate4sd3_1
Xhold53 _0072_ VPWR VGND net422 sg13g2_dlygate4sd3_1
Xhold86 s0.was_valid_out\[9\][0] VPWR VGND net455 sg13g2_dlygate4sd3_1
XFILLER_21_1012 VPWR VGND sg13g2_decap_8
Xhold97 s0.data_out\[16\]\[3\] VPWR VGND net466 sg13g2_dlygate4sd3_1
XFILLER_28_140 VPWR VGND sg13g2_decap_4
XFILLER_29_641 VPWR VGND sg13g2_fill_2
XFILLER_29_663 VPWR VGND sg13g2_fill_2
Xhold75 _2115_ VPWR VGND net444 sg13g2_dlygate4sd3_1
XFILLER_16_302 VPWR VGND sg13g2_fill_2
XFILLER_31_305 VPWR VGND sg13g2_fill_1
XFILLER_32_839 VPWR VGND sg13g2_fill_1
XFILLER_43_198 VPWR VGND sg13g2_fill_1
XFILLER_4_762 VPWR VGND sg13g2_fill_2
XFILLER_39_427 VPWR VGND sg13g2_fill_2
XFILLER_13_4 VPWR VGND sg13g2_fill_2
X_6860_ net1261 net1349 _2670_ VPWR VGND sg13g2_nor2b_1
X_7880__130 VPWR VGND net130 sg13g2_tiehi
X_6791_ _2592_ _2608_ _2611_ _2612_ _2613_ VPWR VGND sg13g2_and4_1
X_5811_ VPWR _0262_ _1729_ VGND sg13g2_inv_1
XFILLER_35_699 VPWR VGND sg13g2_fill_2
X_5742_ _1667_ s0.data_out\[14\]\[7\] net1420 VPWR VGND sg13g2_nand2b_1
X_5673_ _0248_ _1604_ _1605_ _3469_ net1622 VPWR VGND sg13g2_a22oi_1
XFILLER_30_371 VPWR VGND sg13g2_decap_4
X_4624_ VGND VPWR net1523 _0654_ _0657_ _0656_ sg13g2_a21oi_1
X_7412_ _3161_ _3162_ _3171_ _3173_ _3174_ VPWR VGND sg13g2_nor4_1
X_4555_ _0593_ VPWR _0594_ VGND net1184 _0592_ sg13g2_o21ai_1
X_7343_ net1714 net380 _0074_ VPWR VGND sg13g2_and2_1
X_4486_ s0.data_out\[25\]\[7\] s0.data_out\[24\]\[7\] net1528 _0531_ VPWR VGND sg13g2_mux2_1
X_7274_ VGND VPWR net440 _3045_ _3048_ _3047_ sg13g2_a21oi_1
X_6225_ s0.data_out\[11\]\[0\] s0.data_out\[10\]\[0\] net1361 _2102_ VPWR VGND sg13g2_mux2_1
XFILLER_44_1023 VPWR VGND sg13g2_decap_4
X_6156_ _2031_ VPWR _2045_ VGND _2041_ _2042_ sg13g2_o21ai_1
X_5107_ _1091_ VPWR _1092_ VGND net1465 _3448_ sg13g2_o21ai_1
XFILLER_39_950 VPWR VGND sg13g2_decap_8
X_6087_ net1367 net1350 _1976_ VPWR VGND sg13g2_nor2b_1
X_5038_ VGND VPWR net1178 _0962_ _1034_ net1616 sg13g2_a21oi_1
XFILLER_41_614 VPWR VGND sg13g2_fill_1
XFILLER_41_636 VPWR VGND sg13g2_fill_2
XFILLER_40_124 VPWR VGND sg13g2_fill_1
X_6989_ VGND VPWR net1250 _2785_ _2787_ _2786_ sg13g2_a21oi_1
XFILLER_41_669 VPWR VGND sg13g2_fill_1
Xoutput10 net10 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput8 net8 uo_out[5] VPWR VGND sg13g2_buf_1
X_7657__27 VPWR VGND net27 sg13g2_tiehi
XFILLER_0_220 VPWR VGND sg13g2_decap_8
XFILLER_1_754 VPWR VGND sg13g2_decap_8
XFILLER_49_703 VPWR VGND sg13g2_decap_8
XFILLER_37_909 VPWR VGND sg13g2_fill_1
XFILLER_45_942 VPWR VGND sg13g2_decap_8
XFILLER_17_644 VPWR VGND sg13g2_fill_1
XFILLER_17_677 VPWR VGND sg13g2_fill_2
XFILLER_16_198 VPWR VGND sg13g2_fill_2
XFILLER_31_168 VPWR VGND sg13g2_fill_2
XFILLER_8_331 VPWR VGND sg13g2_fill_2
X_7725__298 VPWR VGND net298 sg13g2_tiehi
X_4340_ _0397_ s0.data_out\[25\]\[1\] net1557 VPWR VGND sg13g2_nand2b_1
X_4271_ VGND VPWR _3635_ _3624_ net1668 sg13g2_or2_1
X_6010_ _1911_ net1387 net723 VPWR VGND sg13g2_nand2_1
X_7961_ net230 VGND VPWR _0095_ s0.data_out\[1\]\[7\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_6912_ _2719_ _2721_ net1679 _2722_ VPWR VGND sg13g2_nand3_1
X_7892_ net117 VGND VPWR _0026_ s0.genblk1\[5\].modules.bubble clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_36_986 VPWR VGND sg13g2_decap_8
X_6843_ net1727 net378 _0026_ VPWR VGND sg13g2_and2_1
X_6774_ VGND VPWR net1276 _2595_ _2596_ _2593_ sg13g2_a21oi_1
XFILLER_22_135 VPWR VGND sg13g2_fill_1
X_3986_ VPWR _3362_ net423 VGND sg13g2_inv_1
X_5725_ _1650_ net1573 _1648_ VPWR VGND sg13g2_xnor2_1
X_5656_ VGND VPWR _1588_ _1591_ _0244_ _1592_ sg13g2_a21oi_1
X_4607_ _0640_ s0.data_out\[23\]\[3\] net1531 VPWR VGND sg13g2_nand2b_1
Xhold320 s0.data_out\[17\]\[0\] VPWR VGND net689 sg13g2_dlygate4sd3_1
X_5587_ VGND VPWR net1424 _1521_ _1524_ _1523_ sg13g2_a21oi_1
Xhold331 s0.data_out\[18\]\[5\] VPWR VGND net700 sg13g2_dlygate4sd3_1
X_4538_ _0138_ _0579_ _0580_ _3421_ net1581 VPWR VGND sg13g2_a22oi_1
X_7326_ VPWR _0070_ _3092_ VGND sg13g2_inv_1
Xhold342 s0.data_out\[22\]\[2\] VPWR VGND net711 sg13g2_dlygate4sd3_1
Xhold353 _3180_ VPWR VGND net722 sg13g2_dlygate4sd3_1
Xhold364 s0.data_out\[1\]\[5\] VPWR VGND net733 sg13g2_dlygate4sd3_1
Xhold386 s0.data_out\[22\]\[5\] VPWR VGND net755 sg13g2_dlygate4sd3_1
X_4469_ _0514_ net1185 _0513_ VPWR VGND sg13g2_nand2_1
Xhold375 s0.data_out\[3\]\[2\] VPWR VGND net744 sg13g2_dlygate4sd3_1
X_7257_ _3028_ _3030_ _3031_ VPWR VGND sg13g2_and2_1
X_6208_ net1613 _2080_ _0302_ VPWR VGND sg13g2_nor2_1
Xhold397 _0260_ VPWR VGND net766 sg13g2_dlygate4sd3_1
X_7188_ VGND VPWR net1244 net616 _2969_ _2920_ sg13g2_a21oi_1
X_6139_ _2028_ net639 net1387 VPWR VGND sg13g2_nand2b_1
XFILLER_45_238 VPWR VGND sg13g2_fill_2
XFILLER_26_32 VPWR VGND sg13g2_fill_1
XFILLER_27_942 VPWR VGND sg13g2_fill_2
XFILLER_42_989 VPWR VGND sg13g2_decap_8
XFILLER_10_820 VPWR VGND sg13g2_decap_8
XFILLER_42_75 VPWR VGND sg13g2_fill_1
XFILLER_42_97 VPWR VGND sg13g2_fill_2
X_7679__348 VPWR VGND net348 sg13g2_tiehi
XFILLER_49_500 VPWR VGND sg13g2_fill_2
XFILLER_49_577 VPWR VGND sg13g2_decap_8
X_7731__291 VPWR VGND net291 sg13g2_tiehi
XFILLER_45_750 VPWR VGND sg13g2_decap_8
XFILLER_17_452 VPWR VGND sg13g2_fill_1
XFILLER_44_271 VPWR VGND sg13g2_fill_2
XFILLER_33_967 VPWR VGND sg13g2_decap_8
X_5510_ _1459_ _3375_ _1458_ VPWR VGND sg13g2_nand2_1
X_6490_ VGND VPWR net1295 _2334_ _2336_ _2335_ sg13g2_a21oi_1
X_5441_ _1391_ _1392_ _1393_ VPWR VGND sg13g2_nor2_1
X_5372_ net1666 _1324_ _1333_ VPWR VGND sg13g2_nor2_1
X_4323_ _0380_ VPWR _0383_ VGND net1549 _0382_ sg13g2_o21ai_1
X_7111_ net1570 _2896_ _2897_ VPWR VGND sg13g2_and2_1
X_7042_ _2765_ VPWR _2840_ VGND _2816_ _2818_ sg13g2_o21ai_1
X_4254_ net1564 s0.data_out\[26\]\[5\] _3618_ VPWR VGND sg13g2_nor2_1
X_4185_ net1724 net382 _0108_ VPWR VGND sg13g2_and2_1
X_7644__41 VPWR VGND net41 sg13g2_tiehi
X_7944_ net61 VGND VPWR _0078_ s0.data_out\[2\]\[2\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_7875_ net136 VGND VPWR _0009_ s0.data_out\[8\]\[5\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_6826_ _2640_ net1729 _2641_ VPWR VGND _2587_ sg13g2_nand3b_1
X_6757_ _2579_ s0.data_out\[6\]\[7\] net1291 VPWR VGND sg13g2_nand2b_1
X_5708_ VGND VPWR _1526_ _1632_ _1633_ net1412 sg13g2_a21oi_1
X_6688_ net1177 _3515_ _2518_ VPWR VGND sg13g2_nor2_1
X_5639_ s0.data_out\[16\]\[5\] s0.data_out\[15\]\[5\] net1421 _1576_ VPWR VGND sg13g2_mux2_1
XFILLER_3_805 VPWR VGND sg13g2_decap_8
Xhold150 _2750_ VPWR VGND net519 sg13g2_dlygate4sd3_1
XFILLER_2_348 VPWR VGND sg13g2_fill_2
Xhold161 s0.data_out\[22\]\[3\] VPWR VGND net530 sg13g2_dlygate4sd3_1
X_7309_ VPWR _0066_ net745 VGND sg13g2_inv_1
Xhold172 _0300_ VPWR VGND net541 sg13g2_dlygate4sd3_1
Xfanout1606 net1607 net1606 VPWR VGND sg13g2_buf_8
Xhold183 s0.data_out\[22\]\[6\] VPWR VGND net552 sg13g2_dlygate4sd3_1
Xhold194 s0.data_out\[20\]\[4\] VPWR VGND net563 sg13g2_dlygate4sd3_1
Xfanout1639 net1642 net1639 VPWR VGND sg13g2_buf_8
Xfanout1617 net1621 net1617 VPWR VGND sg13g2_buf_8
Xfanout1628 net1631 net1628 VPWR VGND sg13g2_buf_8
X_7685__341 VPWR VGND net341 sg13g2_tiehi
XFILLER_42_764 VPWR VGND sg13g2_fill_1
XFILLER_15_989 VPWR VGND sg13g2_decap_8
XFILLER_30_948 VPWR VGND sg13g2_fill_2
XFILLER_5_164 VPWR VGND sg13g2_fill_2
XFILLER_2_882 VPWR VGND sg13g2_decap_8
X_5990_ _1889_ _1890_ _1891_ VPWR VGND _1881_ sg13g2_nand3b_1
X_4941_ net1643 _3392_ _0941_ VPWR VGND sg13g2_nor2_1
XFILLER_33_720 VPWR VGND sg13g2_fill_2
X_4872_ _0881_ _0880_ net1663 _0873_ net1653 VPWR VGND sg13g2_a22oi_1
X_7660_ net24 VGND VPWR net708 s0.data_out\[25\]\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_6611_ net1283 net1355 _2445_ VPWR VGND sg13g2_nor2b_1
X_7591_ _3328_ VPWR _3329_ VGND _3393_ net1353 sg13g2_o21ai_1
X_6542_ VGND VPWR _2373_ _2375_ _2388_ net1670 sg13g2_a21oi_1
XFILLER_9_470 VPWR VGND sg13g2_fill_1
X_6473_ _2319_ net1301 net674 VPWR VGND sg13g2_nand2_1
X_5424_ net1439 s0.data_out\[17\]\[5\] _1379_ VPWR VGND sg13g2_and2_1
X_5355_ _1316_ net1693 _1315_ VPWR VGND sg13g2_nand2_1
X_4306_ _0118_ _0367_ _0368_ _3405_ net1575 VPWR VGND sg13g2_a22oi_1
X_5286_ net1619 _1190_ _1257_ VPWR VGND sg13g2_nor2_1
X_4237_ s0.data_out\[27\]\[7\] s0.data_out\[26\]\[7\] net1554 _3601_ VPWR VGND sg13g2_mux2_1
X_7025_ _2823_ s0.data_out\[4\]\[4\] net1268 VPWR VGND sg13g2_nand2b_1
X_4168_ s0.was_valid_out\[27\][0] net1560 _3544_ VPWR VGND sg13g2_nor2_2
XFILLER_28_558 VPWR VGND sg13g2_fill_2
X_4099_ VPWR _3475_ net702 VGND sg13g2_inv_1
X_7669__358 VPWR VGND net358 sg13g2_tiehi
XFILLER_15_219 VPWR VGND sg13g2_fill_2
X_7927_ net79 VGND VPWR _0061_ s0.valid_out\[3\][0] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_7858_ net154 VGND VPWR _0336_ s0.data_out\[9\]\[0\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_6809_ _0018_ _2626_ _2627_ _3516_ net1598 VPWR VGND sg13g2_a22oi_1
X_7789_ net228 VGND VPWR _0267_ s0.genblk1\[13\].modules.bubble clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
XFILLER_11_447 VPWR VGND sg13g2_fill_2
XFILLER_7_418 VPWR VGND sg13g2_fill_1
XFILLER_20_970 VPWR VGND sg13g2_decap_8
XFILLER_23_88 VPWR VGND sg13g2_decap_4
XFILLER_23_99 VPWR VGND sg13g2_fill_1
Xfanout1414 net468 net1414 VPWR VGND sg13g2_buf_2
Xfanout1403 net474 net1403 VPWR VGND sg13g2_buf_2
Xfanout1447 net1448 net1447 VPWR VGND sg13g2_buf_8
Xfanout1436 net1437 net1436 VPWR VGND sg13g2_buf_8
Xfanout1425 net1431 net1425 VPWR VGND sg13g2_buf_8
XFILLER_24_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_801 VPWR VGND sg13g2_decap_8
Xfanout1469 net1477 net1469 VPWR VGND sg13g2_buf_2
Xfanout1458 net1460 net1458 VPWR VGND sg13g2_buf_2
XFILLER_47_878 VPWR VGND sg13g2_decap_8
XFILLER_46_355 VPWR VGND sg13g2_fill_1
XFILLER_14_252 VPWR VGND sg13g2_fill_1
XFILLER_30_778 VPWR VGND sg13g2_fill_1
XFILLER_7_941 VPWR VGND sg13g2_decap_8
X_7954__321 VPWR VGND net321 sg13g2_tiehi
X_5140_ _1125_ net1466 s0.data_out\[19\]\[5\] VPWR VGND sg13g2_nand2_1
X_5071_ _1059_ net1635 net1464 VPWR VGND sg13g2_nand2_1
X_4022_ VPWR _3398_ net557 VGND sg13g2_inv_1
XFILLER_25_506 VPWR VGND sg13g2_decap_4
X_5973_ net1378 net1359 _1874_ VPWR VGND sg13g2_nor2b_1
X_7712_ net312 VGND VPWR _0190_ s0.data_out\[21\]\[6\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_4924_ _0900_ _0927_ net1734 _0928_ VPWR VGND sg13g2_nand3_1
X_7643_ net43 VGND VPWR _0121_ s0.was_valid_out\[26\][0] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4855_ VGND VPWR net1500 _0861_ _0864_ _0863_ sg13g2_a21oi_1
X_7574_ VPWR _0095_ net728 VGND sg13g2_inv_1
X_4786_ VGND VPWR net1183 _0736_ _0804_ net1595 sg13g2_a21oi_1
XFILLER_20_255 VPWR VGND sg13g2_decap_4
X_6525_ net1296 net1339 _2371_ VPWR VGND sg13g2_nor2b_1
X_6456_ net1323 VPWR _2306_ VGND _2239_ _2305_ sg13g2_o21ai_1
X_6387_ s0.data_out\[10\]\[6\] s0.data_out\[9\]\[6\] net1317 _2245_ VPWR VGND sg13g2_mux2_1
X_5407_ VGND VPWR net1203 _1297_ _1366_ net1619 sg13g2_a21oi_1
XFILLER_0_638 VPWR VGND sg13g2_decap_8
X_5338_ _1296_ _1298_ net1708 _1299_ VPWR VGND sg13g2_nand3_1
X_5269_ _1242_ net1683 _1241_ VPWR VGND sg13g2_nand2_1
X_7008_ _2806_ s0.data_out\[4\]\[7\] net1267 VPWR VGND sg13g2_nand2b_1
XFILLER_18_11 VPWR VGND sg13g2_decap_8
XFILLER_18_22 VPWR VGND sg13g2_fill_1
XFILLER_29_845 VPWR VGND sg13g2_fill_2
XFILLER_44_848 VPWR VGND sg13g2_decap_8
XFILLER_43_336 VPWR VGND sg13g2_fill_2
X_7682__344 VPWR VGND net344 sg13g2_tiehi
XFILLER_34_87 VPWR VGND sg13g2_fill_1
XFILLER_8_727 VPWR VGND sg13g2_decap_8
XFILLER_12_767 VPWR VGND sg13g2_fill_2
XFILLER_4_955 VPWR VGND sg13g2_decap_8
Xfanout1211 net1212 net1211 VPWR VGND sg13g2_buf_2
Xfanout1200 net1201 net1200 VPWR VGND sg13g2_buf_8
Xfanout1222 net1223 net1222 VPWR VGND sg13g2_buf_1
Xfanout1255 net1257 net1255 VPWR VGND sg13g2_buf_8
Xfanout1244 net440 net1244 VPWR VGND sg13g2_buf_2
Xfanout1233 net1234 net1233 VPWR VGND sg13g2_buf_8
XFILLER_47_620 VPWR VGND sg13g2_fill_2
Xfanout1299 net1300 net1299 VPWR VGND sg13g2_buf_2
Xfanout1288 s0.shift_out\[7\][0] net1288 VPWR VGND sg13g2_buf_2
Xfanout1277 net445 net1277 VPWR VGND sg13g2_buf_1
Xfanout1266 net1267 net1266 VPWR VGND sg13g2_buf_8
XFILLER_47_675 VPWR VGND sg13g2_decap_8
XFILLER_46_196 VPWR VGND sg13g2_fill_1
X_4640_ VGND VPWR net1524 _0670_ _0673_ _0672_ sg13g2_a21oi_1
X_6310_ net1325 s0.data_out\[10\]\[6\] _2180_ VPWR VGND sg13g2_and2_1
X_4571_ net409 net1515 _0607_ VPWR VGND sg13g2_nor2_1
X_7290_ _3049_ _3059_ _3064_ VPWR VGND sg13g2_nor2_1
X_6241_ _2117_ VPWR _2118_ VGND _2108_ _2109_ sg13g2_o21ai_1
X_6172_ net1376 VPWR _2058_ VGND _1976_ _2057_ sg13g2_o21ai_1
X_5123_ s0.data_out\[20\]\[7\] s0.data_out\[19\]\[7\] net1464 _1108_ VPWR VGND sg13g2_mux2_1
XFILLER_34_0 VPWR VGND sg13g2_fill_2
X_5054_ _1046_ VPWR _1047_ VGND net1736 net680 sg13g2_o21ai_1
X_4005_ _3381_ net1404 VPWR VGND sg13g2_inv_2
XFILLER_34_870 VPWR VGND sg13g2_fill_1
X_5956_ net1750 net377 _0279_ VPWR VGND sg13g2_and2_1
X_4907_ _0914_ VPWR _0915_ VGND net1735 net759 sg13g2_o21ai_1
X_5887_ VGND VPWR net1394 _1798_ _1800_ _1799_ sg13g2_a21oi_1
X_7626_ VGND VPWR net1722 _3326_ _0105_ _3357_ sg13g2_a21oi_1
X_4838_ _0847_ s0.data_out\[21\]\[1\] net1506 VPWR VGND sg13g2_nand2b_1
X_7557_ _3301_ VPWR _3302_ VGND net1200 _3300_ sg13g2_o21ai_1
X_4769_ _0770_ _0786_ _0787_ _0788_ _0790_ VPWR VGND sg13g2_nor4_1
X_7488_ net1211 net1347 _3238_ VPWR VGND sg13g2_nor2b_1
X_6508_ _2352_ net1298 _2353_ _2354_ VPWR VGND sg13g2_a21o_1
X_6439_ net1609 _2233_ _2293_ VPWR VGND sg13g2_nor2_1
XFILLER_1_936 VPWR VGND sg13g2_decap_8
XFILLER_0_424 VPWR VGND sg13g2_decap_4
Xhold21 s0.genblk1\[11\].modules.bubble VPWR VGND net390 sg13g2_dlygate4sd3_1
Xhold10 s0.genblk1\[25\].modules.bubble VPWR VGND net379 sg13g2_dlygate4sd3_1
Xhold32 _0048_ VPWR VGND net401 sg13g2_dlygate4sd3_1
Xhold65 s0.data_out\[0\]\[4\] VPWR VGND net434 sg13g2_dlygate4sd3_1
Xhold43 s0.was_valid_out\[21\][0] VPWR VGND net412 sg13g2_dlygate4sd3_1
Xhold54 s0.was_valid_out\[5\][0] VPWR VGND net423 sg13g2_dlygate4sd3_1
Xhold87 _0332_ VPWR VGND net456 sg13g2_dlygate4sd3_1
Xhold76 s0.shift_out\[6\][0] VPWR VGND net445 sg13g2_dlygate4sd3_1
Xhold98 _0248_ VPWR VGND net467 sg13g2_dlygate4sd3_1
XFILLER_28_152 VPWR VGND sg13g2_fill_2
XFILLER_44_645 VPWR VGND sg13g2_decap_8
XFILLER_31_317 VPWR VGND sg13g2_fill_1
XFILLER_8_557 VPWR VGND sg13g2_fill_2
XFILLER_48_984 VPWR VGND sg13g2_decap_8
X_6790_ _2612_ net1680 _2599_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_829 VPWR VGND sg13g2_decap_8
X_5810_ _1728_ VPWR _1729_ VGND net1748 net644 sg13g2_o21ai_1
X_5741_ _1664_ net1405 _1665_ _1666_ VPWR VGND sg13g2_a21o_1
XFILLER_31_873 VPWR VGND sg13g2_fill_1
X_5672_ net1622 _1547_ _1605_ VPWR VGND sg13g2_nor2_1
X_7411_ _3172_ VPWR _3173_ VGND net1686 _3136_ sg13g2_o21ai_1
X_4623_ VGND VPWR _0537_ _0655_ _0656_ net1523 sg13g2_a21oi_1
X_4554_ VGND VPWR net1184 _0554_ _0593_ net1589 sg13g2_a21oi_1
X_7342_ net1582 _3098_ _3099_ _0073_ VPWR VGND sg13g2_nor3_1
X_7273_ VGND VPWR _2909_ _3046_ _3047_ net1243 sg13g2_a21oi_1
X_4485_ _0530_ net1530 net525 VPWR VGND sg13g2_nand2_1
X_6224_ VGND VPWR net1365 _2098_ _2101_ _2100_ sg13g2_a21oi_1
XFILLER_44_1002 VPWR VGND sg13g2_decap_8
X_6155_ _2040_ _2041_ _2005_ _2044_ VPWR VGND _2043_ sg13g2_nand4_1
X_5106_ _1091_ net1465 net814 VPWR VGND sg13g2_nand2_1
X_6086_ s0.data_out\[12\]\[2\] s0.data_out\[11\]\[2\] net1373 _1975_ VPWR VGND sg13g2_mux2_1
X_5037_ VGND VPWR net1471 net497 _1033_ _0957_ sg13g2_a21oi_1
XFILLER_38_483 VPWR VGND sg13g2_fill_2
XFILLER_13_306 VPWR VGND sg13g2_fill_1
X_6988_ net1250 net1357 _2786_ VPWR VGND sg13g2_nor2b_1
X_5939_ VPWR _0275_ net697 VGND sg13g2_inv_1
X_7609_ _3347_ _3343_ net1678 _3326_ net1669 VPWR VGND sg13g2_a22oi_1
XFILLER_5_527 VPWR VGND sg13g2_fill_1
X_7857__155 VPWR VGND net155 sg13g2_tiehi
Xoutput9 net9 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_1_711 VPWR VGND sg13g2_decap_4
XFILLER_1_733 VPWR VGND sg13g2_decap_8
XFILLER_49_759 VPWR VGND sg13g2_decap_8
XFILLER_0_265 VPWR VGND sg13g2_fill_2
XFILLER_45_921 VPWR VGND sg13g2_decap_8
XFILLER_17_623 VPWR VGND sg13g2_decap_4
X_7864__148 VPWR VGND net148 sg13g2_tiehi
XFILLER_45_998 VPWR VGND sg13g2_decap_8
XFILLER_13_862 VPWR VGND sg13g2_fill_1
X_4270_ net1677 _3633_ _3634_ VPWR VGND sg13g2_and2_1
XFILLER_48_781 VPWR VGND sg13g2_decap_8
X_7960_ net243 VGND VPWR _0094_ s0.data_out\[1\]\[6\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_7891_ net118 VGND VPWR _0025_ s0.valid_out\[6\][0] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_6911_ _2721_ net1174 _2720_ VPWR VGND sg13g2_nand2_1
XFILLER_36_965 VPWR VGND sg13g2_decap_8
XFILLER_36_943 VPWR VGND sg13g2_decap_4
X_6842_ net1729 _2648_ _0025_ VPWR VGND sg13g2_and2_1
X_6773_ _2594_ VPWR _2595_ VGND net1281 _3518_ sg13g2_o21ai_1
X_3985_ VPWR _3361_ net400 VGND sg13g2_inv_1
XFILLER_22_169 VPWR VGND sg13g2_decap_8
X_5724_ VGND VPWR _1649_ _1648_ net1573 sg13g2_or2_1
X_5655_ VGND VPWR _1592_ net1567 net391 sg13g2_or2_1
XFILLER_11_1012 VPWR VGND sg13g2_decap_8
X_4606_ _0637_ net1510 _0638_ _0639_ VPWR VGND sg13g2_a21o_1
X_5586_ VGND VPWR _1413_ _1522_ _1523_ net1425 sg13g2_a21oi_1
X_7325_ _3091_ VPWR _3092_ VGND net1714 net812 sg13g2_o21ai_1
Xhold310 s0.data_out\[15\]\[0\] VPWR VGND net679 sg13g2_dlygate4sd3_1
Xhold343 s0.data_out\[7\]\[5\] VPWR VGND net712 sg13g2_dlygate4sd3_1
Xhold332 _0226_ VPWR VGND net701 sg13g2_dlygate4sd3_1
X_4537_ net1580 _0499_ _0580_ VPWR VGND sg13g2_nor2_1
Xhold321 _1482_ VPWR VGND net690 sg13g2_dlygate4sd3_1
Xhold365 _3307_ VPWR VGND net734 sg13g2_dlygate4sd3_1
Xhold354 s0.data_out\[12\]\[6\] VPWR VGND net723 sg13g2_dlygate4sd3_1
Xhold387 s0.data_out\[2\]\[2\] VPWR VGND net756 sg13g2_dlygate4sd3_1
X_4468_ _0385_ VPWR _0513_ VGND net1543 _3430_ sg13g2_o21ai_1
Xhold376 _3079_ VPWR VGND net745 sg13g2_dlygate4sd3_1
X_7256_ _3030_ net1190 _3029_ VPWR VGND sg13g2_nand2_1
X_6207_ _2081_ _2086_ _0301_ VPWR VGND sg13g2_nor2_1
Xhold398 s0.data_out\[18\]\[6\] VPWR VGND net767 sg13g2_dlygate4sd3_1
X_7187_ _0055_ _2967_ _2968_ _3533_ net1586 VPWR VGND sg13g2_a22oi_1
X_6138_ _2025_ net1370 _2026_ _2027_ VPWR VGND sg13g2_a21o_1
X_4399_ _0435_ _0450_ _0456_ VPWR VGND sg13g2_nor2_1
X_6069_ net1629 _1923_ _1962_ VPWR VGND sg13g2_nor2_1
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_42_968 VPWR VGND sg13g2_decap_8
XFILLER_13_125 VPWR VGND sg13g2_fill_1
XFILLER_14_659 VPWR VGND sg13g2_fill_2
X_7870__141 VPWR VGND net141 sg13g2_tiehi
XFILLER_49_556 VPWR VGND sg13g2_decap_8
XFILLER_29_280 VPWR VGND sg13g2_fill_1
XFILLER_33_924 VPWR VGND sg13g2_fill_2
XFILLER_20_629 VPWR VGND sg13g2_decap_4
XFILLER_34_1012 VPWR VGND sg13g2_decap_8
X_5440_ VGND VPWR net1635 net1445 _1392_ net1440 sg13g2_a21oi_1
X_5371_ _1332_ _1331_ net1654 _1324_ net1664 VPWR VGND sg13g2_a22oi_1
X_4322_ net419 net1556 _0382_ VPWR VGND sg13g2_nor2_1
X_7110_ _2895_ VPWR _2896_ VGND net1170 _2893_ sg13g2_o21ai_1
X_4253_ net461 net1563 _3617_ VPWR VGND sg13g2_nor2b_1
X_7041_ _2819_ _2833_ _2835_ _2839_ VPWR VGND sg13g2_nor3_1
X_4184_ _3552_ VPWR net10 VGND _3399_ net1165 sg13g2_o21ai_1
X_7943_ net62 VGND VPWR _0077_ s0.data_out\[2\]\[1\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_7874_ net137 VGND VPWR _0008_ s0.data_out\[8\]\[4\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_6825_ net1285 VPWR _2640_ VGND _2584_ _2639_ sg13g2_o21ai_1
XFILLER_24_979 VPWR VGND sg13g2_decap_8
X_6756_ _2576_ net1276 _2577_ _2578_ VPWR VGND sg13g2_a21o_1
X_5707_ _1632_ net603 net1419 VPWR VGND sg13g2_nand2b_1
X_6687_ _0006_ _2516_ _2517_ _3512_ net1599 VPWR VGND sg13g2_a22oi_1
X_5638_ _1575_ net1420 s0.data_out\[15\]\[5\] VPWR VGND sg13g2_nand2_1
X_5569_ _1509_ net1635 net1421 VPWR VGND sg13g2_nand2_1
Xhold151 s0.data_out\[2\]\[4\] VPWR VGND net520 sg13g2_dlygate4sd3_1
Xhold140 s0.data_out\[20\]\[5\] VPWR VGND net509 sg13g2_dlygate4sd3_1
Xhold162 _0176_ VPWR VGND net531 sg13g2_dlygate4sd3_1
X_7308_ _3078_ VPWR _3079_ VGND net1715 net744 sg13g2_o21ai_1
Xhold184 _0179_ VPWR VGND net553 sg13g2_dlygate4sd3_1
Xhold173 s0.data_out\[17\]\[3\] VPWR VGND net542 sg13g2_dlygate4sd3_1
Xhold195 s0.data_out\[15\]\[7\] VPWR VGND net564 sg13g2_dlygate4sd3_1
Xfanout1629 net1631 net1629 VPWR VGND sg13g2_buf_8
Xfanout1618 net1621 net1618 VPWR VGND sg13g2_buf_1
Xfanout1607 net1616 net1607 VPWR VGND sg13g2_buf_8
X_7239_ _3013_ _3005_ net1570 _2998_ _3415_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_401 VPWR VGND sg13g2_fill_1
XFILLER_15_946 VPWR VGND sg13g2_fill_2
XFILLER_2_861 VPWR VGND sg13g2_decap_8
X_7641__45 VPWR VGND net45 sg13g2_tiehi
X_4940_ net1483 VPWR _0940_ VGND net1643 net1468 sg13g2_o21ai_1
XFILLER_17_261 VPWR VGND sg13g2_fill_1
X_4871_ VGND VPWR net1499 _0877_ _0880_ _0879_ sg13g2_a21oi_1
X_7590_ net430 net1214 net1208 _3328_ VPWR VGND sg13g2_a21o_1
XFILLER_21_927 VPWR VGND sg13g2_fill_1
X_6610_ s0.data_out\[8\]\[1\] s0.data_out\[7\]\[1\] net1289 _2444_ VPWR VGND sg13g2_mux2_1
X_6541_ VGND VPWR _2382_ _2384_ _2387_ net1685 sg13g2_a21oi_1
X_6472_ net1732 net376 _0334_ VPWR VGND sg13g2_and2_1
X_5423_ _0225_ _1377_ _1378_ _3459_ net1624 VPWR VGND sg13g2_a22oi_1
X_5354_ VGND VPWR net1449 _1312_ _1315_ _1314_ sg13g2_a21oi_1
X_4305_ net1576 _3619_ _0368_ VPWR VGND sg13g2_nor2_1
X_5285_ net1459 VPWR _1256_ VGND _1187_ _1255_ sg13g2_o21ai_1
X_4236_ _3600_ net1556 net557 VPWR VGND sg13g2_nand2_1
X_7024_ _2820_ net1252 _2821_ _2822_ VPWR VGND sg13g2_a21o_1
X_4167_ VPWR _3543_ s0.data_out\[0\]\[3\] VGND sg13g2_inv_1
X_4098_ VPWR _3474_ net606 VGND sg13g2_inv_1
X_7926_ net81 VGND VPWR net403 s0.was_valid_out\[3\][0] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_7857_ net155 VGND VPWR _0335_ s0.shift_out\[9\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_23_220 VPWR VGND sg13g2_fill_1
XFILLER_23_231 VPWR VGND sg13g2_fill_1
X_6808_ net1598 _2548_ _2627_ VPWR VGND sg13g2_nor2_1
X_7788_ net229 VGND VPWR _0266_ s0.valid_out\[14\][0] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_6739_ _2561_ net1284 _2560_ VPWR VGND sg13g2_nand2b_1
XFILLER_3_603 VPWR VGND sg13g2_fill_1
Xfanout1404 net1407 net1404 VPWR VGND sg13g2_buf_8
Xfanout1448 net1452 net1448 VPWR VGND sg13g2_buf_8
Xfanout1437 net1438 net1437 VPWR VGND sg13g2_buf_1
Xfanout1426 net1430 net1426 VPWR VGND sg13g2_buf_8
XFILLER_24_1000 VPWR VGND sg13g2_decap_8
Xfanout1415 net1418 net1415 VPWR VGND sg13g2_buf_8
Xfanout1459 net1460 net1459 VPWR VGND sg13g2_buf_1
XFILLER_47_857 VPWR VGND sg13g2_decap_8
XFILLER_9_25 VPWR VGND sg13g2_fill_2
XFILLER_14_264 VPWR VGND sg13g2_fill_1
XFILLER_7_997 VPWR VGND sg13g2_decap_8
XFILLER_9_1016 VPWR VGND sg13g2_decap_8
XFILLER_9_1027 VPWR VGND sg13g2_fill_2
X_5070_ net1474 VPWR _1058_ VGND net1644 net1457 sg13g2_o21ai_1
X_4021_ VPWR _3397_ net1249 VGND sg13g2_inv_1
X_5972_ s0.data_out\[13\]\[0\] s0.data_out\[12\]\[0\] net1388 _1873_ VPWR VGND sg13g2_mux2_1
XFILLER_46_890 VPWR VGND sg13g2_decap_8
X_7711_ net313 VGND VPWR _0189_ s0.data_out\[21\]\[5\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_4923_ net1500 VPWR _0927_ VGND _0894_ _0926_ sg13g2_o21ai_1
X_7642_ net44 VGND VPWR net516 s0.data_out\[27\]\[7\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4854_ VGND VPWR _0742_ _0862_ _0863_ net1502 sg13g2_a21oi_1
X_7573_ _3314_ VPWR _3315_ VGND net1721 net727 sg13g2_o21ai_1
X_4785_ VGND VPWR net1495 s0.data_out\[22\]\[2\] _0803_ _0734_ sg13g2_a21oi_1
X_6524_ s0.data_out\[9\]\[5\] s0.data_out\[8\]\[5\] net1303 _2370_ VPWR VGND sg13g2_mux2_1
X_6455_ net1311 net483 _2305_ VPWR VGND sg13g2_and2_1
XFILLER_47_1011 VPWR VGND sg13g2_decap_8
X_6386_ _2244_ net1316 net731 VPWR VGND sg13g2_nand2_1
X_5406_ VGND VPWR net1436 s0.data_out\[17\]\[1\] _1365_ _1294_ sg13g2_a21oi_1
X_7675__352 VPWR VGND net352 sg13g2_tiehi
XFILLER_0_617 VPWR VGND sg13g2_decap_8
X_5337_ _1298_ net1203 _1297_ VPWR VGND sg13g2_nand2_1
X_5268_ VGND VPWR net1461 _1238_ _1241_ _1240_ sg13g2_a21oi_1
X_4219_ VGND VPWR net1546 _3582_ _3583_ _3580_ sg13g2_a21oi_1
X_7007_ _2803_ net1251 _2804_ _2805_ VPWR VGND sg13g2_a21o_1
X_5199_ VGND VPWR net1198 _1059_ _1175_ _1170_ sg13g2_a21oi_1
XFILLER_44_805 VPWR VGND sg13g2_fill_1
X_7909_ net99 VGND VPWR _0043_ s0.data_out\[5\]\[3\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_4_934 VPWR VGND sg13g2_decap_8
XFILLER_3_444 VPWR VGND sg13g2_fill_2
Xfanout1223 s0.shift_out\[1\][0] net1223 VPWR VGND sg13g2_buf_1
Xfanout1212 net1213 net1212 VPWR VGND sg13g2_buf_8
Xfanout1201 net1202 net1201 VPWR VGND sg13g2_buf_8
Xfanout1245 net1246 net1245 VPWR VGND sg13g2_buf_8
Xfanout1234 s0.shift_out\[2\][0] net1234 VPWR VGND sg13g2_buf_1
Xfanout1256 net1257 net1256 VPWR VGND sg13g2_buf_1
XFILLER_19_323 VPWR VGND sg13g2_fill_2
Xfanout1267 net1269 net1267 VPWR VGND sg13g2_buf_8
Xfanout1278 net1279 net1278 VPWR VGND sg13g2_buf_8
Xfanout1289 net1290 net1289 VPWR VGND sg13g2_buf_8
XFILLER_34_304 VPWR VGND sg13g2_fill_1
XFILLER_42_381 VPWR VGND sg13g2_fill_1
XFILLER_30_510 VPWR VGND sg13g2_fill_2
X_4570_ _0605_ VPWR _0606_ VGND net1523 _0486_ sg13g2_o21ai_1
X_6240_ _2117_ _2116_ net1690 _2093_ net1697 VPWR VGND sg13g2_a22oi_1
X_6171_ _3383_ _3494_ _2057_ VPWR VGND sg13g2_nor2_1
X_5122_ _1107_ net1466 net672 VPWR VGND sg13g2_nand2_1
XFILLER_27_0 VPWR VGND sg13g2_fill_1
X_5053_ _1045_ VPWR _1046_ VGND net1180 _1044_ sg13g2_o21ai_1
X_4004_ _3380_ net1417 VPWR VGND sg13g2_inv_2
XFILLER_26_816 VPWR VGND sg13g2_fill_2
X_5955_ net1628 _1850_ _1851_ _0278_ VPWR VGND sg13g2_nor3_1
XFILLER_40_307 VPWR VGND sg13g2_fill_1
XFILLER_25_359 VPWR VGND sg13g2_fill_1
X_4906_ _0855_ _0913_ net1735 _0914_ VPWR VGND sg13g2_nand3_1
X_5886_ net1394 net1345 _1799_ VPWR VGND sg13g2_nor2b_1
X_7625_ net1723 net439 _3357_ VPWR VGND sg13g2_nor2_1
X_4837_ _0844_ net1487 _0845_ _0846_ VPWR VGND sg13g2_a21o_1
XFILLER_21_576 VPWR VGND sg13g2_decap_8
X_7556_ VGND VPWR net1200 _3268_ _3301_ net1587 sg13g2_a21oi_1
X_4768_ _0777_ _0775_ net1671 _0789_ VPWR VGND sg13g2_a21o_1
X_7487_ s0.data_out\[1\]\[3\] s0.data_out\[0\]\[3\] net1215 _3237_ VPWR VGND sg13g2_mux2_1
X_6507_ net1298 net1329 _2353_ VPWR VGND sg13g2_nor2b_1
X_4699_ net1495 net1355 _0720_ VPWR VGND sg13g2_nor2b_1
X_6438_ net1320 VPWR _2292_ VGND _2230_ _2291_ sg13g2_o21ai_1
XFILLER_1_915 VPWR VGND sg13g2_decap_8
X_6369_ VPWR VGND _2225_ net1711 _2223_ net1705 _2227_ _2219_ sg13g2_a221oi_1
Xhold11 s0.genblk1\[27\].modules.bubble VPWR VGND net380 sg13g2_dlygate4sd3_1
XFILLER_0_458 VPWR VGND sg13g2_fill_2
Xhold22 s0.genblk1\[16\].modules.bubble VPWR VGND net391 sg13g2_dlygate4sd3_1
Xhold55 s0.shift_out\[22\][0] VPWR VGND net424 sg13g2_dlygate4sd3_1
Xhold44 _0181_ VPWR VGND net413 sg13g2_dlygate4sd3_1
Xhold33 s0.was_valid_out\[3\][0] VPWR VGND net402 sg13g2_dlygate4sd3_1
Xhold66 s0.data_out\[19\]\[4\] VPWR VGND net435 sg13g2_dlygate4sd3_1
Xhold88 s0.data_out\[16\]\[5\] VPWR VGND net457 sg13g2_dlygate4sd3_1
Xhold99 s0.shift_out\[15\][0] VPWR VGND net468 sg13g2_dlygate4sd3_1
XFILLER_29_643 VPWR VGND sg13g2_fill_1
Xhold77 s0.data_out\[9\]\[4\] VPWR VGND net446 sg13g2_dlygate4sd3_1
XFILLER_17_838 VPWR VGND sg13g2_fill_1
XFILLER_32_808 VPWR VGND sg13g2_fill_2
XFILLER_6_59 VPWR VGND sg13g2_fill_2
XFILLER_4_742 VPWR VGND sg13g2_fill_2
XFILLER_4_764 VPWR VGND sg13g2_fill_1
XFILLER_3_263 VPWR VGND sg13g2_fill_2
XFILLER_6_1008 VPWR VGND sg13g2_decap_8
XFILLER_0_992 VPWR VGND sg13g2_decap_8
XFILLER_48_963 VPWR VGND sg13g2_decap_8
XFILLER_37_1010 VPWR VGND sg13g2_decap_8
XFILLER_23_808 VPWR VGND sg13g2_decap_8
X_5740_ net1405 net1330 _1665_ VPWR VGND sg13g2_nor2b_1
X_5671_ net1425 VPWR _1604_ VGND _1544_ _1603_ sg13g2_o21ai_1
X_7410_ VGND VPWR _3172_ _3169_ net1678 sg13g2_or2_1
X_4622_ _0655_ s0.data_out\[23\]\[6\] net1530 VPWR VGND sg13g2_nand2b_1
X_4553_ VGND VPWR net1519 net407 _0592_ _0551_ sg13g2_a21oi_1
X_7341_ VGND VPWR _3359_ _3100_ _0072_ _3105_ sg13g2_a21oi_1
X_4484_ _0528_ VPWR _0529_ VGND _0516_ _0526_ sg13g2_o21ai_1
X_7272_ _3046_ s0.data_out\[2\]\[5\] net1245 VPWR VGND sg13g2_nand2b_1
X_6223_ VGND VPWR _1983_ _2099_ _2100_ net1365 sg13g2_a21oi_1
X_6154_ _2023_ _2032_ _2042_ _2043_ VPWR VGND sg13g2_nor3_1
X_7672__355 VPWR VGND net355 sg13g2_tiehi
X_5105_ _1075_ VPWR _1090_ VGND net1706 _1082_ sg13g2_o21ai_1
X_6085_ _1974_ net1372 net551 VPWR VGND sg13g2_nand2_1
X_5036_ VPWR _0184_ net684 VGND sg13g2_inv_1
XFILLER_39_985 VPWR VGND sg13g2_decap_8
X_6987_ s0.data_out\[5\]\[0\] s0.data_out\[4\]\[0\] net1255 _2785_ VPWR VGND sg13g2_mux2_1
X_5938_ _1843_ VPWR _1844_ VGND net1749 net696 sg13g2_o21ai_1
XFILLER_41_638 VPWR VGND sg13g2_fill_1
X_5869_ _1782_ net575 net1411 VPWR VGND sg13g2_nand2b_1
X_7608_ _3341_ _3337_ _3345_ _3346_ VPWR VGND sg13g2_a21o_1
X_7539_ _3287_ VPWR _3288_ VGND net1720 net799 sg13g2_o21ai_1
XFILLER_49_738 VPWR VGND sg13g2_decap_8
XFILLER_1_789 VPWR VGND sg13g2_decap_8
XFILLER_29_440 VPWR VGND sg13g2_fill_2
XFILLER_45_900 VPWR VGND sg13g2_decap_8
XFILLER_17_602 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_368 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_45_977 VPWR VGND sg13g2_decap_8
XFILLER_44_465 VPWR VGND sg13g2_fill_2
XFILLER_16_134 VPWR VGND sg13g2_fill_2
XFILLER_17_679 VPWR VGND sg13g2_fill_1
XFILLER_12_340 VPWR VGND sg13g2_fill_2
XFILLER_48_760 VPWR VGND sg13g2_decap_8
X_7890_ net120 VGND VPWR net399 s0.was_valid_out\[6\][0] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_6910_ _2594_ VPWR _2720_ VGND net1280 _3527_ sg13g2_o21ai_1
X_6841_ VGND VPWR _3363_ _2648_ _0024_ _2653_ sg13g2_a21oi_1
XFILLER_35_498 VPWR VGND sg13g2_fill_2
X_6772_ _2594_ net1281 s0.data_out\[6\]\[4\] VPWR VGND sg13g2_nand2_1
X_3984_ VPWR _3360_ net402 VGND sg13g2_inv_1
X_5723_ _1647_ VPWR _1648_ VGND net1197 _1645_ sg13g2_o21ai_1
X_5654_ _1511_ _1589_ _1590_ _1591_ VPWR VGND sg13g2_nor3_1
X_4605_ net1510 net1347 _0638_ VPWR VGND sg13g2_nor2b_1
Xhold311 s0.data_out\[21\]\[4\] VPWR VGND net680 sg13g2_dlygate4sd3_1
X_5585_ _1522_ net606 net1435 VPWR VGND sg13g2_nand2b_1
X_7324_ _3030_ _3090_ net1718 _3091_ VPWR VGND sg13g2_nand3_1
Xhold300 _0044_ VPWR VGND net669 sg13g2_dlygate4sd3_1
Xhold344 _2638_ VPWR VGND net713 sg13g2_dlygate4sd3_1
X_4536_ net1539 VPWR _0579_ VGND _0496_ _0578_ sg13g2_o21ai_1
Xhold322 s0.data_out\[20\]\[0\] VPWR VGND net691 sg13g2_dlygate4sd3_1
Xhold333 s0.data_out\[15\]\[1\] VPWR VGND net702 sg13g2_dlygate4sd3_1
Xhold355 _2073_ VPWR VGND net724 sg13g2_dlygate4sd3_1
Xhold377 s0.data_out\[12\]\[5\] VPWR VGND net746 sg13g2_dlygate4sd3_1
Xhold366 s0.data_out\[2\]\[3\] VPWR VGND net735 sg13g2_dlygate4sd3_1
X_4467_ VGND VPWR net1522 _0511_ _0512_ _0509_ sg13g2_a21oi_1
X_7255_ s0.data_out\[2\]\[6\] s0.data_out\[3\]\[6\] net1247 _3029_ VPWR VGND sg13g2_mux2_1
X_6206_ net1739 VPWR _2086_ VGND _2083_ _2085_ sg13g2_o21ai_1
Xhold388 s0.data_out\[13\]\[3\] VPWR VGND net757 sg13g2_dlygate4sd3_1
Xhold399 _1385_ VPWR VGND net768 sg13g2_dlygate4sd3_1
X_4398_ _0435_ _0451_ _0452_ _0454_ _0455_ VPWR VGND sg13g2_nor4_1
X_7186_ net1586 _2905_ _2968_ VPWR VGND sg13g2_nor2_1
X_6137_ net1370 net1340 _2026_ VPWR VGND sg13g2_nor2b_1
X_6068_ net1395 VPWR _1961_ VGND _1920_ _1960_ sg13g2_o21ai_1
X_5019_ _1014_ _1016_ net1682 _1017_ VPWR VGND sg13g2_nand3_1
XFILLER_27_922 VPWR VGND sg13g2_fill_2
XFILLER_26_56 VPWR VGND sg13g2_decap_8
XFILLER_42_947 VPWR VGND sg13g2_decap_8
XFILLER_27_999 VPWR VGND sg13g2_decap_8
XFILLER_21_170 VPWR VGND sg13g2_decap_4
XFILLER_42_99 VPWR VGND sg13g2_fill_1
XFILLER_10_899 VPWR VGND sg13g2_decap_4
XFILLER_27_1020 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_fill_2
XFILLER_49_535 VPWR VGND sg13g2_decap_8
X_7653__32 VPWR VGND net32 sg13g2_tiehi
XFILLER_17_443 VPWR VGND sg13g2_decap_8
XFILLER_18_988 VPWR VGND sg13g2_decap_8
XFILLER_9_653 VPWR VGND sg13g2_fill_1
X_5370_ VGND VPWR net1452 _1328_ _1331_ _1330_ sg13g2_a21oi_1
X_4321_ net1533 _0375_ _0381_ VPWR VGND sg13g2_nor2_1
X_4252_ _3615_ _3613_ _3616_ VPWR VGND _3614_ sg13g2_nand3b_1
X_7040_ _2838_ _2801_ _2837_ VPWR VGND sg13g2_nand2_1
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_1017 VPWR VGND sg13g2_decap_8
X_4183_ _3552_ net1647 net1165 VPWR VGND sg13g2_nand2_1
XFILLER_28_719 VPWR VGND sg13g2_decap_4
X_7942_ net63 VGND VPWR _0076_ s0.data_out\[2\]\[0\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_7847__166 VPWR VGND net166 sg13g2_tiehi
X_7873_ net138 VGND VPWR net548 s0.data_out\[8\]\[3\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_6824_ net1174 _3520_ _2639_ VPWR VGND sg13g2_nor2_1
XFILLER_23_435 VPWR VGND sg13g2_fill_2
X_6755_ net1276 net1329 _2577_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_479 VPWR VGND sg13g2_fill_2
X_5706_ _1629_ net1401 _1630_ _1631_ VPWR VGND sg13g2_a21o_1
Xclkbuf_leaf_30_clk clknet_3_5__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_6686_ net1599 _2440_ _2517_ VPWR VGND sg13g2_nor2_1
X_5637_ VGND VPWR net1426 _1571_ _1574_ _1573_ sg13g2_a21oi_1
X_5568_ net1428 VPWR _1508_ VGND net1644 net1416 sg13g2_o21ai_1
Xhold152 _0080_ VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold130 s0.data_out\[18\]\[4\] VPWR VGND net499 sg13g2_dlygate4sd3_1
Xhold141 _0202_ VPWR VGND net510 sg13g2_dlygate4sd3_1
X_4519_ _0561_ _0563_ net1679 _0564_ VPWR VGND sg13g2_nand3_1
X_7307_ _3077_ VPWR _3078_ VGND net1191 _3076_ sg13g2_o21ai_1
X_7854__159 VPWR VGND net159 sg13g2_tiehi
X_5499_ _1448_ _1447_ net1664 _1440_ net1654 VPWR VGND sg13g2_a22oi_1
Xhold174 _0236_ VPWR VGND net543 sg13g2_dlygate4sd3_1
Xhold163 s0.data_out\[6\]\[2\] VPWR VGND net532 sg13g2_dlygate4sd3_1
Xhold185 s0.data_out\[7\]\[2\] VPWR VGND net554 sg13g2_dlygate4sd3_1
X_7238_ net1695 _3011_ _3012_ VPWR VGND sg13g2_nor2_1
Xfanout1619 net1621 net1619 VPWR VGND sg13g2_buf_8
Xhold196 _0264_ VPWR VGND net565 sg13g2_dlygate4sd3_1
Xfanout1608 net1610 net1608 VPWR VGND sg13g2_buf_8
X_7169_ VGND VPWR net1241 s0.data_out\[3\]\[0\] _2954_ _2892_ sg13g2_a21oi_1
XFILLER_2_1022 VPWR VGND sg13g2_decap_8
X_7650__35 VPWR VGND net35 sg13g2_tiehi
XFILLER_27_741 VPWR VGND sg13g2_fill_1
XFILLER_42_733 VPWR VGND sg13g2_fill_2
XFILLER_23_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_21_clk clknet_3_7__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_5_166 VPWR VGND sg13g2_fill_1
XFILLER_2_840 VPWR VGND sg13g2_decap_8
XFILLER_18_763 VPWR VGND sg13g2_fill_1
XFILLER_17_240 VPWR VGND sg13g2_fill_2
X_4870_ VGND VPWR _0760_ _0878_ _0879_ net1499 sg13g2_a21oi_1
X_7929__77 VPWR VGND net77 sg13g2_tiehi
X_6540_ _2386_ _2377_ _2385_ VPWR VGND sg13g2_nand2_1
XFILLER_32_276 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_12_clk clknet_3_2__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_6471_ net1610 _2312_ _0333_ VPWR VGND sg13g2_nor2_1
X_5422_ net1624 _1341_ _1378_ VPWR VGND sg13g2_nor2_1
X_5353_ VGND VPWR _1200_ _1313_ _1314_ net1449 sg13g2_a21oi_1
X_4304_ net1559 VPWR _0367_ VGND _3622_ _0366_ sg13g2_o21ai_1
X_5284_ net1447 s0.data_out\[18\]\[1\] _1255_ VPWR VGND sg13g2_and2_1
X_4235_ net1558 _3597_ _3598_ _3599_ VPWR VGND sg13g2_nor3_1
X_7023_ net1252 net1343 _2821_ VPWR VGND sg13g2_nor2b_1
X_4166_ VPWR _3542_ net769 VGND sg13g2_inv_1
X_4097_ VPWR _3473_ net765 VGND sg13g2_inv_1
X_7925_ net82 VGND VPWR _0059_ s0.data_out\[4\]\[7\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_7856_ net156 VGND VPWR _0334_ s0.genblk1\[8\].modules.bubble clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_6807_ net1284 VPWR _2626_ VGND _2545_ _2625_ sg13g2_o21ai_1
X_4999_ VGND VPWR net1483 _0994_ _0997_ _0996_ sg13g2_a21oi_1
XFILLER_23_287 VPWR VGND sg13g2_fill_1
XFILLER_23_298 VPWR VGND sg13g2_fill_1
X_7860__152 VPWR VGND net152 sg13g2_tiehi
X_7787_ net231 VGND VPWR _0265_ s0.was_valid_out\[14\][0] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_6738_ VGND VPWR net1271 _2558_ _2560_ _2559_ sg13g2_a21oi_1
X_6669_ _2466_ _2484_ _2502_ _2503_ VPWR VGND sg13g2_or3_1
X_7717__306 VPWR VGND net306 sg13g2_tiehi
Xfanout1405 net1407 net1405 VPWR VGND sg13g2_buf_1
Xfanout1438 net460 net1438 VPWR VGND sg13g2_buf_1
Xfanout1427 net1430 net1427 VPWR VGND sg13g2_buf_1
Xfanout1416 net1418 net1416 VPWR VGND sg13g2_buf_1
Xfanout1449 net1452 net1449 VPWR VGND sg13g2_buf_8
XFILLER_47_836 VPWR VGND sg13g2_decap_8
XFILLER_46_313 VPWR VGND sg13g2_fill_1
XFILLER_46_335 VPWR VGND sg13g2_fill_2
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_7_976 VPWR VGND sg13g2_decap_8
X_7837__176 VPWR VGND net176 sg13g2_tiehi
X_4020_ _3396_ net1274 VPWR VGND sg13g2_inv_2
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_38_858 VPWR VGND sg13g2_fill_1
X_5971_ _1869_ _1871_ net1708 _1872_ VPWR VGND sg13g2_nand3_1
X_4922_ net1486 s0.data_out\[21\]\[4\] _0926_ VPWR VGND sg13g2_and2_1
X_7710_ net314 VGND VPWR _0188_ s0.data_out\[21\]\[4\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_33_530 VPWR VGND sg13g2_fill_2
X_7844__169 VPWR VGND net169 sg13g2_tiehi
X_7641_ net45 VGND VPWR net473 s0.data_out\[27\]\[6\] clknet_leaf_0_clk sg13g2_dfrbpq_2
X_4853_ _0862_ s0.data_out\[21\]\[3\] net1506 VPWR VGND sg13g2_nand2b_1
X_7572_ _3313_ VPWR _3314_ VGND net1202 _3312_ sg13g2_o21ai_1
X_4784_ _0162_ _0801_ _0802_ _3436_ net1595 VPWR VGND sg13g2_a22oi_1
X_7959__256 VPWR VGND net256 sg13g2_tiehi
X_6523_ _2369_ net1303 net426 VPWR VGND sg13g2_nand2_1
X_6454_ VPWR _0330_ _2304_ VGND sg13g2_inv_1
X_5405_ VPWR _0221_ _1364_ VGND sg13g2_inv_1
X_6385_ VGND VPWR net1323 _2240_ _2243_ _2242_ sg13g2_a21oi_1
X_5336_ _1185_ VPWR _1297_ VGND net1453 _3465_ sg13g2_o21ai_1
X_5267_ VGND VPWR _1118_ _1239_ _1240_ net1461 sg13g2_a21oi_1
X_4218_ s0.data_out\[27\]\[0\] s0.data_out\[26\]\[0\] net1555 _3582_ VPWR VGND sg13g2_mux2_1
X_7006_ net1251 net1328 _2804_ VPWR VGND sg13g2_nor2b_1
X_5198_ _1174_ _1171_ _1173_ VPWR VGND sg13g2_nand2_1
XFILLER_18_57 VPWR VGND sg13g2_fill_1
X_4149_ VPWR _3525_ net584 VGND sg13g2_inv_1
XFILLER_29_858 VPWR VGND sg13g2_fill_2
XFILLER_44_828 VPWR VGND sg13g2_decap_8
X_7908_ net100 VGND VPWR net581 s0.data_out\[5\]\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_2
XFILLER_24_563 VPWR VGND sg13g2_fill_1
X_7839_ net174 VGND VPWR _0317_ s0.data_new_delayed\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_2
XFILLER_34_78 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_3_3__leaf_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_11_268 VPWR VGND sg13g2_fill_2
X_7916__91 VPWR VGND net91 sg13g2_tiehi
XFILLER_4_913 VPWR VGND sg13g2_decap_8
Xfanout1213 s0.shift_out\[0\][0] net1213 VPWR VGND sg13g2_buf_2
Xfanout1202 _3378_ net1202 VPWR VGND sg13g2_buf_8
XFILLER_3_489 VPWR VGND sg13g2_fill_2
Xfanout1224 net1227 net1224 VPWR VGND sg13g2_buf_8
Xfanout1235 net828 net1235 VPWR VGND sg13g2_buf_8
Xfanout1246 net824 net1246 VPWR VGND sg13g2_buf_8
Xfanout1257 s0.valid_out\[4\][0] net1257 VPWR VGND sg13g2_buf_2
Xfanout1268 net1269 net1268 VPWR VGND sg13g2_buf_8
Xfanout1279 s0.valid_out\[6\][0] net1279 VPWR VGND sg13g2_buf_1
XFILLER_47_644 VPWR VGND sg13g2_decap_4
XFILLER_35_806 VPWR VGND sg13g2_fill_1
XFILLER_46_165 VPWR VGND sg13g2_fill_2
X_7908__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_43_872 VPWR VGND sg13g2_decap_8
X_7798__219 VPWR VGND net219 sg13g2_tiehi
X_6170_ _0294_ _2055_ _2056_ _3491_ net1614 VPWR VGND sg13g2_a22oi_1
X_5121_ VGND VPWR net1473 _1103_ _1106_ _1105_ sg13g2_a21oi_1
XFILLER_34_2 VPWR VGND sg13g2_fill_1
X_5052_ VGND VPWR net1180 _1015_ _1045_ net1606 sg13g2_a21oi_1
X_4003_ VPWR _3379_ net1462 VGND sg13g2_inv_1
XFILLER_37_165 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_20 VPWR VGND uio_out[4] sg13g2_tielo
X_5954_ VGND VPWR _3364_ _1852_ _0277_ _1857_ sg13g2_a21oi_1
XFILLER_40_319 VPWR VGND sg13g2_fill_1
X_4905_ net1501 VPWR _0913_ VGND _0851_ _0912_ sg13g2_o21ai_1
X_5885_ _1797_ VPWR _1798_ VGND net1400 _3478_ sg13g2_o21ai_1
X_7624_ VGND VPWR net1722 _3343_ _0104_ _3356_ sg13g2_a21oi_1
X_4836_ net1487 net1355 _0845_ VPWR VGND sg13g2_nor2b_1
X_7555_ VGND VPWR net1211 net434 _3300_ _3271_ sg13g2_a21oi_1
X_6506_ s0.data_out\[9\]\[7\] s0.data_out\[8\]\[7\] net1304 _2352_ VPWR VGND sg13g2_mux2_1
X_4767_ VGND VPWR _0775_ _0777_ _0788_ net1671 sg13g2_a21oi_1
X_7486_ _3130_ VPWR _3236_ VGND net1226 _3543_ sg13g2_o21ai_1
X_4698_ _0718_ VPWR _0719_ VGND net1504 _3436_ sg13g2_o21ai_1
X_6437_ net1308 net544 _2291_ VPWR VGND sg13g2_and2_1
X_6368_ _2212_ VPWR _2226_ VGND net1705 _2219_ sg13g2_o21ai_1
X_5319_ VGND VPWR _1283_ net1456 net428 sg13g2_or2_1
Xhold23 s0.genblk1\[18\].modules.bubble VPWR VGND net392 sg13g2_dlygate4sd3_1
Xhold12 s0.genblk1\[3\].modules.bubble VPWR VGND net381 sg13g2_dlygate4sd3_1
X_6299_ net1366 VPWR _2172_ VGND _2112_ _2171_ sg13g2_o21ai_1
Xhold45 s0.data_out\[7\]\[7\] VPWR VGND net414 sg13g2_dlygate4sd3_1
Xhold56 s0.was_valid_out\[22\][0] VPWR VGND net425 sg13g2_dlygate4sd3_1
Xhold34 _0060_ VPWR VGND net403 sg13g2_dlygate4sd3_1
XFILLER_29_45 VPWR VGND sg13g2_fill_1
XFILLER_29_56 VPWR VGND sg13g2_fill_1
Xhold78 s0.data_out\[0\]\[7\] VPWR VGND net447 sg13g2_dlygate4sd3_1
Xhold67 _1123_ VPWR VGND net436 sg13g2_dlygate4sd3_1
Xhold89 _1580_ VPWR VGND net458 sg13g2_dlygate4sd3_1
XFILLER_21_1026 VPWR VGND sg13g2_fill_2
XFILLER_44_625 VPWR VGND sg13g2_decap_8
XFILLER_16_316 VPWR VGND sg13g2_fill_2
XFILLER_12_511 VPWR VGND sg13g2_fill_1
XFILLER_8_504 VPWR VGND sg13g2_decap_8
XFILLER_40_875 VPWR VGND sg13g2_fill_2
XFILLER_8_559 VPWR VGND sg13g2_fill_1
XFILLER_12_599 VPWR VGND sg13g2_fill_1
XFILLER_3_231 VPWR VGND sg13g2_fill_2
XFILLER_0_971 VPWR VGND sg13g2_decap_8
XFILLER_48_942 VPWR VGND sg13g2_decap_8
XFILLER_19_143 VPWR VGND sg13g2_fill_2
XFILLER_35_636 VPWR VGND sg13g2_fill_1
X_7665__363 VPWR VGND net363 sg13g2_tiehi
X_5670_ net1197 _3473_ _1603_ VPWR VGND sg13g2_nor2_1
XFILLER_30_330 VPWR VGND sg13g2_fill_2
XFILLER_31_864 VPWR VGND sg13g2_decap_4
X_4621_ _0652_ net1509 _0653_ _0654_ VPWR VGND sg13g2_a21o_1
XFILLER_31_886 VPWR VGND sg13g2_fill_1
X_4552_ VPWR _0141_ _0591_ VGND sg13g2_inv_1
X_7340_ net1718 VPWR _3105_ VGND _3102_ _3104_ sg13g2_o21ai_1
XFILLER_7_592 VPWR VGND sg13g2_fill_2
X_4483_ _0528_ net1687 _0525_ VPWR VGND sg13g2_nand2_1
X_7271_ _3043_ net1232 _3044_ _3045_ VPWR VGND sg13g2_a21o_1
X_6222_ _2099_ net589 net1372 VPWR VGND sg13g2_nand2b_1
X_6153_ net1675 _2030_ _2042_ VPWR VGND sg13g2_nor2_1
X_6084_ net1739 net390 _0291_ VPWR VGND sg13g2_and2_1
X_5104_ VPWR VGND _1088_ net1712 _1086_ net1706 _1089_ _1082_ sg13g2_a221oi_1
XFILLER_39_964 VPWR VGND sg13g2_decap_8
X_5035_ _1031_ VPWR _1032_ VGND net1735 net683 sg13g2_o21ai_1
XFILLER_38_441 VPWR VGND sg13g2_fill_1
XFILLER_41_606 VPWR VGND sg13g2_fill_1
X_6986_ VGND VPWR net1260 _2781_ _2784_ _2783_ sg13g2_a21oi_1
XFILLER_25_135 VPWR VGND sg13g2_fill_2
XFILLER_25_157 VPWR VGND sg13g2_fill_1
XFILLER_26_669 VPWR VGND sg13g2_fill_1
X_5937_ _1842_ net1749 _1843_ VPWR VGND _1790_ sg13g2_nand3b_1
XFILLER_41_628 VPWR VGND sg13g2_fill_2
X_5868_ _1779_ net1395 _1780_ _1781_ VPWR VGND sg13g2_a21o_1
X_7607_ _3344_ VPWR _3345_ VGND net1689 _3340_ sg13g2_o21ai_1
X_4819_ net412 net1505 _0831_ VPWR VGND sg13g2_nor2_1
X_5799_ net1414 VPWR _1720_ VGND _1654_ _1719_ sg13g2_o21ai_1
X_7538_ _3228_ _3286_ net1720 _3287_ VPWR VGND sg13g2_nand3_1
XFILLER_5_507 VPWR VGND sg13g2_fill_2
X_7469_ net1201 _3218_ _3219_ VPWR VGND sg13g2_nor2_1
XFILLER_1_702 VPWR VGND sg13g2_fill_1
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_1_768 VPWR VGND sg13g2_decap_8
XFILLER_49_717 VPWR VGND sg13g2_decap_8
X_7968__119 VPWR VGND net119 sg13g2_tiehi
X_7788__229 VPWR VGND net229 sg13g2_tiehi
Xheichips25_top_sorter_369 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_29_452 VPWR VGND sg13g2_fill_1
XFILLER_45_956 VPWR VGND sg13g2_decap_8
XFILLER_44_400 VPWR VGND sg13g2_fill_1
XFILLER_31_105 VPWR VGND sg13g2_fill_2
X_7905__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_40_672 VPWR VGND sg13g2_fill_2
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
X_6840_ net1729 VPWR _2653_ VGND _2650_ _2652_ sg13g2_o21ai_1
X_6771_ net1276 s0.data_new_delayed\[4\] _2593_ VPWR VGND sg13g2_nor2b_1
X_3983_ VPWR _3359_ net421 VGND sg13g2_inv_1
X_5722_ _1647_ net1197 _1646_ VPWR VGND sg13g2_nand2_1
X_5653_ _1564_ _1565_ _1590_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_694 VPWR VGND sg13g2_fill_2
X_4604_ s0.data_out\[24\]\[3\] s0.data_out\[23\]\[3\] net1518 _0637_ VPWR VGND sg13g2_mux2_1
X_5584_ _1519_ net1413 _1520_ _1521_ VPWR VGND sg13g2_a21o_1
X_4535_ net1522 net481 _0578_ VPWR VGND sg13g2_and2_1
X_7323_ net1239 VPWR _3090_ VGND _3026_ _3089_ sg13g2_o21ai_1
Xhold301 s0.data_out\[4\]\[4\] VPWR VGND net670 sg13g2_dlygate4sd3_1
Xhold312 s0.data_out\[17\]\[4\] VPWR VGND net681 sg13g2_dlygate4sd3_1
Xhold323 s0.data_out\[12\]\[0\] VPWR VGND net692 sg13g2_dlygate4sd3_1
Xhold334 _0258_ VPWR VGND net703 sg13g2_dlygate4sd3_1
Xhold345 s0.data_out\[1\]\[4\] VPWR VGND net714 sg13g2_dlygate4sd3_1
Xhold367 _0079_ VPWR VGND net736 sg13g2_dlygate4sd3_1
X_4466_ _0510_ VPWR _0511_ VGND net1529 _3423_ sg13g2_o21ai_1
X_7254_ _3028_ net1239 _3027_ VPWR VGND sg13g2_nand2b_1
Xhold378 s0.data_out\[10\]\[4\] VPWR VGND net747 sg13g2_dlygate4sd3_1
Xhold356 s0.data_out\[2\]\[6\] VPWR VGND net725 sg13g2_dlygate4sd3_1
X_6205_ _2084_ VPWR _2085_ VGND _2079_ _2082_ sg13g2_o21ai_1
X_4397_ _0453_ VPWR _0454_ VGND net1677 _0442_ sg13g2_o21ai_1
X_7185_ net1249 VPWR _2967_ VGND _2902_ _2966_ sg13g2_o21ai_1
Xhold389 _0284_ VPWR VGND net758 sg13g2_dlygate4sd3_1
X_6136_ s0.data_out\[12\]\[5\] s0.data_out\[11\]\[5\] net1375 _2025_ VPWR VGND sg13g2_mux2_1
XFILLER_46_709 VPWR VGND sg13g2_decap_8
X_6067_ net1383 net540 _1960_ VPWR VGND sg13g2_and2_1
XFILLER_39_750 VPWR VGND sg13g2_fill_1
X_5018_ _1016_ net1180 _1015_ VPWR VGND sg13g2_nand2_1
XFILLER_26_444 VPWR VGND sg13g2_decap_4
XFILLER_27_978 VPWR VGND sg13g2_decap_8
XFILLER_42_926 VPWR VGND sg13g2_decap_8
X_6969_ net1726 VPWR _2770_ VGND _2767_ _2769_ sg13g2_o21ai_1
XFILLER_18_945 VPWR VGND sg13g2_fill_1
XFILLER_45_764 VPWR VGND sg13g2_decap_8
XFILLER_45_786 VPWR VGND sg13g2_decap_4
X_7662__366 VPWR VGND net366 sg13g2_tiehi
X_4320_ _0377_ VPWR _0380_ VGND net419 net1540 sg13g2_o21ai_1
XFILLER_5_893 VPWR VGND sg13g2_decap_4
X_4251_ VGND VPWR _3615_ _3612_ net1658 sg13g2_or2_1
X_4182_ VGND VPWR _3402_ net1165 net9 _3551_ sg13g2_a21oi_1
X_7941_ net64 VGND VPWR _0075_ s0.shift_out\[2\][0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_7872_ net139 VGND VPWR _0006_ s0.data_out\[8\]\[2\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_6823_ VPWR _0021_ net713 VGND sg13g2_inv_1
X_6754_ s0.data_out\[7\]\[7\] s0.data_out\[6\]\[7\] net1281 _2576_ VPWR VGND sg13g2_mux2_1
X_6685_ net1293 VPWR _2516_ VGND _2437_ _2515_ sg13g2_o21ai_1
X_5705_ net1401 s0.data_new_delayed\[1\] _1630_ VPWR VGND sg13g2_nor2b_1
X_5636_ VGND VPWR _1462_ _1572_ _1573_ net1427 sg13g2_a21oi_1
XFILLER_3_819 VPWR VGND sg13g2_decap_8
X_5567_ _0240_ _1506_ _1507_ _3462_ net1623 VPWR VGND sg13g2_a22oi_1
Xhold153 s0.data_out\[10\]\[7\] VPWR VGND net522 sg13g2_dlygate4sd3_1
X_4518_ _0563_ net1184 _0562_ VPWR VGND sg13g2_nand2_1
Xhold120 s0.data_out\[24\]\[6\] VPWR VGND net489 sg13g2_dlygate4sd3_1
Xhold131 _0213_ VPWR VGND net500 sg13g2_dlygate4sd3_1
X_5498_ VGND VPWR net1440 _1444_ _1447_ _1446_ sg13g2_a21oi_1
Xhold142 s0.data_out\[21\]\[2\] VPWR VGND net511 sg13g2_dlygate4sd3_1
X_7306_ VGND VPWR net1191 _3010_ _3077_ net1582 sg13g2_a21oi_1
X_4449_ _0494_ net1528 net481 VPWR VGND sg13g2_nand2_1
Xhold164 _2743_ VPWR VGND net533 sg13g2_dlygate4sd3_1
Xhold186 _0018_ VPWR VGND net555 sg13g2_dlygate4sd3_1
X_7237_ VGND VPWR net1191 _3010_ _3011_ _3009_ sg13g2_a21oi_1
Xhold175 s0.data_out\[9\]\[3\] VPWR VGND net544 sg13g2_dlygate4sd3_1
Xhold197 s0.data_out\[5\]\[7\] VPWR VGND net566 sg13g2_dlygate4sd3_1
Xfanout1609 net1610 net1609 VPWR VGND sg13g2_buf_1
X_7168_ _2952_ _2953_ _0051_ VPWR VGND sg13g2_and2_1
X_6119_ net1371 net1335 _2008_ VPWR VGND sg13g2_nor2b_1
X_7099_ net1240 net1352 _2885_ VPWR VGND sg13g2_nor2b_1
XFILLER_19_709 VPWR VGND sg13g2_fill_2
XFILLER_37_45 VPWR VGND sg13g2_fill_2
XFILLER_37_34 VPWR VGND sg13g2_fill_1
XFILLER_2_1001 VPWR VGND sg13g2_decap_8
XFILLER_18_208 VPWR VGND sg13g2_fill_2
XFILLER_27_720 VPWR VGND sg13g2_fill_1
XFILLER_26_241 VPWR VGND sg13g2_fill_2
XFILLER_26_252 VPWR VGND sg13g2_fill_1
XFILLER_18_1009 VPWR VGND sg13g2_decap_8
XFILLER_23_970 VPWR VGND sg13g2_decap_8
XFILLER_30_907 VPWR VGND sg13g2_fill_2
XFILLER_10_664 VPWR VGND sg13g2_fill_2
XFILLER_6_657 VPWR VGND sg13g2_fill_2
XFILLER_2_896 VPWR VGND sg13g2_decap_8
XFILLER_45_561 VPWR VGND sg13g2_fill_1
XFILLER_14_981 VPWR VGND sg13g2_decap_8
XFILLER_20_428 VPWR VGND sg13g2_fill_1
XFILLER_9_462 VPWR VGND sg13g2_decap_4
X_6470_ _2313_ _2318_ _0332_ VPWR VGND sg13g2_nor2_1
X_5421_ net1450 VPWR _1377_ VGND _1338_ _1376_ sg13g2_o21ai_1
X_5352_ _1313_ s0.data_out\[17\]\[3\] net1456 VPWR VGND sg13g2_nand2b_1
X_4303_ net1545 s0.data_out\[26\]\[5\] _0366_ VPWR VGND sg13g2_and2_1
X_7853__160 VPWR VGND net160 sg13g2_tiehi
XFILLER_4_60 VPWR VGND sg13g2_fill_2
X_5283_ VPWR _0209_ net648 VGND sg13g2_inv_1
X_7022_ s0.data_out\[5\]\[4\] s0.data_out\[4\]\[4\] net1256 _2820_ VPWR VGND sg13g2_mux2_1
X_4234_ net1563 s0.data_out\[26\]\[7\] _3598_ VPWR VGND sg13g2_nor2_1
X_4165_ VPWR _3541_ s0.data_out\[1\]\[5\] VGND sg13g2_inv_1
XFILLER_28_506 VPWR VGND sg13g2_decap_8
X_4096_ VPWR _3472_ net564 VGND sg13g2_inv_1
XFILLER_36_550 VPWR VGND sg13g2_fill_1
X_7924_ net83 VGND VPWR net537 s0.data_out\[4\]\[6\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_7855_ net157 VGND VPWR _0333_ s0.valid_out\[9\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_36_583 VPWR VGND sg13g2_decap_4
X_6806_ net1175 _3522_ _2625_ VPWR VGND sg13g2_nor2_1
XFILLER_24_767 VPWR VGND sg13g2_fill_2
X_4998_ VGND VPWR _0874_ _0995_ _0996_ net1483 sg13g2_a21oi_1
X_7786_ net232 VGND VPWR net565 s0.data_out\[15\]\[7\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_23_69 VPWR VGND sg13g2_fill_2
X_6737_ net1271 net1357 _2559_ VPWR VGND sg13g2_nor2b_1
X_6668_ _2502_ _2497_ _2501_ VPWR VGND sg13g2_nand2_1
XFILLER_20_984 VPWR VGND sg13g2_decap_8
X_6599_ net1601 _2428_ _0001_ VPWR VGND sg13g2_nor2_1
X_5619_ VGND VPWR net1428 _1553_ _1556_ _1555_ sg13g2_a21oi_1
Xfanout1406 net1407 net1406 VPWR VGND sg13g2_buf_8
Xfanout1439 net1442 net1439 VPWR VGND sg13g2_buf_8
Xfanout1428 net1430 net1428 VPWR VGND sg13g2_buf_8
Xfanout1417 net1418 net1417 VPWR VGND sg13g2_buf_8
XFILLER_47_815 VPWR VGND sg13g2_decap_8
XFILLER_34_509 VPWR VGND sg13g2_fill_2
XFILLER_15_734 VPWR VGND sg13g2_fill_1
XFILLER_30_726 VPWR VGND sg13g2_decap_8
XFILLER_7_900 VPWR VGND sg13g2_fill_1
XFILLER_11_940 VPWR VGND sg13g2_fill_2
XFILLER_14_299 VPWR VGND sg13g2_fill_1
XFILLER_31_1006 VPWR VGND sg13g2_decap_8
XFILLER_11_984 VPWR VGND sg13g2_decap_8
XFILLER_7_955 VPWR VGND sg13g2_decap_8
XFILLER_13_91 VPWR VGND sg13g2_fill_1
XFILLER_37_369 VPWR VGND sg13g2_fill_1
X_5970_ _1871_ net1192 _1870_ VPWR VGND sg13g2_nand2_1
X_4921_ _0176_ _0924_ _0925_ _3439_ net1605 VPWR VGND sg13g2_a22oi_1
XFILLER_18_572 VPWR VGND sg13g2_decap_4
X_7640_ net46 VGND VPWR net462 s0.data_out\[27\]\[5\] clknet_leaf_0_clk sg13g2_dfrbpq_2
X_4852_ _0860_ net1486 _0858_ _0861_ VPWR VGND sg13g2_a21o_1
X_7571_ VGND VPWR net1202 _3244_ _3313_ net1583 sg13g2_a21oi_1
X_4783_ net1595 _0723_ _0802_ VPWR VGND sg13g2_nor2_1
X_6522_ _2365_ _2366_ _2368_ VPWR VGND _2367_ sg13g2_nand3b_1
X_6453_ net833 VPWR _2304_ VGND net1741 net720 sg13g2_o21ai_1
XFILLER_9_281 VPWR VGND sg13g2_fill_1
X_5404_ _1363_ VPWR _1364_ VGND net1743 net779 sg13g2_o21ai_1
X_6384_ VGND VPWR _2126_ _2241_ _2242_ net1323 sg13g2_a21oi_1
X_5335_ _1296_ net1448 _1295_ VPWR VGND sg13g2_nand2b_1
X_5266_ _1239_ net499 net1466 VPWR VGND sg13g2_nand2b_1
X_4217_ _3581_ net1557 s0.data_out\[26\]\[0\] VPWR VGND sg13g2_nand2_1
X_7005_ s0.data_out\[5\]\[7\] s0.data_out\[4\]\[7\] net1255 _2803_ VPWR VGND sg13g2_mux2_1
X_5197_ net1198 VPWR _1173_ VGND s0.was_valid_out\[18\][0] net1466 sg13g2_o21ai_1
XFILLER_29_826 VPWR VGND sg13g2_fill_2
X_4148_ VPWR _3524_ net566 VGND sg13g2_inv_1
X_4079_ VPWR _3455_ net634 VGND sg13g2_inv_1
XFILLER_43_328 VPWR VGND sg13g2_fill_2
X_7907_ net101 VGND VPWR _0041_ s0.data_out\[5\]\[1\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_24_531 VPWR VGND sg13g2_fill_1
X_7723__300 VPWR VGND net300 sg13g2_tiehi
X_7838_ net175 VGND VPWR _0316_ s0.data_new_delayed\[1\] clknet_leaf_2_clk sg13g2_dfrbpq_2
X_7769_ net250 VGND VPWR net656 s0.data_out\[16\]\[2\] clknet_leaf_29_clk sg13g2_dfrbpq_1
Xclkload1 clknet_3_5__leaf_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_20_792 VPWR VGND sg13g2_fill_1
XFILLER_4_969 VPWR VGND sg13g2_decap_8
XFILLER_3_446 VPWR VGND sg13g2_fill_1
Xfanout1214 net1216 net1214 VPWR VGND sg13g2_buf_8
Xfanout1203 net1205 net1203 VPWR VGND sg13g2_buf_8
Xfanout1225 net1227 net1225 VPWR VGND sg13g2_buf_1
Xfanout1247 s0.valid_out\[3\][0] net1247 VPWR VGND sg13g2_buf_8
Xfanout1236 s0.valid_out\[2\][0] net1236 VPWR VGND sg13g2_buf_2
Xfanout1269 net827 net1269 VPWR VGND sg13g2_buf_8
Xfanout1258 net1259 net1258 VPWR VGND sg13g2_buf_8
XFILLER_47_689 VPWR VGND sg13g2_decap_8
XFILLER_30_512 VPWR VGND sg13g2_fill_1
X_7843__170 VPWR VGND net170 sg13g2_tiehi
XFILLER_30_567 VPWR VGND sg13g2_decap_8
XFILLER_30_578 VPWR VGND sg13g2_fill_2
X_5120_ VGND VPWR _0991_ _1104_ _1105_ net1474 sg13g2_a21oi_1
XFILLER_3_991 VPWR VGND sg13g2_decap_8
X_5051_ VGND VPWR net1469 net563 _1044_ _1012_ sg13g2_a21oi_1
X_4002_ VPWR _3378_ net1220 VGND sg13g2_inv_1
XFILLER_38_612 VPWR VGND sg13g2_fill_1
X_7850__163 VPWR VGND net163 sg13g2_tiehi
XFILLER_37_122 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_21 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_26_818 VPWR VGND sg13g2_fill_1
XFILLER_37_188 VPWR VGND sg13g2_fill_2
XFILLER_18_380 VPWR VGND sg13g2_fill_2
X_5953_ net1747 VPWR _1857_ VGND _1854_ _1856_ sg13g2_o21ai_1
X_7707__317 VPWR VGND net317 sg13g2_tiehi
X_4904_ net1487 s0.data_out\[21\]\[0\] _0912_ VPWR VGND sg13g2_and2_1
X_5884_ _1797_ net1400 net574 VPWR VGND sg13g2_nand2_1
X_7623_ net1722 net434 _3356_ VPWR VGND sg13g2_nor2_1
X_4835_ _0843_ VPWR _0844_ VGND net1491 _3440_ sg13g2_o21ai_1
X_7554_ VPWR _0091_ net615 VGND sg13g2_inv_1
X_4766_ VGND VPWR _0782_ _0784_ _0787_ net1679 sg13g2_a21oi_1
XFILLER_14_1023 VPWR VGND sg13g2_decap_4
X_6505_ _2351_ net1303 net561 VPWR VGND sg13g2_nand2_1
X_7485_ _3233_ VPWR _3235_ VGND net1695 _3220_ sg13g2_o21ai_1
X_4697_ _0718_ net1503 net599 VPWR VGND sg13g2_nand2_1
X_7913__95 VPWR VGND net95 sg13g2_tiehi
X_6436_ _0326_ _2289_ _2290_ _3500_ net1608 VPWR VGND sg13g2_a22oi_1
X_6367_ _2225_ _2224_ net1319 VPWR VGND sg13g2_nand2b_1
X_5318_ net1439 _1277_ _1282_ VPWR VGND sg13g2_nor2_1
Xhold13 s0.module0.bubble VPWR VGND net382 sg13g2_dlygate4sd3_1
X_6298_ net1322 net443 _2171_ VPWR VGND sg13g2_and2_1
Xhold46 _2580_ VPWR VGND net415 sg13g2_dlygate4sd3_1
Xhold35 s0.data_out\[0\]\[6\] VPWR VGND net404 sg13g2_dlygate4sd3_1
X_5249_ VGND VPWR net1461 _1219_ _1222_ _1221_ sg13g2_a21oi_1
Xhold24 s0.genblk1\[17\].modules.bubble VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold57 s0.data_out\[8\]\[5\] VPWR VGND net426 sg13g2_dlygate4sd3_1
Xhold68 s0.was_valid_out\[19\][0] VPWR VGND net437 sg13g2_dlygate4sd3_1
Xhold79 s0.data_out\[27\]\[3\] VPWR VGND net448 sg13g2_dlygate4sd3_1
XFILLER_21_1005 VPWR VGND sg13g2_decap_8
XFILLER_28_133 VPWR VGND sg13g2_decap_8
XFILLER_29_689 VPWR VGND sg13g2_fill_1
XFILLER_28_199 VPWR VGND sg13g2_decap_8
XFILLER_45_67 VPWR VGND sg13g2_fill_1
XFILLER_40_821 VPWR VGND sg13g2_fill_1
X_7827__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_25_884 VPWR VGND sg13g2_decap_4
X_7797__220 VPWR VGND net220 sg13g2_tiehi
XFILLER_8_549 VPWR VGND sg13g2_fill_2
XFILLER_0_950 VPWR VGND sg13g2_decap_8
XFILLER_48_921 VPWR VGND sg13g2_decap_8
XFILLER_48_998 VPWR VGND sg13g2_decap_8
XFILLER_16_840 VPWR VGND sg13g2_fill_1
XFILLER_42_191 VPWR VGND sg13g2_fill_1
X_4620_ net1508 net1334 _0653_ VPWR VGND sg13g2_nor2b_1
X_4551_ _0590_ VPWR _0591_ VGND net1725 net431 sg13g2_o21ai_1
XFILLER_7_571 VPWR VGND sg13g2_decap_8
X_4482_ _0508_ _0517_ _0518_ _0526_ _0527_ VPWR VGND sg13g2_nor4_1
X_7270_ net1233 net1339 _3044_ VPWR VGND sg13g2_nor2b_1
X_7910__98 VPWR VGND net98 sg13g2_tiehi
X_6221_ _2096_ net1321 _2097_ _2098_ VPWR VGND sg13g2_a21o_1
X_6152_ _2037_ _2039_ net1684 _2041_ VPWR VGND sg13g2_nand3_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_44_1016 VPWR VGND sg13g2_decap_8
X_5103_ _1088_ _1087_ net1472 VPWR VGND sg13g2_nand2b_1
XFILLER_32_0 VPWR VGND sg13g2_fill_1
X_6083_ net1628 _1967_ _0290_ VPWR VGND sg13g2_nor2_1
XFILLER_39_943 VPWR VGND sg13g2_decap_8
X_5034_ _1030_ VPWR _1031_ VGND net1178 _1029_ sg13g2_o21ai_1
X_6985_ VGND VPWR _2654_ _2782_ _2783_ net1260 sg13g2_a21oi_1
X_5936_ net1407 VPWR _1842_ VGND _1787_ _1841_ sg13g2_o21ai_1
X_7606_ _3344_ _3406_ _3343_ VPWR VGND sg13g2_nand2b_1
X_5867_ net1394 net1331 _1780_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_331 VPWR VGND sg13g2_fill_1
XFILLER_21_342 VPWR VGND sg13g2_fill_1
X_4818_ net1482 _0824_ _0830_ VPWR VGND sg13g2_nor2_1
X_7720__303 VPWR VGND net303 sg13g2_tiehi
X_5798_ net1195 _3479_ _1719_ VPWR VGND sg13g2_nor2_1
X_7537_ net1220 VPWR _3286_ VGND _3230_ _3285_ sg13g2_o21ai_1
X_4749_ _0767_ _0768_ _0770_ VPWR VGND _0769_ sg13g2_nand3b_1
XFILLER_5_519 VPWR VGND sg13g2_fill_2
X_7468_ VGND VPWR net1212 _3216_ _3218_ _3217_ sg13g2_a21oi_1
X_6419_ _2254_ _2276_ _2277_ VPWR VGND sg13g2_nor2b_1
X_7399_ _3403_ _3160_ _3161_ VPWR VGND sg13g2_and2_1
XFILLER_0_235 VPWR VGND sg13g2_decap_4
XFILLER_1_747 VPWR VGND sg13g2_decap_8
XFILLER_5_1021 VPWR VGND sg13g2_decap_8
XFILLER_45_935 VPWR VGND sg13g2_decap_8
XFILLER_13_810 VPWR VGND sg13g2_fill_1
XFILLER_16_169 VPWR VGND sg13g2_fill_1
XFILLER_31_117 VPWR VGND sg13g2_fill_2
XFILLER_31_139 VPWR VGND sg13g2_fill_1
XFILLER_40_684 VPWR VGND sg13g2_fill_2
XFILLER_12_386 VPWR VGND sg13g2_fill_1
X_7840__173 VPWR VGND net173 sg13g2_tiehi
XFILLER_48_795 VPWR VGND sg13g2_decap_8
XFILLER_36_979 VPWR VGND sg13g2_decap_8
X_6770_ _2592_ _2589_ _2590_ _2591_ VPWR VGND sg13g2_and3_1
XFILLER_15_180 VPWR VGND sg13g2_fill_1
XFILLER_16_692 VPWR VGND sg13g2_fill_1
X_5721_ _1518_ VPWR _1646_ VGND net1422 _3480_ sg13g2_o21ai_1
X_5652_ _1567_ _1582_ _1585_ _1589_ VPWR VGND sg13g2_nor3_1
X_4603_ _0636_ net1517 net810 VPWR VGND sg13g2_nand2_1
X_5583_ net1412 net1350 _1520_ VPWR VGND sg13g2_nor2b_1
XFILLER_11_1026 VPWR VGND sg13g2_fill_2
X_4534_ _0137_ _0576_ _0577_ _3420_ net1580 VPWR VGND sg13g2_a22oi_1
X_7322_ net1228 s0.data_out\[2\]\[6\] _3089_ VPWR VGND sg13g2_and2_1
Xhold302 _2972_ VPWR VGND net671 sg13g2_dlygate4sd3_1
Xhold335 s0.shift_out\[9\][0] VPWR VGND net704 sg13g2_dlygate4sd3_1
Xhold313 _1496_ VPWR VGND net682 sg13g2_dlygate4sd3_1
Xhold324 s0.data_out\[5\]\[3\] VPWR VGND net693 sg13g2_dlygate4sd3_1
Xhold368 s0.data_out\[1\]\[6\] VPWR VGND net737 sg13g2_dlygate4sd3_1
Xhold346 s0.was_valid_out\[1\][0] VPWR VGND net715 sg13g2_dlygate4sd3_1
Xhold357 s0.data_out\[14\]\[5\] VPWR VGND net726 sg13g2_dlygate4sd3_1
X_4465_ _0510_ net1528 net601 VPWR VGND sg13g2_nand2_1
X_7253_ VGND VPWR net1228 _3025_ _3027_ _3026_ sg13g2_a21oi_1
Xhold379 s0.was_valid_out\[8\][0] VPWR VGND net748 sg13g2_dlygate4sd3_1
X_6204_ _3383_ VPWR _2084_ VGND net441 net1374 sg13g2_o21ai_1
X_4396_ VGND VPWR _0453_ _0449_ net1668 sg13g2_or2_1
X_7184_ net1191 _3534_ _2966_ VPWR VGND sg13g2_nor2_1
X_6135_ _2024_ net1374 net639 VPWR VGND sg13g2_nand2_1
X_6066_ VPWR _0287_ net739 VGND sg13g2_inv_1
X_5017_ _0895_ VPWR _1015_ VGND net1489 _3447_ sg13g2_o21ai_1
XFILLER_39_784 VPWR VGND sg13g2_fill_2
XFILLER_27_924 VPWR VGND sg13g2_fill_1
X_6968_ _2766_ VPWR _2769_ VGND net1258 _2768_ sg13g2_o21ai_1
XFILLER_35_990 VPWR VGND sg13g2_decap_8
X_6899_ net1265 net1339 _2709_ VPWR VGND sg13g2_nor2b_1
X_5919_ net1402 VPWR _1829_ VGND _1748_ _1828_ sg13g2_o21ai_1
XFILLER_10_813 VPWR VGND sg13g2_fill_2
XFILLER_22_695 VPWR VGND sg13g2_fill_1
XFILLER_5_305 VPWR VGND sg13g2_fill_2
X_7794__223 VPWR VGND net223 sg13g2_tiehi
XFILLER_1_511 VPWR VGND sg13g2_fill_1
XFILLER_45_743 VPWR VGND sg13g2_decap_8
XFILLER_41_982 VPWR VGND sg13g2_decap_8
XFILLER_13_695 VPWR VGND sg13g2_fill_2
XFILLER_34_1026 VPWR VGND sg13g2_fill_2
XFILLER_8_154 VPWR VGND sg13g2_decap_4
XFILLER_5_872 VPWR VGND sg13g2_decap_8
X_4250_ net1647 _3604_ _3614_ VPWR VGND sg13g2_nor2_1
X_4181_ s0.data_out\[27\]\[6\] net1166 _3551_ VPWR VGND sg13g2_nor2_1
X_7940_ net65 VGND VPWR _0074_ s0.genblk1\[27\].modules.bubble clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
XFILLER_48_592 VPWR VGND sg13g2_decap_8
X_7871_ net140 VGND VPWR net650 s0.data_out\[8\]\[1\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_6822_ _2637_ VPWR _2638_ VGND net1729 net712 sg13g2_o21ai_1
XFILLER_17_990 VPWR VGND sg13g2_decap_8
XFILLER_23_437 VPWR VGND sg13g2_fill_1
X_6753_ _2575_ net1280 net630 VPWR VGND sg13g2_nand2_1
X_6684_ net1177 _3516_ _2515_ VPWR VGND sg13g2_nor2_1
X_5704_ _1628_ VPWR _1629_ VGND net1408 _3475_ sg13g2_o21ai_1
XFILLER_32_982 VPWR VGND sg13g2_decap_8
X_7970__93 VPWR VGND net93 sg13g2_tiehi
X_5635_ _1572_ net777 net1433 VPWR VGND sg13g2_nand2b_1
X_5566_ net1623 _1439_ _1507_ VPWR VGND sg13g2_nor2_1
Xhold110 _0152_ VPWR VGND net479 sg13g2_dlygate4sd3_1
X_4517_ net432 VPWR _0562_ VGND net1543 _3428_ sg13g2_o21ai_1
Xhold121 _0155_ VPWR VGND net490 sg13g2_dlygate4sd3_1
X_5497_ VGND VPWR _1318_ _1445_ _1446_ net1440 sg13g2_a21oi_1
Xhold132 s0.data_out\[25\]\[3\] VPWR VGND net501 sg13g2_dlygate4sd3_1
Xhold143 _1040_ VPWR VGND net512 sg13g2_dlygate4sd3_1
X_7305_ VGND VPWR net1234 s0.data_out\[2\]\[2\] _3076_ _3007_ sg13g2_a21oi_1
X_4448_ net1727 net374 _0135_ VPWR VGND sg13g2_and2_1
Xhold165 s0.data_out\[21\]\[3\] VPWR VGND net534 sg13g2_dlygate4sd3_1
X_7236_ s0.data_out\[2\]\[2\] s0.data_out\[3\]\[2\] net1247 _3010_ VPWR VGND sg13g2_mux2_1
Xhold154 s0.data_out\[10\]\[2\] VPWR VGND net523 sg13g2_dlygate4sd3_1
Xhold176 _2292_ VPWR VGND net545 sg13g2_dlygate4sd3_1
Xhold187 s0.data_out\[25\]\[7\] VPWR VGND net556 sg13g2_dlygate4sd3_1
Xhold198 _0047_ VPWR VGND net567 sg13g2_dlygate4sd3_1
X_4379_ _0436_ net1542 s0.data_out\[25\]\[4\] VPWR VGND sg13g2_nand2_1
X_7167_ net384 net1565 _2953_ VPWR VGND sg13g2_nor2_1
X_6118_ s0.data_out\[12\]\[6\] s0.data_out\[11\]\[6\] net1374 _2007_ VPWR VGND sg13g2_mux2_1
X_7098_ s0.data_out\[4\]\[1\] s0.data_out\[3\]\[1\] net1246 _2884_ VPWR VGND sg13g2_mux2_1
X_6049_ VPWR _0283_ net625 VGND sg13g2_inv_1
XFILLER_37_68 VPWR VGND sg13g2_fill_2
XFILLER_27_765 VPWR VGND sg13g2_fill_2
XFILLER_42_724 VPWR VGND sg13g2_fill_1
X_7938__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_14_459 VPWR VGND sg13g2_fill_1
X_7902__107 VPWR VGND net107 sg13g2_tiehi
XFILLER_2_875 VPWR VGND sg13g2_decap_8
XFILLER_17_242 VPWR VGND sg13g2_fill_1
XFILLER_45_584 VPWR VGND sg13g2_decap_4
XFILLER_17_297 VPWR VGND sg13g2_fill_2
X_5420_ net1439 net681 _1376_ VPWR VGND sg13g2_and2_1
X_5351_ _1310_ net1438 _1311_ _1312_ VPWR VGND sg13g2_a21o_1
X_4302_ _0117_ _0364_ _0365_ _3408_ net1575 VPWR VGND sg13g2_a22oi_1
X_5282_ _1253_ VPWR _1254_ VGND net1737 net647 sg13g2_o21ai_1
X_4233_ net515 net1563 _3597_ VPWR VGND sg13g2_nor2b_1
X_7021_ _2816_ _2817_ _2819_ VPWR VGND _2818_ sg13g2_nand3b_1
X_4164_ VPWR _3540_ net735 VGND sg13g2_inv_1
X_4095_ VPWR _3471_ net495 VGND sg13g2_inv_1
X_7923_ net84 VGND VPWR _0057_ s0.data_out\[4\]\[5\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_7964__178 VPWR VGND net178 sg13g2_tiehi
X_7854_ net159 VGND VPWR net456 s0.was_valid_out\[9\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_6805_ _0017_ _2623_ _2624_ _3514_ net1598 VPWR VGND sg13g2_a22oi_1
X_7785_ net233 VGND VPWR _0263_ s0.data_out\[15\]\[6\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4997_ _0995_ net835 net1489 VPWR VGND sg13g2_nand2b_1
X_6736_ s0.data_out\[7\]\[0\] s0.data_out\[6\]\[0\] net1278 _2558_ VPWR VGND sg13g2_mux2_1
XFILLER_23_59 VPWR VGND sg13g2_fill_1
X_6667_ _2498_ _2499_ _2500_ _2501_ VPWR VGND sg13g2_nor3_1
X_6598_ _2433_ _2434_ _0000_ VPWR VGND sg13g2_nor2_1
X_5618_ VGND VPWR _1434_ _1554_ _1555_ net1428 sg13g2_a21oi_1
X_5549_ VGND VPWR net1426 s0.data_out\[16\]\[4\] _1493_ _1461_ sg13g2_a21oi_1
X_7791__226 VPWR VGND net226 sg13g2_tiehi
Xfanout1429 net1430 net1429 VPWR VGND sg13g2_buf_2
X_7219_ s0.data_out\[3\]\[1\] s0.data_out\[2\]\[1\] net1235 _2993_ VPWR VGND sg13g2_mux2_1
Xfanout1418 net468 net1418 VPWR VGND sg13g2_buf_8
Xfanout1407 net474 net1407 VPWR VGND sg13g2_buf_8
XFILLER_48_67 VPWR VGND sg13g2_fill_2
XFILLER_24_1014 VPWR VGND sg13g2_decap_8
XFILLER_42_510 VPWR VGND sg13g2_fill_1
XFILLER_14_223 VPWR VGND sg13g2_fill_1
XFILLER_10_473 VPWR VGND sg13g2_fill_2
XFILLER_2_694 VPWR VGND sg13g2_fill_2
XFILLER_1_160 VPWR VGND sg13g2_fill_1
XFILLER_45_381 VPWR VGND sg13g2_fill_2
X_4920_ net1605 _0863_ _0925_ VPWR VGND sg13g2_nor2_1
X_4851_ _0859_ VPWR _0860_ VGND net1491 _3439_ sg13g2_o21ai_1
XFILLER_33_532 VPWR VGND sg13g2_fill_1
XFILLER_21_738 VPWR VGND sg13g2_fill_2
X_7570_ VGND VPWR net1210 net447 _3312_ _3246_ sg13g2_a21oi_1
X_4782_ net1514 VPWR _0801_ VGND _0720_ _0800_ sg13g2_o21ai_1
X_6521_ net1667 _2364_ _2367_ VPWR VGND sg13g2_nor2_1
XFILLER_9_260 VPWR VGND sg13g2_decap_4
X_7925__82 VPWR VGND net82 sg13g2_tiehi
X_6452_ _2302_ net1738 _2303_ VPWR VGND _2249_ sg13g2_nand3b_1
X_5403_ _1362_ VPWR _1363_ VGND net1203 _1361_ sg13g2_o21ai_1
X_6383_ _2241_ net483 net1362 VPWR VGND sg13g2_nand2b_1
XFILLER_47_1025 VPWR VGND sg13g2_decap_4
X_5334_ VGND VPWR net1436 _1293_ _1295_ _1294_ sg13g2_a21oi_1
X_5265_ _1237_ net1449 _1235_ _1238_ VPWR VGND sg13g2_a21o_1
X_5196_ net1448 _1169_ _1172_ VPWR VGND sg13g2_nor2_1
X_4216_ net1546 net1356 _3580_ VPWR VGND sg13g2_nor2b_1
X_7004_ _2802_ net1253 net780 VPWR VGND sg13g2_nand2_1
X_4147_ VPWR _3523_ net694 VGND sg13g2_inv_1
X_4078_ VPWR _3454_ net814 VGND sg13g2_inv_1
XFILLER_43_318 VPWR VGND sg13g2_fill_1
X_7906_ net102 VGND VPWR _0040_ s0.data_out\[5\]\[0\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_7837_ net176 VGND VPWR _0315_ s0.data_new_delayed\[0\] clknet_leaf_7_clk sg13g2_dfrbpq_2
XFILLER_12_716 VPWR VGND sg13g2_fill_1
X_7768_ net251 VGND VPWR net496 s0.data_out\[16\]\[1\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_6719_ net1601 _2536_ _0013_ VPWR VGND sg13g2_nor2_1
X_7699_ net326 VGND VPWR _0177_ s0.data_out\[22\]\[4\] clknet_leaf_40_clk sg13g2_dfrbpq_2
Xclkload2 clknet_3_7__leaf_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_20_782 VPWR VGND sg13g2_decap_4
XFILLER_4_948 VPWR VGND sg13g2_decap_8
Xfanout1204 net1205 net1204 VPWR VGND sg13g2_buf_1
Xfanout1215 net1216 net1215 VPWR VGND sg13g2_buf_8
Xfanout1226 net1227 net1226 VPWR VGND sg13g2_buf_8
Xfanout1237 net1238 net1237 VPWR VGND sg13g2_buf_8
Xfanout1248 net1249 net1248 VPWR VGND sg13g2_buf_8
Xfanout1259 net480 net1259 VPWR VGND sg13g2_buf_8
XFILLER_47_668 VPWR VGND sg13g2_decap_8
XFILLER_46_167 VPWR VGND sg13g2_fill_1
XFILLER_27_370 VPWR VGND sg13g2_fill_1
X_7922__85 VPWR VGND net85 sg13g2_tiehi
XFILLER_3_970 VPWR VGND sg13g2_decap_8
X_5050_ _0187_ _1042_ _1043_ _3443_ net1605 VPWR VGND sg13g2_a22oi_1
X_4001_ VPWR _3377_ net1451 VGND sg13g2_inv_1
XFILLER_1_40 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_22 VPWR VGND uio_out[6] sg13g2_tielo
Xheichips25_top_sorter_11 VPWR VGND uio_oe[0] sg13g2_tielo
X_5952_ _1856_ _1853_ _1855_ VPWR VGND sg13g2_nand2_1
X_4903_ VGND VPWR _0907_ _0910_ _0172_ _0911_ sg13g2_a21oi_1
XFILLER_18_392 VPWR VGND sg13g2_fill_2
X_5883_ _1793_ _1794_ _1792_ _1796_ VPWR VGND sg13g2_nand3_1
X_7622_ VGND VPWR net1722 _3340_ _0103_ _3355_ sg13g2_a21oi_1
X_4834_ _0843_ net1491 s0.data_out\[21\]\[1\] VPWR VGND sg13g2_nand2_1
X_7553_ _3298_ VPWR _3299_ VGND net1722 net614 sg13g2_o21ai_1
X_4765_ _0786_ _0778_ _0785_ VPWR VGND sg13g2_nand2_1
XFILLER_14_1002 VPWR VGND sg13g2_decap_8
X_6504_ VPWR VGND net1691 _2342_ _2349_ net1699 _2350_ _2325_ sg13g2_a221oi_1
X_7484_ VPWR VGND _3232_ net1710 _3228_ net1702 _3234_ _3226_ sg13g2_a221oi_1
X_4696_ net1727 net385 _0159_ VPWR VGND sg13g2_and2_1
X_6435_ net1608 _2210_ _2290_ VPWR VGND sg13g2_nor2_1
X_6366_ s0.data_out\[9\]\[0\] s0.data_out\[10\]\[0\] net1360 _2224_ VPWR VGND sg13g2_mux2_1
X_5317_ VGND VPWR _1281_ net1444 net428 sg13g2_or2_1
XFILLER_0_417 VPWR VGND sg13g2_decap_8
XFILLER_0_428 VPWR VGND sg13g2_fill_2
XFILLER_1_929 VPWR VGND sg13g2_decap_8
Xhold14 s0.genblk1\[7\].modules.bubble VPWR VGND net383 sg13g2_dlygate4sd3_1
X_6297_ _0307_ _2169_ _2170_ _3494_ net1611 VPWR VGND sg13g2_a22oi_1
Xhold25 s0.genblk1\[9\].modules.bubble VPWR VGND net394 sg13g2_dlygate4sd3_1
Xhold47 s0.was_valid_out\[13\][0] VPWR VGND net416 sg13g2_dlygate4sd3_1
X_5248_ VGND VPWR _1107_ _1220_ _1221_ net1461 sg13g2_a21oi_1
Xhold36 s0.was_valid_out\[15\][0] VPWR VGND net405 sg13g2_dlygate4sd3_1
Xhold58 _2495_ VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold69 _0205_ VPWR VGND net438 sg13g2_dlygate4sd3_1
X_5179_ _0201_ _1157_ _1158_ _3447_ net1606 VPWR VGND sg13g2_a22oi_1
XFILLER_21_1028 VPWR VGND sg13g2_fill_1
XFILLER_16_318 VPWR VGND sg13g2_fill_1
XFILLER_12_502 VPWR VGND sg13g2_fill_2
XFILLER_3_288 VPWR VGND sg13g2_fill_2
XFILLER_48_900 VPWR VGND sg13g2_decap_8
XFILLER_48_977 VPWR VGND sg13g2_decap_8
XFILLER_16_830 VPWR VGND sg13g2_fill_1
XFILLER_37_1024 VPWR VGND sg13g2_decap_4
X_4550_ _0589_ VPWR _0590_ VGND net1184 _0588_ sg13g2_o21ai_1
X_4481_ net1687 _0525_ _0526_ VPWR VGND sg13g2_nor2_1
X_6220_ net1321 net1354 _2097_ VPWR VGND sg13g2_nor2b_1
X_6151_ _2039_ _2037_ net1684 _2040_ VPWR VGND sg13g2_a21o_1
X_5102_ s0.data_out\[19\]\[0\] s0.data_out\[20\]\[0\] net1479 _1087_ VPWR VGND sg13g2_mux2_1
X_6082_ _1968_ _1973_ _0289_ VPWR VGND sg13g2_nor2_1
X_7713__311 VPWR VGND net311 sg13g2_tiehi
XFILLER_25_0 VPWR VGND sg13g2_fill_2
X_5033_ VGND VPWR net1179 _0969_ _1030_ net1607 sg13g2_a21oi_1
XFILLER_38_432 VPWR VGND sg13g2_decap_8
Xfanout1590 net1591 net1590 VPWR VGND sg13g2_buf_8
XFILLER_39_999 VPWR VGND sg13g2_decap_8
X_6984_ _2782_ net716 net1266 VPWR VGND sg13g2_nand2b_1
XFILLER_25_137 VPWR VGND sg13g2_fill_1
X_5935_ net1395 s0.data_out\[13\]\[6\] _1841_ VPWR VGND sg13g2_and2_1
XFILLER_15_27 VPWR VGND sg13g2_fill_1
X_5866_ s0.data_out\[14\]\[7\] s0.data_out\[13\]\[7\] net1399 _1779_ VPWR VGND sg13g2_mux2_1
X_7605_ _3342_ VPWR _3343_ VGND _3393_ net1343 sg13g2_o21ai_1
X_4817_ _0826_ VPWR _0829_ VGND net412 net1490 sg13g2_o21ai_1
XFILLER_22_899 VPWR VGND sg13g2_decap_4
X_5797_ VPWR _0259_ net607 VGND sg13g2_inv_1
X_7536_ net1208 net570 _3285_ VPWR VGND sg13g2_and2_1
X_4748_ net1650 _0759_ _0769_ VPWR VGND sg13g2_nor2_1
X_7467_ net1212 net1348 _3217_ VPWR VGND sg13g2_nor2b_1
X_4679_ net1523 VPWR _0705_ VGND _0653_ _0704_ sg13g2_o21ai_1
X_6418_ _2271_ VPWR _2276_ VGND _2262_ _2270_ sg13g2_o21ai_1
XFILLER_1_726 VPWR VGND sg13g2_decap_8
X_7398_ _3159_ VPWR _3160_ VGND net1188 _3157_ sg13g2_o21ai_1
X_6349_ net1307 net1351 _2207_ VPWR VGND sg13g2_nor2b_1
X_7833__181 VPWR VGND net181 sg13g2_tiehi
XFILLER_5_1000 VPWR VGND sg13g2_decap_8
XFILLER_45_914 VPWR VGND sg13g2_decap_8
XFILLER_17_616 VPWR VGND sg13g2_fill_2
XFILLER_31_107 VPWR VGND sg13g2_fill_1
XFILLER_48_774 VPWR VGND sg13g2_decap_8
XFILLER_36_947 VPWR VGND sg13g2_fill_2
XFILLER_36_958 VPWR VGND sg13g2_decap_8
XFILLER_23_608 VPWR VGND sg13g2_fill_2
X_5720_ VGND VPWR net1403 _1643_ _1645_ _1644_ sg13g2_a21oi_1
Xclkbuf_leaf_42_clk clknet_3_1__leaf_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
XFILLER_31_630 VPWR VGND sg13g2_fill_1
X_5651_ _1549_ _1567_ _1587_ _1588_ VPWR VGND sg13g2_or3_1
XFILLER_11_1005 VPWR VGND sg13g2_decap_8
X_4602_ _0619_ _0633_ _0634_ _0635_ VPWR VGND sg13g2_nor3_1
X_5582_ s0.data_out\[16\]\[2\] s0.data_out\[15\]\[2\] net1419 _1519_ VPWR VGND sg13g2_mux2_1
XFILLER_8_870 VPWR VGND sg13g2_fill_1
X_4533_ VGND VPWR net1185 _0501_ _0577_ net1580 sg13g2_a21oi_1
X_7321_ _0069_ _3087_ _3088_ _3536_ net1586 VPWR VGND sg13g2_a22oi_1
Xhold303 s0.data_out\[19\]\[7\] VPWR VGND net672 sg13g2_dlygate4sd3_1
Xhold314 s0.data_out\[21\]\[0\] VPWR VGND net683 sg13g2_dlygate4sd3_1
Xhold325 s0.data_out\[6\]\[1\] VPWR VGND net694 sg13g2_dlygate4sd3_1
X_7252_ net1228 net1334 _3026_ VPWR VGND sg13g2_nor2b_1
Xhold358 s0.data_out\[1\]\[7\] VPWR VGND net727 sg13g2_dlygate4sd3_1
Xhold369 s0.data_out\[13\]\[6\] VPWR VGND net738 sg13g2_dlygate4sd3_1
X_6203_ net1325 _2077_ _2083_ VPWR VGND sg13g2_nor2_1
X_4464_ net1522 net1348 _0509_ VPWR VGND sg13g2_nor2b_1
Xhold336 s0.data_out\[17\]\[2\] VPWR VGND net705 sg13g2_dlygate4sd3_1
Xhold347 s0.data_out\[4\]\[1\] VPWR VGND net716 sg13g2_dlygate4sd3_1
X_4395_ net1687 _0414_ _0452_ VPWR VGND sg13g2_nor2_1
X_7183_ VPWR _0054_ net686 VGND sg13g2_inv_1
X_6134_ _2022_ _2020_ _2023_ VPWR VGND _2021_ sg13g2_nand3b_1
X_7817__198 VPWR VGND net198 sg13g2_tiehi
X_6065_ _1958_ VPWR _1959_ VGND net1747 net738 sg13g2_o21ai_1
XFILLER_39_730 VPWR VGND sg13g2_decap_8
X_5016_ _1014_ net1484 _1013_ VPWR VGND sg13g2_nand2b_1
X_7967__132 VPWR VGND net132 sg13g2_tiehi
X_7787__231 VPWR VGND net231 sg13g2_tiehi
XFILLER_14_619 VPWR VGND sg13g2_fill_2
X_6967_ net400 net1267 _2768_ VPWR VGND sg13g2_nor2_1
X_5918_ net1193 _3486_ _1828_ VPWR VGND sg13g2_nor2_1
X_6898_ s0.data_out\[6\]\[5\] s0.data_out\[5\]\[5\] net1268 _2708_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_33_clk clknet_3_5__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
XFILLER_42_58 VPWR VGND sg13g2_fill_2
XFILLER_21_162 VPWR VGND sg13g2_fill_2
XFILLER_22_685 VPWR VGND sg13g2_fill_1
X_5849_ net1390 net1359 _1762_ VPWR VGND sg13g2_nor2b_1
X_7519_ _3269_ net1200 _3268_ VPWR VGND sg13g2_nand2_1
XFILLER_49_549 VPWR VGND sg13g2_decap_8
XFILLER_45_700 VPWR VGND sg13g2_decap_8
XFILLER_26_991 VPWR VGND sg13g2_decap_8
XFILLER_32_427 VPWR VGND sg13g2_decap_4
XFILLER_41_961 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_24_clk clknet_3_7__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_34_1005 VPWR VGND sg13g2_decap_8
XFILLER_9_612 VPWR VGND sg13g2_fill_1
XFILLER_9_678 VPWR VGND sg13g2_fill_2
X_4180_ VGND VPWR _3403_ net1166 net8 _3550_ sg13g2_a21oi_1
XFILLER_48_571 VPWR VGND sg13g2_decap_8
X_7710__314 VPWR VGND net314 sg13g2_tiehi
X_7870_ net141 VGND VPWR _0004_ s0.data_out\[8\]\[0\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_6821_ _2636_ VPWR _2637_ VGND net1176 _2635_ sg13g2_o21ai_1
X_7947__58 VPWR VGND net58 sg13g2_tiehi
XFILLER_24_917 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_15_clk clknet_3_3__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_6752_ _2573_ VPWR _2574_ VGND _2564_ _2565_ sg13g2_o21ai_1
X_6683_ _0005_ _2513_ _2514_ _3513_ net1599 VPWR VGND sg13g2_a22oi_1
X_5703_ _1628_ net1408 net603 VPWR VGND sg13g2_nand2_1
X_5634_ _1569_ net1415 _1570_ _1571_ VPWR VGND sg13g2_a21o_1
Xhold100 s0.data_out\[27\]\[4\] VPWR VGND net469 sg13g2_dlygate4sd3_1
X_5565_ net1441 VPWR _1506_ VGND _1436_ _1505_ sg13g2_o21ai_1
X_7304_ VPWR _0065_ _3075_ VGND sg13g2_inv_1
Xhold122 s0.data_out\[26\]\[5\] VPWR VGND net491 sg13g2_dlygate4sd3_1
X_4516_ _0561_ net1537 _0560_ VPWR VGND sg13g2_nand2b_1
Xhold133 _0128_ VPWR VGND net502 sg13g2_dlygate4sd3_1
X_5496_ _1445_ s0.data_out\[16\]\[6\] net1444 VPWR VGND sg13g2_nand2b_1
Xhold144 s0.data_out\[12\]\[1\] VPWR VGND net513 sg13g2_dlygate4sd3_1
Xhold111 s0.shift_out\[5\][0] VPWR VGND net480 sg13g2_dlygate4sd3_1
Xhold155 s0.was_valid_out\[26\][0] VPWR VGND net524 sg13g2_dlygate4sd3_1
X_4447_ net1716 _0488_ _0134_ VPWR VGND sg13g2_and2_1
Xhold166 _0187_ VPWR VGND net535 sg13g2_dlygate4sd3_1
X_7235_ net1191 _3008_ _3009_ VPWR VGND sg13g2_nor2_1
Xhold177 _0327_ VPWR VGND net546 sg13g2_dlygate4sd3_1
Xhold188 s0.data_out\[26\]\[7\] VPWR VGND net557 sg13g2_dlygate4sd3_1
X_7166_ _2951_ VPWR _2952_ VGND _2929_ _2948_ sg13g2_o21ai_1
Xhold199 s0.data_out\[2\]\[7\] VPWR VGND net568 sg13g2_dlygate4sd3_1
X_6117_ _2006_ net1374 net687 VPWR VGND sg13g2_nand2_1
X_4378_ _0434_ _0431_ _0435_ VPWR VGND _0432_ sg13g2_nand3b_1
X_7097_ _2882_ VPWR _2883_ VGND net1171 _2880_ sg13g2_o21ai_1
X_6048_ _1945_ VPWR _1946_ VGND net1747 net624 sg13g2_o21ai_1
X_7830__184 VPWR VGND net184 sg13g2_tiehi
XFILLER_15_917 VPWR VGND sg13g2_fill_1
XFILLER_14_416 VPWR VGND sg13g2_fill_1
XFILLER_6_659 VPWR VGND sg13g2_fill_1
XFILLER_5_158 VPWR VGND sg13g2_fill_1
XFILLER_2_854 VPWR VGND sg13g2_decap_8
XFILLER_18_788 VPWR VGND sg13g2_fill_2
XFILLER_27_80 VPWR VGND sg13g2_fill_1
XFILLER_20_408 VPWR VGND sg13g2_decap_4
XFILLER_9_442 VPWR VGND sg13g2_fill_1
X_7777__241 VPWR VGND net241 sg13g2_tiehi
X_5350_ net1438 net1347 _1311_ VPWR VGND sg13g2_nor2b_1
X_4301_ net1575 _3628_ _0365_ VPWR VGND sg13g2_nor2_1
X_5281_ _1252_ VPWR _1253_ VGND net1199 _1251_ sg13g2_o21ai_1
X_4232_ VPWR _3596_ _3595_ VGND sg13g2_inv_1
X_7020_ net1650 _2808_ _2818_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_4_clk clknet_3_1__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ VPWR _3539_ net520 VGND sg13g2_inv_1
X_4094_ VPWR _3470_ net655 VGND sg13g2_inv_1
X_7922_ net85 VGND VPWR _0056_ s0.data_out\[4\]\[4\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_7784__234 VPWR VGND net234 sg13g2_tiehi
X_7853_ net160 VGND VPWR _0331_ s0.data_out\[10\]\[7\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_4996_ _0992_ net1469 _0993_ _0994_ VPWR VGND sg13g2_a21o_1
XFILLER_24_769 VPWR VGND sg13g2_fill_1
X_6804_ net1598 _2556_ _2624_ VPWR VGND sg13g2_nor2_1
X_7784_ net234 VGND VPWR _0262_ s0.data_out\[15\]\[5\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_17_1011 VPWR VGND sg13g2_decap_8
X_6735_ VGND VPWR net1282 _2554_ _2557_ _2556_ sg13g2_a21oi_1
X_6666_ net1691 _2465_ _2500_ VPWR VGND sg13g2_nor2_1
X_6597_ net1731 VPWR _2434_ VGND net748 _2428_ sg13g2_o21ai_1
X_5617_ _1554_ s0.data_out\[15\]\[7\] net1434 VPWR VGND sg13g2_nand2b_1
X_5548_ _0236_ _1491_ _1492_ _3463_ net1622 VPWR VGND sg13g2_a22oi_1
XFILLER_2_106 VPWR VGND sg13g2_fill_2
X_5479_ VGND VPWR _1309_ _1427_ _1428_ net1438 sg13g2_a21oi_1
X_7218_ _2992_ net1236 s0.data_out\[2\]\[1\] VPWR VGND sg13g2_nand2_1
Xfanout1419 net1422 net1419 VPWR VGND sg13g2_buf_8
Xfanout1408 net1409 net1408 VPWR VGND sg13g2_buf_8
X_7149_ VGND VPWR _2802_ _2934_ _2935_ net1248 sg13g2_a21oi_1
XFILLER_19_508 VPWR VGND sg13g2_fill_1
XFILLER_42_555 VPWR VGND sg13g2_fill_2
XFILLER_14_257 VPWR VGND sg13g2_decap_8
X_7934__72 VPWR VGND net72 sg13g2_tiehi
XFILLER_6_401 VPWR VGND sg13g2_fill_2
XFILLER_9_1009 VPWR VGND sg13g2_decap_8
XFILLER_37_327 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_46_883 VPWR VGND sg13g2_decap_8
X_4850_ _0859_ net1491 net534 VPWR VGND sg13g2_nand2_1
XFILLER_33_566 VPWR VGND sg13g2_fill_1
X_6520_ VGND VPWR _2366_ _2357_ net1657 sg13g2_or2_1
X_4781_ net1495 net599 _0800_ VPWR VGND sg13g2_and2_1
X_6451_ net1323 VPWR _2302_ VGND _2246_ _2301_ sg13g2_o21ai_1
X_6382_ _2238_ net1311 _2239_ _2240_ VPWR VGND sg13g2_a21o_1
X_5402_ VGND VPWR net1203 _1303_ _1362_ net1619 sg13g2_a21oi_1
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
X_5333_ net1436 net1354 _1294_ VPWR VGND sg13g2_nor2b_1
X_5264_ s0.data_out\[19\]\[4\] s0.data_out\[18\]\[4\] net1453 _1237_ VPWR VGND sg13g2_mux2_1
X_5195_ _1170_ VPWR _1171_ VGND s0.was_valid_out\[18\][0] net1453 sg13g2_o21ai_1
X_4215_ VGND VPWR net1564 _3419_ _3579_ _3578_ sg13g2_a21oi_1
X_7003_ _2800_ VPWR _2801_ VGND _2791_ _2792_ sg13g2_o21ai_1
X_4146_ VPWR _3522_ net532 VGND sg13g2_inv_1
XFILLER_29_806 VPWR VGND sg13g2_fill_2
XFILLER_29_828 VPWR VGND sg13g2_fill_1
X_4077_ VPWR _3453_ net435 VGND sg13g2_inv_1
XFILLER_24_500 VPWR VGND sg13g2_fill_1
X_7905_ net103 VGND VPWR _0039_ s0.shift_out\[5\][0] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_7836_ net177 VGND VPWR _0314_ s0.valid_out\[10\][0] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_11_216 VPWR VGND sg13g2_fill_1
X_4979_ _0975_ net1471 _0976_ _0977_ VPWR VGND sg13g2_a21o_1
X_7767_ net252 VGND VPWR _0245_ s0.data_out\[16\]\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_2
XFILLER_24_599 VPWR VGND sg13g2_fill_2
X_6718_ _2537_ _2542_ _0012_ VPWR VGND sg13g2_nor2_1
X_7698_ net327 VGND VPWR net531 s0.data_out\[22\]\[3\] clknet_leaf_40_clk sg13g2_dfrbpq_2
Xclkload3 VPWR clkload3/Y clknet_leaf_2_clk VGND sg13g2_inv_1
X_6649_ VGND VPWR _2483_ _2480_ net1651 sg13g2_or2_1
X_7931__75 VPWR VGND net75 sg13g2_tiehi
XFILLER_4_927 VPWR VGND sg13g2_decap_8
Xfanout1205 _3377_ net1205 VPWR VGND sg13g2_buf_1
Xfanout1216 net571 net1216 VPWR VGND sg13g2_buf_8
Xfanout1227 s0.valid_out\[1\][0] net1227 VPWR VGND sg13g2_buf_8
Xfanout1238 s0.valid_out\[2\][0] net1238 VPWR VGND sg13g2_buf_2
Xfanout1249 net454 net1249 VPWR VGND sg13g2_buf_8
XFILLER_28_861 VPWR VGND sg13g2_fill_2
XFILLER_43_886 VPWR VGND sg13g2_fill_1
XFILLER_11_761 VPWR VGND sg13g2_fill_2
X_4000_ VPWR _3376_ net1434 VGND sg13g2_inv_1
Xfanout1750 net1751 net1750 VPWR VGND sg13g2_buf_8
XFILLER_37_124 VPWR VGND sg13g2_fill_1
XFILLER_38_658 VPWR VGND sg13g2_fill_1
Xheichips25_top_sorter_23 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_19_861 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_12 VPWR VGND uio_oe[1] sg13g2_tielo
X_5951_ net1194 VPWR _1855_ VGND s0.was_valid_out\[12\][0] net1398 sg13g2_o21ai_1
X_4902_ VGND VPWR _0911_ net1567 net385 sg13g2_or2_1
XFILLER_18_382 VPWR VGND sg13g2_fill_1
X_5882_ _1795_ _1792_ _1793_ _1794_ VPWR VGND sg13g2_and3_1
X_7781__237 VPWR VGND net237 sg13g2_tiehi
X_7621_ net1722 net433 _3355_ VPWR VGND sg13g2_nor2_1
X_4833_ _0840_ _0838_ net1699 _0842_ VPWR VGND sg13g2_a21o_1
X_7552_ _3297_ VPWR _3298_ VGND net1200 _3296_ sg13g2_o21ai_1
X_4764_ _0782_ _0784_ net1679 _0785_ VPWR VGND sg13g2_nand3_1
X_7483_ VGND VPWR _3233_ _3226_ net1702 sg13g2_or2_1
X_6503_ VGND VPWR net1306 _2346_ _2349_ _2348_ sg13g2_a21oi_1
X_4695_ net1727 _0712_ _0158_ VPWR VGND sg13g2_and2_1
X_6434_ net1319 VPWR _2289_ VGND _2207_ _2288_ sg13g2_o21ai_1
XFILLER_1_908 VPWR VGND sg13g2_decap_8
X_6365_ _2223_ net1319 _2222_ VPWR VGND sg13g2_nand2b_1
X_5316_ net821 _1278_ net476 _1280_ VPWR VGND sg13g2_nor3_1
X_6296_ net1611 _2092_ _2170_ VPWR VGND sg13g2_nor2_1
X_5247_ _1220_ s0.data_out\[18\]\[7\] net1466 VPWR VGND sg13g2_nand2b_1
Xhold26 s0.genblk1\[14\].modules.bubble VPWR VGND net395 sg13g2_dlygate4sd3_1
Xhold15 s0.genblk1\[4\].modules.bubble VPWR VGND net384 sg13g2_dlygate4sd3_1
XFILLER_29_37 VPWR VGND sg13g2_fill_2
Xhold37 _0253_ VPWR VGND net406 sg13g2_dlygate4sd3_1
Xhold48 _0277_ VPWR VGND net417 sg13g2_dlygate4sd3_1
X_5178_ net1606 net436 _1158_ VPWR VGND sg13g2_nor2_1
Xhold59 s0.was_valid_out\[17\][0] VPWR VGND net428 sg13g2_dlygate4sd3_1
XFILLER_28_102 VPWR VGND sg13g2_fill_2
XFILLER_29_669 VPWR VGND sg13g2_fill_2
X_4129_ VPWR _3505_ net485 VGND sg13g2_inv_1
X_7819_ net196 VGND VPWR _0297_ s0.data_out\[12\]\[4\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_0_985 VPWR VGND sg13g2_decap_8
XFILLER_48_956 VPWR VGND sg13g2_decap_8
XFILLER_35_606 VPWR VGND sg13g2_fill_1
XFILLER_37_1003 VPWR VGND sg13g2_decap_8
XFILLER_31_812 VPWR VGND sg13g2_fill_1
XFILLER_43_694 VPWR VGND sg13g2_fill_1
XFILLER_7_551 VPWR VGND sg13g2_decap_4
XFILLER_7_540 VPWR VGND sg13g2_fill_1
X_4480_ VGND VPWR net1538 _0522_ _0525_ _0524_ sg13g2_a21oi_1
X_6150_ _2039_ _2038_ net1380 VPWR VGND sg13g2_nand2b_1
X_5101_ _1086_ net1475 _1085_ VPWR VGND sg13g2_nand2b_1
X_6081_ net1739 VPWR _1973_ VGND _1970_ _1972_ sg13g2_o21ai_1
X_5032_ VGND VPWR net1470 s0.data_out\[20\]\[0\] _1029_ _0967_ sg13g2_a21oi_1
XFILLER_39_978 VPWR VGND sg13g2_decap_8
XFILLER_38_455 VPWR VGND sg13g2_decap_4
Xfanout1580 net1588 net1580 VPWR VGND sg13g2_buf_8
Xfanout1591 net1592 net1591 VPWR VGND sg13g2_buf_2
X_6983_ _2779_ net1250 _2780_ _2781_ VPWR VGND sg13g2_a21o_1
X_5934_ _0274_ _1839_ _1840_ _3477_ net1629 VPWR VGND sg13g2_a22oi_1
X_5865_ _1778_ net1399 net575 VPWR VGND sg13g2_nand2_1
XFILLER_22_823 VPWR VGND sg13g2_fill_1
X_7604_ net434 net1216 net1212 _3342_ VPWR VGND sg13g2_a21o_1
X_4816_ _0826_ _0827_ _0828_ VPWR VGND sg13g2_nor2_1
XFILLER_22_856 VPWR VGND sg13g2_fill_2
XFILLER_22_889 VPWR VGND sg13g2_decap_8
X_5796_ _1717_ VPWR _1718_ VGND net1747 net606 sg13g2_o21ai_1
X_7535_ VGND VPWR _3279_ _3283_ _0087_ _3284_ sg13g2_a21oi_1
X_4747_ VGND VPWR _0768_ _0766_ net1660 sg13g2_or2_1
X_7466_ s0.data_out\[1\]\[2\] s0.data_out\[0\]\[2\] net1215 _3216_ VPWR VGND sg13g2_mux2_1
X_4678_ net1181 _3433_ _0704_ VPWR VGND sg13g2_nor2_1
X_6417_ _2262_ _2272_ _2236_ _2275_ VPWR VGND _2274_ sg13g2_nand4_1
X_7397_ _3159_ net1188 _3158_ VPWR VGND sg13g2_nand2_1
X_6348_ s0.data_out\[10\]\[2\] s0.data_out\[9\]\[2\] net1315 _2206_ VPWR VGND sg13g2_mux2_1
X_6279_ _2137_ _2152_ _2154_ _2155_ _2156_ VPWR VGND sg13g2_nor4_1
XFILLER_0_259 VPWR VGND sg13g2_fill_2
XFILLER_31_119 VPWR VGND sg13g2_fill_1
XFILLER_21_71 VPWR VGND sg13g2_fill_2
XFILLER_0_782 VPWR VGND sg13g2_decap_8
XFILLER_48_753 VPWR VGND sg13g2_decap_8
XFILLER_44_981 VPWR VGND sg13g2_decap_8
X_5650_ _1587_ _1582_ _1586_ VPWR VGND sg13g2_nand2_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_4601_ VPWR VGND _0632_ net1710 _0630_ net1703 _0634_ _0626_ sg13g2_a221oi_1
X_5581_ _1518_ net1419 s0.data_out\[15\]\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
X_4532_ net1539 VPWR _0576_ VGND _0503_ _0575_ sg13g2_o21ai_1
X_7320_ net1585 _3047_ _3088_ VPWR VGND sg13g2_nor2_1
Xhold304 _0216_ VPWR VGND net673 sg13g2_dlygate4sd3_1
X_4463_ VPWR VGND _0507_ net1710 _0502_ net1703 _0508_ _0500_ sg13g2_a221oi_1
Xhold315 _1032_ VPWR VGND net684 sg13g2_dlygate4sd3_1
Xhold326 _0029_ VPWR VGND net695 sg13g2_dlygate4sd3_1
X_7251_ s0.data_out\[3\]\[6\] s0.data_out\[2\]\[6\] net1235 _3025_ VPWR VGND sg13g2_mux2_1
Xhold359 _3315_ VPWR VGND net728 sg13g2_dlygate4sd3_1
X_6202_ net441 net1363 _2082_ VPWR VGND sg13g2_nor2_1
Xhold337 s0.data_out\[26\]\[6\] VPWR VGND net706 sg13g2_dlygate4sd3_1
Xhold348 _2961_ VPWR VGND net717 sg13g2_dlygate4sd3_1
X_4394_ VPWR _0451_ _0450_ VGND sg13g2_inv_1
X_7182_ _2964_ VPWR _2965_ VGND net1716 net685 sg13g2_o21ai_1
X_6133_ VGND VPWR _2022_ _2019_ net1655 sg13g2_or2_1
X_6064_ _1957_ net1747 _1958_ VPWR VGND _1916_ sg13g2_nand3b_1
X_5015_ VGND VPWR net1469 _1011_ _1013_ _1012_ sg13g2_a21oi_1
XFILLER_39_786 VPWR VGND sg13g2_fill_1
XFILLER_14_609 VPWR VGND sg13g2_fill_1
X_6966_ net1251 _2761_ _2767_ VPWR VGND sg13g2_nor2_1
X_5917_ _0270_ _1826_ _1827_ _3481_ net1627 VPWR VGND sg13g2_a22oi_1
X_6897_ _2707_ net1268 net666 VPWR VGND sg13g2_nand2_1
X_5848_ s0.data_out\[14\]\[0\] s0.data_out\[13\]\[0\] net1397 _1761_ VPWR VGND sg13g2_mux2_1
XFILLER_21_174 VPWR VGND sg13g2_fill_2
X_5779_ VGND VPWR _1689_ _1697_ _1704_ _1681_ sg13g2_a21oi_1
X_7518_ s0.data_out\[0\]\[4\] s0.data_out\[1\]\[4\] net1226 _3268_ VPWR VGND sg13g2_mux2_1
X_7449_ net1219 s0.data_out\[1\]\[7\] _3203_ VPWR VGND sg13g2_and2_1
XFILLER_49_506 VPWR VGND sg13g2_fill_2
XFILLER_27_1013 VPWR VGND sg13g2_decap_8
XFILLER_49_528 VPWR VGND sg13g2_decap_8
XFILLER_1_579 VPWR VGND sg13g2_fill_1
XFILLER_45_712 VPWR VGND sg13g2_decap_4
XFILLER_17_436 VPWR VGND sg13g2_decap_8
XFILLER_45_778 VPWR VGND sg13g2_decap_4
XFILLER_41_940 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
X_7703__322 VPWR VGND net322 sg13g2_tiehi
XFILLER_13_697 VPWR VGND sg13g2_fill_1
XFILLER_0_590 VPWR VGND sg13g2_decap_4
XFILLER_48_550 VPWR VGND sg13g2_decap_8
X_6820_ VGND VPWR net1177 _2606_ _2636_ net1601 sg13g2_a21oi_1
X_6751_ _2573_ _2572_ net1688 _2549_ net1696 VPWR VGND sg13g2_a22oi_1
X_5702_ net1749 net395 _0255_ VPWR VGND sg13g2_and2_1
X_6682_ net1598 _2448_ _2514_ VPWR VGND sg13g2_nor2_1
XFILLER_31_461 VPWR VGND sg13g2_fill_1
X_5633_ net1415 net1345 _1570_ VPWR VGND sg13g2_nor2b_1
X_7823__192 VPWR VGND net192 sg13g2_tiehi
X_5564_ net1429 net527 _1505_ VPWR VGND sg13g2_and2_1
X_4515_ VGND VPWR net1519 _0559_ _0560_ _0557_ sg13g2_a21oi_1
Xhold101 _0117_ VPWR VGND net470 sg13g2_dlygate4sd3_1
X_7303_ _3074_ VPWR _3075_ VGND net1715 net770 sg13g2_o21ai_1
Xhold123 _0130_ VPWR VGND net492 sg13g2_dlygate4sd3_1
X_5495_ _1442_ net1429 _1443_ _1444_ VPWR VGND sg13g2_a21o_1
Xhold112 s0.data_out\[24\]\[1\] VPWR VGND net481 sg13g2_dlygate4sd3_1
Xhold134 s0.data_out\[3\]\[5\] VPWR VGND net503 sg13g2_dlygate4sd3_1
X_4446_ VGND VPWR _3371_ _0488_ _0133_ _0493_ sg13g2_a21oi_1
Xhold156 s0.data_out\[24\]\[7\] VPWR VGND net525 sg13g2_dlygate4sd3_1
Xhold167 s0.data_out\[4\]\[6\] VPWR VGND net536 sg13g2_dlygate4sd3_1
Xhold145 _0294_ VPWR VGND net514 sg13g2_dlygate4sd3_1
X_7234_ VGND VPWR net1234 _3006_ _3008_ _3007_ sg13g2_a21oi_1
X_4377_ VGND VPWR _0434_ _0430_ net1652 sg13g2_or2_1
Xhold189 s0.data_out\[22\]\[7\] VPWR VGND net558 sg13g2_dlygate4sd3_1
X_7165_ VGND VPWR _2947_ _2949_ _2951_ _2950_ sg13g2_a21oi_1
Xhold178 s0.data_out\[8\]\[3\] VPWR VGND net547 sg13g2_dlygate4sd3_1
X_6116_ _2004_ VPWR _2005_ VGND _1995_ _1996_ sg13g2_o21ai_1
X_7096_ _2882_ net1171 _2881_ VPWR VGND sg13g2_nand2_1
X_6047_ _1944_ VPWR _1945_ VGND net1193 _1943_ sg13g2_o21ai_1
XFILLER_39_594 VPWR VGND sg13g2_fill_2
XFILLER_2_1015 VPWR VGND sg13g2_decap_8
XFILLER_42_715 VPWR VGND sg13g2_fill_1
X_6949_ _2752_ VPWR _2753_ VGND net1174 _2751_ sg13g2_o21ai_1
XFILLER_23_984 VPWR VGND sg13g2_decap_8
XFILLER_5_137 VPWR VGND sg13g2_decap_8
XFILLER_2_833 VPWR VGND sg13g2_decap_8
XFILLER_17_233 VPWR VGND sg13g2_decap_8
XFILLER_32_269 VPWR VGND sg13g2_fill_2
XFILLER_14_995 VPWR VGND sg13g2_decap_8
X_4300_ net1559 VPWR _0364_ VGND _3631_ _0363_ sg13g2_o21ai_1
X_5280_ VGND VPWR net1199 _1196_ _1252_ net1619 sg13g2_a21oi_1
X_4231_ _3595_ _3594_ net1687 _3568_ net1695 VPWR VGND sg13g2_a22oi_1
X_4162_ VPWR _3538_ net568 VGND sg13g2_inv_1
X_4093_ VPWR _3469_ net466 VGND sg13g2_inv_1
XFILLER_49_892 VPWR VGND sg13g2_decap_8
X_7921_ net86 VGND VPWR net506 s0.data_out\[4\]\[3\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_7852_ net161 VGND VPWR _0330_ s0.data_out\[10\]\[6\] clknet_leaf_20_clk sg13g2_dfrbpq_2
XFILLER_24_737 VPWR VGND sg13g2_fill_2
X_4995_ net1469 net1335 _0993_ VPWR VGND sg13g2_nor2b_1
X_6803_ net1284 VPWR _2623_ VGND _2553_ _2622_ sg13g2_o21ai_1
X_7783_ net235 VGND VPWR _0261_ s0.data_out\[15\]\[4\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_6734_ VGND VPWR _2443_ _2555_ _2556_ net1282 sg13g2_a21oi_1
X_7943__62 VPWR VGND net62 sg13g2_tiehi
X_6665_ net1672 _2496_ _2499_ VPWR VGND sg13g2_nor2_1
X_6596_ _2430_ _2432_ _2433_ VPWR VGND sg13g2_nor2_1
XFILLER_20_998 VPWR VGND sg13g2_decap_8
X_5616_ _1551_ net1415 _1552_ _1553_ VPWR VGND sg13g2_a21o_1
X_5547_ net1622 _1428_ _1492_ VPWR VGND sg13g2_nor2_1
X_5478_ _1427_ net466 net1446 VPWR VGND sg13g2_nand2b_1
X_4429_ net1549 VPWR _0479_ VGND _0419_ _0478_ sg13g2_o21ai_1
X_7217_ net1720 net371 _0062_ VPWR VGND sg13g2_and2_1
XFILLER_48_14 VPWR VGND sg13g2_decap_4
Xfanout1409 s0.valid_out\[14\][0] net1409 VPWR VGND sg13g2_buf_2
X_7148_ _2934_ net604 net1253 VPWR VGND sg13g2_nand2b_1
XFILLER_47_829 VPWR VGND sg13g2_decap_8
X_7079_ net1248 VPWR _2868_ VGND net1639 net1241 sg13g2_o21ai_1
XFILLER_39_380 VPWR VGND sg13g2_fill_1
XFILLER_14_236 VPWR VGND sg13g2_decap_4
XFILLER_22_280 VPWR VGND sg13g2_fill_2
XFILLER_7_936 VPWR VGND sg13g2_fill_1
XFILLER_11_998 VPWR VGND sg13g2_decap_8
XFILLER_7_969 VPWR VGND sg13g2_decap_8
X_7700__325 VPWR VGND net325 sg13g2_tiehi
XFILLER_37_317 VPWR VGND sg13g2_fill_1
XFILLER_46_862 VPWR VGND sg13g2_decap_8
XFILLER_33_523 VPWR VGND sg13g2_fill_2
X_7963__191 VPWR VGND net191 sg13g2_tiehi
X_4780_ VPWR _0161_ net741 VGND sg13g2_inv_1
X_6450_ net1311 s0.data_out\[9\]\[6\] _2301_ VPWR VGND sg13g2_and2_1
X_7940__65 VPWR VGND net65 sg13g2_tiehi
Xclkload10 VPWR clkload10/Y clknet_leaf_23_clk VGND sg13g2_inv_1
X_7820__195 VPWR VGND net195 sg13g2_tiehi
X_6381_ net1311 net1330 _2239_ VPWR VGND sg13g2_nor2b_1
X_5401_ VGND VPWR net1436 net689 _1361_ _1301_ sg13g2_a21oi_1
XFILLER_6_980 VPWR VGND sg13g2_decap_8
X_5332_ s0.data_out\[18\]\[1\] s0.data_out\[17\]\[1\] net1443 _1293_ VPWR VGND sg13g2_mux2_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_5263_ _1236_ net1455 net499 VPWR VGND sg13g2_nand2_1
X_5194_ VGND VPWR net1635 net1453 _1170_ _1169_ sg13g2_a21oi_1
X_4214_ _3386_ VPWR _3578_ VGND s0.valid_out\[27\][0] s0.data_out\[26\]\[0\] sg13g2_o21ai_1
X_7002_ _2800_ _2799_ net1688 _2776_ net1700 VPWR VGND sg13g2_a22oi_1
X_4145_ VPWR _3521_ net796 VGND sg13g2_inv_1
XFILLER_28_317 VPWR VGND sg13g2_fill_1
XFILLER_28_328 VPWR VGND sg13g2_fill_1
X_4076_ VPWR _3452_ net645 VGND sg13g2_inv_1
X_7904_ net104 VGND VPWR _0038_ s0.genblk1\[4\].modules.bubble clknet_leaf_3_clk sg13g2_dfrbpq_1
X_7835_ net179 VGND VPWR net442 s0.was_valid_out\[10\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_24_545 VPWR VGND sg13g2_fill_1
X_4978_ net1471 net1347 _0976_ VPWR VGND sg13g2_nor2b_1
X_7766_ net253 VGND VPWR _0244_ s0.shift_out\[16\][0] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_6717_ net1729 VPWR _2542_ VGND _2539_ _2541_ sg13g2_o21ai_1
X_7697_ net328 VGND VPWR _0175_ s0.data_out\[22\]\[2\] clknet_leaf_37_clk sg13g2_dfrbpq_2
Xclkload4 clkload4/Y clknet_leaf_6_clk VPWR VGND sg13g2_inv_2
X_6648_ VGND VPWR _2482_ _2473_ net1661 sg13g2_or2_1
XFILLER_4_906 VPWR VGND sg13g2_decap_8
X_6579_ _3394_ _3508_ _2418_ VPWR VGND sg13g2_nor2_1
XFILLER_8_1010 VPWR VGND sg13g2_decap_8
Xfanout1206 net1207 net1206 VPWR VGND sg13g2_buf_8
Xfanout1228 net1229 net1228 VPWR VGND sg13g2_buf_2
Xfanout1217 net1218 net1217 VPWR VGND sg13g2_buf_2
Xfanout1239 net440 net1239 VPWR VGND sg13g2_buf_8
XFILLER_47_615 VPWR VGND sg13g2_fill_1
XFILLER_46_114 VPWR VGND sg13g2_fill_1
X_7767__252 VPWR VGND net252 sg13g2_tiehi
XFILLER_43_898 VPWR VGND sg13g2_fill_1
XFILLER_30_548 VPWR VGND sg13g2_fill_2
XFILLER_6_243 VPWR VGND sg13g2_fill_2
XFILLER_11_795 VPWR VGND sg13g2_fill_2
X_7774__245 VPWR VGND net245 sg13g2_tiehi
Xfanout1740 net1741 net1740 VPWR VGND sg13g2_buf_8
Xfanout1751 rst_n net1751 VPWR VGND sg13g2_buf_8
Xheichips25_top_sorter_13 VPWR VGND uio_oe[3] sg13g2_tielo
X_5950_ net1383 _1848_ _1854_ VPWR VGND sg13g2_nor2_1
XFILLER_46_681 VPWR VGND sg13g2_decap_8
X_4901_ VGND VPWR _0885_ _0908_ _0910_ _0909_ sg13g2_a21oi_1
XFILLER_18_394 VPWR VGND sg13g2_fill_1
XFILLER_34_832 VPWR VGND sg13g2_fill_1
X_7620_ VGND VPWR net1721 _3335_ _0102_ _3354_ sg13g2_a21oi_1
XFILLER_45_191 VPWR VGND sg13g2_fill_1
X_5881_ VGND VPWR _1794_ _1791_ net1666 sg13g2_or2_1
X_4832_ _0838_ _0840_ _0841_ VPWR VGND sg13g2_and2_1
X_7551_ VGND VPWR net1200 _3236_ _3297_ net1587 sg13g2_a21oi_1
X_4763_ _0784_ net1181 _0783_ VPWR VGND sg13g2_nand2_1
X_7482_ _3232_ net1218 _3231_ VPWR VGND sg13g2_nand2b_1
X_4694_ VGND VPWR _3370_ _0712_ _0157_ _0717_ sg13g2_a21oi_1
X_6502_ VGND VPWR _2228_ _2347_ _2348_ net1305 sg13g2_a21oi_1
X_6433_ net1307 net485 _2288_ VPWR VGND sg13g2_and2_1
X_6364_ VGND VPWR net1307 _2220_ _2222_ _2221_ sg13g2_a21oi_1
X_5315_ VGND VPWR net1636 net1456 _1279_ net1452 sg13g2_a21oi_1
X_6295_ net1365 VPWR _2169_ VGND _2089_ _2168_ sg13g2_o21ai_1
X_5246_ _1217_ net1449 _1218_ _1219_ VPWR VGND sg13g2_a21o_1
Xhold38 s0.data_out\[24\]\[5\] VPWR VGND net407 sg13g2_dlygate4sd3_1
Xhold16 s0.genblk1\[22\].modules.bubble VPWR VGND net385 sg13g2_dlygate4sd3_1
Xhold27 s0.genblk1\[15\].modules.bubble VPWR VGND net396 sg13g2_dlygate4sd3_1
Xhold49 s0.data_out\[12\]\[4\] VPWR VGND net418 sg13g2_dlygate4sd3_1
X_5177_ net1473 VPWR _1157_ VGND _1120_ _1156_ sg13g2_o21ai_1
XFILLER_21_1019 VPWR VGND sg13g2_decap_8
X_4128_ VPWR _3504_ net544 VGND sg13g2_inv_1
XFILLER_43_106 VPWR VGND sg13g2_fill_1
X_4059_ VPWR _3435_ s0.data_out\[23\]\[2\] VGND sg13g2_inv_1
X_7818_ net197 VGND VPWR net598 s0.data_out\[12\]\[3\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_7749_ net272 VGND VPWR _0227_ s0.data_out\[18\]\[6\] clknet_leaf_32_clk sg13g2_dfrbpq_2
XFILLER_0_964 VPWR VGND sg13g2_decap_8
XFILLER_48_935 VPWR VGND sg13g2_decap_8
XFILLER_43_651 VPWR VGND sg13g2_fill_2
XFILLER_31_879 VPWR VGND sg13g2_fill_2
XFILLER_30_356 VPWR VGND sg13g2_fill_2
X_6080_ _1969_ VPWR _1972_ VGND net1379 _1971_ sg13g2_o21ai_1
XFILLER_3_791 VPWR VGND sg13g2_decap_8
X_5100_ VGND VPWR net1458 _1083_ _1085_ _1084_ sg13g2_a21oi_1
X_5031_ VGND VPWR _1023_ _1027_ _0183_ _1028_ sg13g2_a21oi_1
XFILLER_39_957 VPWR VGND sg13g2_decap_8
Xfanout1581 net1588 net1581 VPWR VGND sg13g2_buf_1
Xfanout1592 net1603 net1592 VPWR VGND sg13g2_buf_2
Xfanout1570 _3418_ net1570 VPWR VGND sg13g2_buf_8
XFILLER_47_990 VPWR VGND sg13g2_decap_8
XFILLER_19_670 VPWR VGND sg13g2_decap_4
X_6982_ net1250 net1353 _2780_ VPWR VGND sg13g2_nor2b_1
X_5933_ net1629 _1809_ _1840_ VPWR VGND sg13g2_nor2_1
X_5864_ _1776_ VPWR _1777_ VGND _1767_ _1768_ sg13g2_o21ai_1
XFILLER_33_161 VPWR VGND sg13g2_fill_1
X_7603_ _3341_ _3340_ net1689 _3335_ net1696 VPWR VGND sg13g2_a22oi_1
X_4815_ VGND VPWR net1635 net1505 _0827_ net1498 sg13g2_a21oi_1
XFILLER_22_846 VPWR VGND sg13g2_fill_1
XFILLER_33_183 VPWR VGND sg13g2_fill_1
X_7534_ VGND VPWR _3284_ net1565 net397 sg13g2_or2_1
X_5795_ _1716_ VPWR _1717_ VGND net1197 _1715_ sg13g2_o21ai_1
X_4746_ _0767_ _0766_ net1660 _0759_ net1650 VPWR VGND sg13g2_a22oi_1
X_7465_ s0.data_out\[0\]\[2\] s0.data_out\[1\]\[2\] net1226 _3215_ VPWR VGND sg13g2_mux2_1
X_4677_ _0154_ net611 _0703_ _3427_ net1592 VPWR VGND sg13g2_a22oi_1
X_6416_ _2254_ _2270_ _2273_ _2274_ VPWR VGND sg13g2_nor3_1
X_7396_ _3042_ VPWR _3158_ VGND net1237 _3541_ sg13g2_o21ai_1
X_6347_ _2205_ net1314 net485 VPWR VGND sg13g2_nand2_1
XFILLER_0_227 VPWR VGND sg13g2_fill_2
X_6278_ net1690 _2116_ _2155_ VPWR VGND sg13g2_nor2_1
X_5229_ net1447 net1168 _1202_ VPWR VGND sg13g2_nor2_1
XFILLER_45_949 VPWR VGND sg13g2_decap_8
XFILLER_13_835 VPWR VGND sg13g2_fill_1
X_7764__255 VPWR VGND net255 sg13g2_tiehi
XFILLER_8_327 VPWR VGND sg13g2_decap_4
X_7771__248 VPWR VGND net248 sg13g2_tiehi
XFILLER_0_761 VPWR VGND sg13g2_decap_8
XFILLER_48_732 VPWR VGND sg13g2_decap_8
XFILLER_11_8 VPWR VGND sg13g2_fill_1
XFILLER_44_960 VPWR VGND sg13g2_decap_8
X_4600_ net1703 _0626_ _0633_ VPWR VGND sg13g2_nor2_1
X_5580_ net1748 net396 _0243_ VPWR VGND sg13g2_and2_1
X_4531_ net1521 net626 _0575_ VPWR VGND sg13g2_and2_1
XFILLER_7_85 VPWR VGND sg13g2_fill_1
X_4462_ _0507_ net1538 _0506_ VPWR VGND sg13g2_nand2b_1
Xhold316 s0.data_out\[4\]\[2\] VPWR VGND net685 sg13g2_dlygate4sd3_1
Xhold305 s0.data_out\[8\]\[2\] VPWR VGND net674 sg13g2_dlygate4sd3_1
X_7250_ _3024_ net1236 s0.data_out\[2\]\[6\] VPWR VGND sg13g2_nand2_1
X_6201_ net463 _2080_ _2081_ VPWR VGND sg13g2_nor2_1
Xhold327 s0.data_out\[14\]\[6\] VPWR VGND net696 sg13g2_dlygate4sd3_1
Xhold349 s0.data_out\[21\]\[6\] VPWR VGND net718 sg13g2_dlygate4sd3_1
Xhold338 s0.data_out\[25\]\[1\] VPWR VGND net707 sg13g2_dlygate4sd3_1
X_4393_ _0450_ _0449_ net1668 _0442_ net1677 VPWR VGND sg13g2_a22oi_1
X_7181_ _2963_ VPWR _2964_ VGND net1171 _2962_ sg13g2_o21ai_1
X_6132_ net1665 _2012_ _2021_ VPWR VGND sg13g2_nor2_1
XFILLER_30_0 VPWR VGND sg13g2_fill_1
X_6063_ net1393 VPWR _1957_ VGND _1913_ _1956_ sg13g2_o21ai_1
X_5014_ net1469 net1346 _1012_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_242 VPWR VGND sg13g2_fill_2
XFILLER_26_404 VPWR VGND sg13g2_fill_2
XFILLER_42_919 VPWR VGND sg13g2_decap_8
XFILLER_42_908 VPWR VGND sg13g2_fill_2
X_6965_ _2763_ VPWR _2766_ VGND net400 net1255 sg13g2_o21ai_1
XFILLER_26_448 VPWR VGND sg13g2_fill_2
X_5916_ net1626 _1759_ _1827_ VPWR VGND sg13g2_nor2_1
X_6896_ _2703_ _2704_ _2706_ VPWR VGND _2705_ sg13g2_nand3b_1
XFILLER_10_827 VPWR VGND sg13g2_fill_2
X_5847_ VGND VPWR net1402 _1757_ _1760_ _1759_ sg13g2_a21oi_1
XFILLER_10_849 VPWR VGND sg13g2_fill_2
XFILLER_21_164 VPWR VGND sg13g2_fill_1
X_5778_ _1702_ VPWR _1703_ VGND _1660_ _1662_ sg13g2_o21ai_1
X_7517_ VPWR _3267_ _3266_ VGND sg13g2_inv_1
X_4729_ _0731_ _0740_ _0741_ _0749_ _0750_ VPWR VGND sg13g2_nor4_1
X_7448_ VPWR _0082_ _3202_ VGND sg13g2_inv_1
X_7379_ _3139_ net1217 _3140_ _3141_ VPWR VGND sg13g2_a21o_1
XFILLER_29_231 VPWR VGND sg13g2_fill_1
XFILLER_44_212 VPWR VGND sg13g2_fill_2
XFILLER_45_757 VPWR VGND sg13g2_decap_8
XFILLER_41_996 VPWR VGND sg13g2_decap_8
XFILLER_5_897 VPWR VGND sg13g2_fill_1
XFILLER_5_886 VPWR VGND sg13g2_fill_2
XFILLER_36_757 VPWR VGND sg13g2_fill_2
XFILLER_24_919 VPWR VGND sg13g2_fill_1
X_6750_ VGND VPWR net1284 _2569_ _2572_ _2571_ sg13g2_a21oi_1
XFILLER_35_267 VPWR VGND sg13g2_fill_2
X_5701_ net1748 _1622_ _0254_ VPWR VGND sg13g2_and2_1
X_6681_ net1293 VPWR _2513_ VGND _2445_ _2512_ sg13g2_o21ai_1
X_5632_ s0.data_out\[16\]\[4\] s0.data_out\[15\]\[4\] net1421 _1569_ VPWR VGND sg13g2_mux2_1
XFILLER_32_996 VPWR VGND sg13g2_decap_8
X_5563_ VPWR _0239_ net754 VGND sg13g2_inv_1
X_4514_ s0.data_out\[25\]\[4\] s0.data_out\[24\]\[4\] net1528 _0559_ VPWR VGND sg13g2_mux2_1
X_7302_ _2997_ _3073_ net1715 _3074_ VPWR VGND sg13g2_nand3_1
Xhold102 s0.was_valid_out\[7\][0] VPWR VGND net471 sg13g2_dlygate4sd3_1
Xhold124 s0.data_out\[10\]\[5\] VPWR VGND net493 sg13g2_dlygate4sd3_1
X_5494_ net1429 net1335 _1443_ VPWR VGND sg13g2_nor2b_1
Xhold113 _0150_ VPWR VGND net482 sg13g2_dlygate4sd3_1
Xhold135 _0069_ VPWR VGND net504 sg13g2_dlygate4sd3_1
X_4445_ net1725 VPWR _0493_ VGND _0490_ _0492_ sg13g2_o21ai_1
Xhold146 s0.data_out\[27\]\[7\] VPWR VGND net515 sg13g2_dlygate4sd3_1
Xhold157 _0156_ VPWR VGND net526 sg13g2_dlygate4sd3_1
Xhold168 _0058_ VPWR VGND net537 sg13g2_dlygate4sd3_1
X_7233_ net1234 net1348 _3007_ VPWR VGND sg13g2_nor2b_1
X_4376_ net1647 _0430_ _0433_ VPWR VGND sg13g2_nor2_1
X_7164_ _2872_ VPWR _2950_ VGND _2943_ _2945_ sg13g2_o21ai_1
Xhold179 _0007_ VPWR VGND net548 sg13g2_dlygate4sd3_1
X_6115_ _2004_ _2003_ net1693 _1980_ net1698 VPWR VGND sg13g2_a22oi_1
X_7095_ s0.data_out\[3\]\[2\] s0.data_out\[4\]\[2\] net1253 _2881_ VPWR VGND sg13g2_mux2_1
X_6046_ VGND VPWR net1192 _1862_ _1944_ net1627 sg13g2_a21oi_1
XFILLER_26_234 VPWR VGND sg13g2_fill_2
XFILLER_27_757 VPWR VGND sg13g2_fill_1
X_6948_ VGND VPWR net1174 _2712_ _2752_ net1597 sg13g2_a21oi_1
X_6879_ _2689_ net1267 net584 VPWR VGND sg13g2_nand2_1
XFILLER_22_473 VPWR VGND sg13g2_decap_4
XFILLER_2_812 VPWR VGND sg13g2_decap_8
XFILLER_2_889 VPWR VGND sg13g2_decap_8
XFILLER_40_1011 VPWR VGND sg13g2_decap_8
XFILLER_32_204 VPWR VGND sg13g2_decap_4
XFILLER_17_289 VPWR VGND sg13g2_fill_2
XFILLER_9_455 VPWR VGND sg13g2_decap_8
X_4230_ VGND VPWR net1560 _3593_ _3594_ _3589_ sg13g2_a21oi_1
X_4161_ VPWR _3537_ net616 VGND sg13g2_inv_1
X_4092_ VPWR _3468_ net791 VGND sg13g2_inv_1
XFILLER_49_871 VPWR VGND sg13g2_decap_8
XFILLER_36_521 VPWR VGND sg13g2_fill_2
X_7920_ net87 VGND VPWR _0054_ s0.data_out\[4\]\[2\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_7851_ net162 VGND VPWR net494 s0.data_out\[10\]\[5\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_6802_ net1175 _3523_ _2622_ VPWR VGND sg13g2_nor2_1
X_4994_ s0.data_out\[21\]\[6\] s0.data_out\[20\]\[6\] net1478 _0992_ VPWR VGND sg13g2_mux2_1
X_7782_ net236 VGND VPWR net766 s0.data_out\[15\]\[3\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_6733_ _2555_ net694 net1289 VPWR VGND sg13g2_nand2b_1
X_6664_ net1680 _2490_ _2498_ VPWR VGND sg13g2_nor2_1
XFILLER_20_977 VPWR VGND sg13g2_decap_8
X_5615_ net1416 net1330 _1552_ VPWR VGND sg13g2_nor2b_1
X_6595_ _2431_ VPWR _2432_ VGND net1287 _2425_ sg13g2_o21ai_1
X_5546_ net1438 VPWR _1491_ VGND _1425_ _1490_ sg13g2_o21ai_1
X_5477_ _1424_ net1431 _1425_ _1426_ VPWR VGND sg13g2_a21o_1
X_4428_ net1533 s0.data_out\[25\]\[6\] _0478_ VPWR VGND sg13g2_and2_1
X_7216_ net1714 _2986_ _0061_ VPWR VGND sg13g2_and2_1
X_4359_ _0415_ VPWR _0416_ VGND _0406_ _0407_ sg13g2_o21ai_1
X_7147_ _2931_ net1241 _2932_ _2933_ VPWR VGND sg13g2_a21o_1
XFILLER_47_808 VPWR VGND sg13g2_decap_8
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
X_7078_ _0047_ _2866_ _2867_ _3524_ net1596 VPWR VGND sg13g2_a22oi_1
X_6029_ _1926_ _1928_ _1925_ _1930_ VPWR VGND sg13g2_nand3_1
XFILLER_27_576 VPWR VGND sg13g2_fill_2
XFILLER_42_524 VPWR VGND sg13g2_decap_8
XFILLER_7_915 VPWR VGND sg13g2_fill_2
XFILLER_11_977 VPWR VGND sg13g2_decap_8
XFILLER_7_948 VPWR VGND sg13g2_decap_8
XFILLER_13_62 VPWR VGND sg13g2_fill_2
XFILLER_8_0 VPWR VGND sg13g2_fill_2
XFILLER_38_70 VPWR VGND sg13g2_fill_1
XFILLER_46_841 VPWR VGND sg13g2_decap_8
X_6380_ s0.data_out\[10\]\[7\] s0.data_out\[9\]\[7\] net1317 _2238_ VPWR VGND sg13g2_mux2_1
X_5400_ VGND VPWR _1356_ _1359_ _0220_ _1360_ sg13g2_a21oi_1
Xclkload11 clkload11/Y clknet_leaf_25_clk VPWR VGND sg13g2_inv_2
X_5331_ _1292_ net1443 net813 VPWR VGND sg13g2_nand2_1
X_5262_ net1449 net1345 _1235_ VPWR VGND sg13g2_nor2b_1
X_7001_ VGND VPWR net1259 _2796_ _2799_ _2798_ sg13g2_a21oi_1
X_4213_ _3577_ net1701 _3576_ VPWR VGND sg13g2_nand2_1
X_5193_ net1461 VPWR _1169_ VGND net1644 net1448 sg13g2_o21ai_1
X_4144_ VPWR _3520_ net719 VGND sg13g2_inv_1
XFILLER_18_18 VPWR VGND sg13g2_decap_4
X_4075_ VPWR _3451_ net672 VGND sg13g2_inv_1
X_7903_ net105 VGND VPWR _0037_ s0.valid_out\[5\][0] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_7834_ net180 VGND VPWR net587 s0.data_out\[11\]\[7\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_7765_ net254 VGND VPWR _0243_ s0.genblk1\[15\].modules.bubble clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_6716_ _2540_ VPWR _2541_ VGND _2535_ _2538_ sg13g2_o21ai_1
X_4977_ s0.data_out\[21\]\[3\] s0.data_out\[20\]\[3\] net1478 _0975_ VPWR VGND sg13g2_mux2_1
Xclkload5 VPWR clkload5/Y clknet_leaf_13_clk VGND sg13g2_inv_1
X_7696_ net329 VGND VPWR net600 s0.data_out\[22\]\[1\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_6647_ _2481_ _2480_ net1651 _2473_ net1661 VPWR VGND sg13g2_a22oi_1
X_6578_ VPWR _0341_ _2417_ VGND sg13g2_inv_1
XFILLER_30_1021 VPWR VGND sg13g2_decap_8
X_5529_ VGND VPWR _1478_ net1567 net393 sg13g2_or2_1
Xfanout1207 _3375_ net1207 VPWR VGND sg13g2_buf_8
Xfanout1229 net1231 net1229 VPWR VGND sg13g2_buf_1
Xfanout1218 net1219 net1218 VPWR VGND sg13g2_buf_8
XFILLER_28_885 VPWR VGND sg13g2_fill_2
XFILLER_27_395 VPWR VGND sg13g2_fill_1
XFILLER_40_60 VPWR VGND sg13g2_fill_1
XFILLER_3_984 VPWR VGND sg13g2_decap_8
Xfanout1730 net1732 net1730 VPWR VGND sg13g2_buf_8
Xfanout1741 net1751 net1741 VPWR VGND sg13g2_buf_8
XFILLER_19_841 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_14 VPWR VGND uio_oe[4] sg13g2_tielo
XFILLER_19_863 VPWR VGND sg13g2_fill_1
X_5880_ VGND VPWR _1793_ _1784_ net1656 sg13g2_or2_1
X_4900_ _0828_ VPWR _0909_ VGND _0881_ _0884_ sg13g2_o21ai_1
X_4831_ _0840_ _0839_ net1500 VPWR VGND sg13g2_nand2b_1
XFILLER_34_899 VPWR VGND sg13g2_fill_1
X_7550_ VGND VPWR net1211 net433 _3296_ _3238_ sg13g2_a21oi_1
X_4762_ s0.data_out\[22\]\[4\] s0.data_out\[23\]\[4\] net1516 _0783_ VPWR VGND sg13g2_mux2_1
XFILLER_21_549 VPWR VGND sg13g2_fill_1
X_7481_ VGND VPWR net1208 _3229_ _3231_ _3230_ sg13g2_a21oi_1
X_4693_ net1727 VPWR _0717_ VGND _0714_ _0716_ sg13g2_o21ai_1
XFILLER_14_1016 VPWR VGND sg13g2_decap_8
XFILLER_14_1027 VPWR VGND sg13g2_fill_2
X_6501_ _2347_ net547 net1314 VPWR VGND sg13g2_nand2b_1
X_6432_ _0325_ _2286_ _2287_ _3498_ net1609 VPWR VGND sg13g2_a22oi_1
X_6363_ net1308 net1359 _2221_ VPWR VGND sg13g2_nor2b_1
X_5314_ VGND VPWR _1277_ _1278_ net1444 net1635 sg13g2_a21oi_2
X_6294_ net1321 net523 _2168_ VPWR VGND sg13g2_and2_1
X_5245_ net1449 net1331 _1218_ VPWR VGND sg13g2_nor2b_1
Xhold17 s0.genblk1\[6\].modules.bubble VPWR VGND net386 sg13g2_dlygate4sd3_1
Xhold28 s0.genblk1\[1\].modules.bubble VPWR VGND net397 sg13g2_dlygate4sd3_1
XFILLER_29_39 VPWR VGND sg13g2_fill_1
Xhold39 _0672_ VPWR VGND net408 sg13g2_dlygate4sd3_1
X_5176_ net1198 _3453_ _1156_ VPWR VGND sg13g2_nor2_1
XFILLER_28_104 VPWR VGND sg13g2_fill_1
X_4127_ VPWR _3503_ net483 VGND sg13g2_inv_1
X_4058_ VPWR _3434_ net810 VGND sg13g2_inv_1
XFILLER_24_321 VPWR VGND sg13g2_decap_8
XFILLER_24_343 VPWR VGND sg13g2_fill_2
X_7817_ net198 VGND VPWR net790 s0.data_out\[12\]\[2\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_7748_ net273 VGND VPWR net701 s0.data_out\[18\]\[5\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_7679_ net348 VGND VPWR net410 s0.was_valid_out\[23\][0] clknet_leaf_42_clk sg13g2_dfrbpq_1
XFILLER_0_943 VPWR VGND sg13g2_decap_8
XFILLER_48_914 VPWR VGND sg13g2_decap_8
XFILLER_43_663 VPWR VGND sg13g2_fill_2
XFILLER_16_855 VPWR VGND sg13g2_fill_2
XFILLER_7_520 VPWR VGND sg13g2_fill_1
XFILLER_44_1009 VPWR VGND sg13g2_decap_8
XFILLER_3_770 VPWR VGND sg13g2_decap_8
X_5030_ VGND VPWR _1028_ net1567 net389 sg13g2_or2_1
XFILLER_39_936 VPWR VGND sg13g2_decap_8
Xfanout1560 net1562 net1560 VPWR VGND sg13g2_buf_8
Xfanout1593 net1595 net1593 VPWR VGND sg13g2_buf_8
Xfanout1582 net1584 net1582 VPWR VGND sg13g2_buf_8
Xfanout1571 net1574 net1571 VPWR VGND sg13g2_buf_8
X_6981_ _2778_ VPWR _2779_ VGND net1255 _3530_ sg13g2_o21ai_1
X_5932_ net1406 VPWR _1839_ VGND _1806_ _1838_ sg13g2_o21ai_1
X_5863_ _1776_ _1775_ net1693 _1752_ net1698 VPWR VGND sg13g2_a22oi_1
X_7602_ _3340_ _3339_ VPWR VGND sg13g2_inv_2
X_4814_ _0824_ _0825_ _0826_ VPWR VGND sg13g2_nor2_1
X_5794_ VGND VPWR net1197 _1646_ _1716_ net1626 sg13g2_a21oi_1
X_7533_ _3209_ _3281_ _3282_ _3283_ VPWR VGND sg13g2_nor3_1
X_4745_ VGND VPWR net1512 _0763_ _0766_ _0765_ sg13g2_a21oi_1
X_4676_ net1589 net408 _0703_ VPWR VGND sg13g2_nor2_1
X_7464_ net1742 net372 _0086_ VPWR VGND sg13g2_and2_1
X_7395_ VGND VPWR net1221 _3155_ _3157_ _3156_ sg13g2_a21oi_1
X_6415_ _2271_ VPWR _2273_ VGND net1691 _2234_ sg13g2_o21ai_1
X_6346_ net1328 net1649 net1 _0322_ VPWR VGND sg13g2_mux2_1
X_7757__263 VPWR VGND net263 sg13g2_tiehi
XFILLER_0_239 VPWR VGND sg13g2_fill_2
X_6277_ _2153_ VPWR _2154_ VGND net1682 _2143_ sg13g2_o21ai_1
XFILLER_5_1014 VPWR VGND sg13g2_decap_8
X_5228_ _1200_ VPWR _1201_ VGND net1454 _3454_ sg13g2_o21ai_1
X_5159_ net1458 s0.data_out\[19\]\[0\] _1143_ VPWR VGND sg13g2_and2_1
XFILLER_45_928 VPWR VGND sg13g2_decap_8
XFILLER_16_118 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_36_clk clknet_3_4__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_12_346 VPWR VGND sg13g2_fill_2
XFILLER_0_740 VPWR VGND sg13g2_decap_8
XFILLER_48_711 VPWR VGND sg13g2_decap_8
XFILLER_48_788 VPWR VGND sg13g2_decap_8
XFILLER_16_641 VPWR VGND sg13g2_fill_2
XFILLER_16_652 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_27_clk clknet_3_4__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_35_449 VPWR VGND sg13g2_fill_2
XFILLER_16_685 VPWR VGND sg13g2_fill_2
XFILLER_31_611 VPWR VGND sg13g2_decap_4
XFILLER_12_880 VPWR VGND sg13g2_fill_2
X_4530_ VGND VPWR _0570_ _0573_ _0136_ _0574_ sg13g2_a21oi_1
XFILLER_11_1019 VPWR VGND sg13g2_decap_8
XFILLER_30_198 VPWR VGND sg13g2_fill_1
X_4461_ VGND VPWR net1521 _0505_ _0506_ _0503_ sg13g2_a21oi_1
Xhold317 _2965_ VPWR VGND net686 sg13g2_dlygate4sd3_1
Xhold306 s0.data_out\[11\]\[1\] VPWR VGND net675 sg13g2_dlygate4sd3_1
Xhold328 _1844_ VPWR VGND net697 sg13g2_dlygate4sd3_1
X_6200_ _2079_ VPWR _2080_ VGND net1369 _1964_ sg13g2_o21ai_1
Xhold339 _0138_ VPWR VGND net708 sg13g2_dlygate4sd3_1
X_7180_ VGND VPWR net1171 _2881_ _2963_ net1581 sg13g2_a21oi_1
X_6131_ _2020_ _2019_ net1655 _2012_ net1665 VPWR VGND sg13g2_a22oi_1
X_4392_ VGND VPWR net1549 _0446_ _0449_ _0448_ sg13g2_a21oi_1
X_6062_ net1383 s0.data_out\[12\]\[6\] _1956_ VPWR VGND sg13g2_and2_1
XFILLER_23_0 VPWR VGND sg13g2_fill_1
X_5013_ s0.data_out\[21\]\[4\] s0.data_out\[20\]\[4\] net1479 _1011_ VPWR VGND sg13g2_mux2_1
Xfanout1390 net1391 net1390 VPWR VGND sg13g2_buf_8
XFILLER_39_799 VPWR VGND sg13g2_fill_2
XFILLER_26_18 VPWR VGND sg13g2_fill_2
XFILLER_26_416 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_18_clk clknet_3_6__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
X_6964_ _2763_ _2764_ _2765_ VPWR VGND sg13g2_nor2_1
X_6895_ net1650 _2702_ _2705_ VPWR VGND sg13g2_nor2_1
XFILLER_22_611 VPWR VGND sg13g2_decap_4
X_5915_ net1401 VPWR _1826_ VGND _1756_ _1825_ sg13g2_o21ai_1
XFILLER_35_983 VPWR VGND sg13g2_decap_8
X_5846_ VGND VPWR _1628_ _1758_ _1759_ net1401 sg13g2_a21oi_1
X_5777_ _1681_ _1698_ _1699_ _1701_ _1702_ VPWR VGND sg13g2_nor4_1
X_7516_ _3261_ _3265_ net1669 _3266_ VPWR VGND sg13g2_nand3_1
X_4728_ net1690 _0748_ _0749_ VPWR VGND sg13g2_nor2_1
X_4659_ net1526 VPWR _0690_ VGND _0622_ _0689_ sg13g2_o21ai_1
X_7447_ _3201_ VPWR _3202_ VGND net1718 net725 sg13g2_o21ai_1
X_7378_ net1217 net1334 _3140_ VPWR VGND sg13g2_nor2b_1
X_6329_ net1738 VPWR _2197_ VGND _2192_ _2194_ sg13g2_o21ai_1
XFILLER_29_221 VPWR VGND sg13g2_fill_1
XFILLER_45_736 VPWR VGND sg13g2_decap_8
XFILLER_29_298 VPWR VGND sg13g2_fill_1
XFILLER_26_961 VPWR VGND sg13g2_fill_1
XFILLER_13_644 VPWR VGND sg13g2_fill_2
XFILLER_41_975 VPWR VGND sg13g2_decap_8
XFILLER_34_1019 VPWR VGND sg13g2_decap_8
XFILLER_40_485 VPWR VGND sg13g2_fill_1
XFILLER_9_637 VPWR VGND sg13g2_fill_1
XFILLER_32_94 VPWR VGND sg13g2_fill_2
XFILLER_4_331 VPWR VGND sg13g2_fill_2
XFILLER_48_585 VPWR VGND sg13g2_decap_8
XFILLER_17_983 VPWR VGND sg13g2_decap_8
XFILLER_35_257 VPWR VGND sg13g2_fill_2
X_5700_ VGND VPWR _3365_ _1622_ _0253_ _1627_ sg13g2_a21oi_1
X_6680_ net1177 _3514_ _2512_ VPWR VGND sg13g2_nor2_1
XFILLER_32_975 VPWR VGND sg13g2_decap_8
XFILLER_31_485 VPWR VGND sg13g2_fill_1
X_5631_ _1568_ net1420 s0.data_out\[15\]\[4\] VPWR VGND sg13g2_nand2_1
X_5562_ _1503_ VPWR _1504_ VGND net1745 net753 sg13g2_o21ai_1
X_4513_ _0558_ net1530 net698 VPWR VGND sg13g2_nand2_1
X_7301_ net1239 VPWR _3073_ VGND _2994_ _3072_ sg13g2_o21ai_1
Xhold125 _0329_ VPWR VGND net494 sg13g2_dlygate4sd3_1
Xhold114 s0.data_out\[9\]\[7\] VPWR VGND net483 sg13g2_dlygate4sd3_1
Xhold103 s0.data_out\[27\]\[6\] VPWR VGND net472 sg13g2_dlygate4sd3_1
X_5493_ s0.data_out\[17\]\[6\] s0.data_out\[16\]\[6\] net1433 _1442_ VPWR VGND sg13g2_mux2_1
X_7232_ s0.data_out\[3\]\[2\] s0.data_out\[2\]\[2\] net1238 _3006_ VPWR VGND sg13g2_mux2_1
X_4444_ _0492_ _0489_ _0491_ VPWR VGND sg13g2_nand2_1
Xhold147 _0120_ VPWR VGND net516 sg13g2_dlygate4sd3_1
Xhold158 s0.data_out\[16\]\[7\] VPWR VGND net527 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_3_2__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold136 s0.data_out\[4\]\[3\] VPWR VGND net505 sg13g2_dlygate4sd3_1
X_4375_ net1658 _0423_ _0432_ VPWR VGND sg13g2_nor2_1
Xhold169 s0.data_out\[21\]\[7\] VPWR VGND net538 sg13g2_dlygate4sd3_1
X_7163_ _2927_ _2919_ _2916_ _2949_ VPWR VGND sg13g2_a21o_1
X_7754__266 VPWR VGND net266 sg13g2_tiehi
X_7094_ VGND VPWR net1240 _2878_ _2880_ _2879_ sg13g2_a21oi_1
X_6114_ VGND VPWR net1377 _2000_ _2003_ _2002_ sg13g2_a21oi_1
X_6045_ VGND VPWR net1381 s0.data_out\[12\]\[2\] _1943_ _1860_ sg13g2_a21oi_1
XFILLER_26_246 VPWR VGND sg13g2_fill_1
XFILLER_26_279 VPWR VGND sg13g2_decap_8
X_6947_ VGND VPWR net1265 net666 _2751_ _2709_ sg13g2_a21oi_1
X_6878_ _2687_ VPWR _2688_ VGND _2675_ _2684_ sg13g2_o21ai_1
X_7761__259 VPWR VGND net259 sg13g2_tiehi
X_5829_ net1749 VPWR _1745_ VGND net663 _1740_ sg13g2_o21ai_1
XFILLER_1_323 VPWR VGND sg13g2_fill_1
XFILLER_49_305 VPWR VGND sg13g2_fill_2
XFILLER_2_868 VPWR VGND sg13g2_decap_8
XFILLER_45_588 VPWR VGND sg13g2_fill_2
XFILLER_14_920 VPWR VGND sg13g2_fill_1
XFILLER_41_761 VPWR VGND sg13g2_fill_1
XFILLER_9_423 VPWR VGND sg13g2_fill_2
XFILLER_9_489 VPWR VGND sg13g2_fill_2
X_4160_ _3536_ net503 VPWR VGND sg13g2_inv_2
XFILLER_49_850 VPWR VGND sg13g2_decap_8
X_4091_ VPWR _3467_ net457 VGND sg13g2_inv_1
XFILLER_48_371 VPWR VGND sg13g2_fill_1
X_7850_ net163 VGND VPWR _0328_ s0.data_out\[10\]\[4\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_6801_ VPWR _0016_ net642 VGND sg13g2_inv_1
X_4993_ _0991_ net1480 net836 VPWR VGND sg13g2_nand2_1
X_7781_ net237 VGND VPWR _0259_ s0.data_out\[15\]\[2\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_6732_ _2552_ net1271 _2553_ _2554_ VPWR VGND sg13g2_a21o_1
XFILLER_32_750 VPWR VGND sg13g2_fill_1
X_6663_ _2497_ _2496_ net1672 _2490_ net1680 VPWR VGND sg13g2_a22oi_1
XFILLER_17_1025 VPWR VGND sg13g2_decap_4
X_5614_ s0.data_out\[16\]\[7\] s0.data_out\[15\]\[7\] net1421 _1551_ VPWR VGND sg13g2_mux2_1
XFILLER_31_293 VPWR VGND sg13g2_fill_2
X_6594_ _3394_ VPWR _2431_ VGND net471 net1303 sg13g2_o21ai_1
X_8333_ s0.was_valid_out\[27\][0] net2 VPWR VGND sg13g2_buf_1
X_5545_ net1431 net466 _1490_ VPWR VGND sg13g2_and2_1
X_5476_ net1425 net1168 _1425_ VPWR VGND sg13g2_nor2_1
X_4427_ _0130_ _0476_ _0477_ _3404_ net1577 VPWR VGND sg13g2_a22oi_1
X_7215_ VGND VPWR _3360_ _2986_ _0060_ _2991_ sg13g2_a21oi_1
X_7146_ net1240 net1328 _2932_ VPWR VGND sg13g2_nor2b_1
X_4358_ _0415_ _0414_ net1687 _0391_ net1695 VPWR VGND sg13g2_a22oi_1
XFILLER_24_1007 VPWR VGND sg13g2_decap_8
X_4289_ net1578 _3571_ _0356_ VPWR VGND sg13g2_nor2_1
X_7077_ net1596 _2807_ _2867_ VPWR VGND sg13g2_nor2_1
X_6028_ _1929_ _1925_ _1926_ _1928_ VPWR VGND sg13g2_and3_1
XFILLER_27_533 VPWR VGND sg13g2_fill_2
XFILLER_42_503 VPWR VGND sg13g2_decap_8
XFILLER_15_717 VPWR VGND sg13g2_fill_2
XFILLER_23_783 VPWR VGND sg13g2_decap_8
XFILLER_2_687 VPWR VGND sg13g2_decap_8
XFILLER_46_820 VPWR VGND sg13g2_decap_8
X_7809__207 VPWR VGND net207 sg13g2_tiehi
XFILLER_45_341 VPWR VGND sg13g2_fill_2
XFILLER_46_897 VPWR VGND sg13g2_decap_8
XFILLER_45_396 VPWR VGND sg13g2_fill_1
XFILLER_9_253 VPWR VGND sg13g2_decap_8
XFILLER_9_264 VPWR VGND sg13g2_fill_2
X_5330_ _1290_ VPWR _1291_ VGND net1204 _1288_ sg13g2_o21ai_1
XFILLER_47_1018 VPWR VGND sg13g2_decap_8
XFILLER_5_481 VPWR VGND sg13g2_fill_1
X_5261_ _1231_ _1233_ net1674 _1234_ VPWR VGND sg13g2_nand3_1
X_4212_ VGND VPWR net1560 _3575_ _3576_ _3571_ sg13g2_a21oi_1
X_7000_ VGND VPWR _2677_ _2797_ _2798_ net1259 sg13g2_a21oi_1
X_5192_ _0204_ _1167_ _1168_ _3445_ net1617 VPWR VGND sg13g2_a22oi_1
X_4143_ VPWR _3519_ net630 VGND sg13g2_inv_1
X_4074_ _3450_ net497 VPWR VGND sg13g2_inv_2
XFILLER_37_831 VPWR VGND sg13g2_fill_2
X_7902_ net107 VGND VPWR _0036_ s0.was_valid_out\[5\][0] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_7833_ net181 VGND VPWR _0311_ s0.data_out\[11\]\[6\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_7764_ net255 VGND VPWR _0242_ s0.valid_out\[16\][0] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_7899__110 VPWR VGND net110 sg13g2_tiehi
X_6715_ net1176 VPWR _2540_ VGND net398 net1291 sg13g2_o21ai_1
X_4976_ _0974_ net1481 net664 VPWR VGND sg13g2_nand2_1
X_7695_ net330 VGND VPWR _0173_ s0.data_out\[22\]\[0\] clknet_leaf_38_clk sg13g2_dfrbpq_2
XFILLER_20_720 VPWR VGND sg13g2_decap_4
X_6646_ VGND VPWR net1297 _2477_ _2480_ _2479_ sg13g2_a21oi_1
Xclkload6 clkload6/Y clknet_leaf_35_clk VPWR VGND sg13g2_inv_2
XFILLER_20_786 VPWR VGND sg13g2_fill_2
XFILLER_30_1000 VPWR VGND sg13g2_decap_8
X_6577_ _2416_ VPWR _2417_ VGND net1732 net804 sg13g2_o21ai_1
X_5528_ VGND VPWR _1471_ _1475_ _1477_ _1476_ sg13g2_a21oi_1
X_5459_ net1423 net1358 _1408_ VPWR VGND sg13g2_nor2b_1
Xfanout1208 net1210 net1208 VPWR VGND sg13g2_buf_2
Xfanout1219 net1220 net1219 VPWR VGND sg13g2_buf_1
X_7129_ _2915_ net1172 _2914_ VPWR VGND sg13g2_nand2_1
XFILLER_47_606 VPWR VGND sg13g2_decap_4
XFILLER_15_547 VPWR VGND sg13g2_fill_2
XFILLER_6_256 VPWR VGND sg13g2_fill_2
XFILLER_6_245 VPWR VGND sg13g2_fill_1
XFILLER_40_94 VPWR VGND sg13g2_decap_8
XFILLER_3_963 VPWR VGND sg13g2_decap_8
X_7815__200 VPWR VGND net200 sg13g2_tiehi
Xfanout1731 net1732 net1731 VPWR VGND sg13g2_buf_8
Xfanout1720 net1721 net1720 VPWR VGND sg13g2_buf_8
Xfanout1742 net1746 net1742 VPWR VGND sg13g2_buf_8
XFILLER_38_628 VPWR VGND sg13g2_fill_1
XFILLER_19_831 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_15 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_46_672 VPWR VGND sg13g2_decap_4
XFILLER_45_171 VPWR VGND sg13g2_fill_2
X_4830_ _0732_ VPWR _0839_ VGND net1506 _3444_ sg13g2_o21ai_1
X_4761_ _0782_ net1512 _0781_ VPWR VGND sg13g2_nand2b_1
X_7480_ net1208 net1356 _3230_ VPWR VGND sg13g2_nor2b_1
X_4692_ _0716_ _0713_ _0715_ VPWR VGND sg13g2_nand2_1
X_6500_ _2344_ net1300 _2345_ _2346_ VPWR VGND sg13g2_a21o_1
X_6431_ net1609 _2218_ _2287_ VPWR VGND sg13g2_nor2_1
X_6362_ s0.data_out\[10\]\[0\] s0.data_out\[9\]\[0\] net1315 _2220_ VPWR VGND sg13g2_mux2_1
X_5313_ net1452 VPWR _1277_ VGND net1644 net1439 sg13g2_o21ai_1
X_6293_ _0306_ _2166_ _2167_ _3492_ net1611 VPWR VGND sg13g2_a22oi_1
X_5244_ s0.data_out\[19\]\[7\] s0.data_out\[18\]\[7\] net1454 _1217_ VPWR VGND sg13g2_mux2_1
Xhold29 s0.was_valid_out\[6\][0] VPWR VGND net398 sg13g2_dlygate4sd3_1
Xhold18 s0.genblk1\[20\].modules.bubble VPWR VGND net387 sg13g2_dlygate4sd3_1
X_5175_ _0200_ _1154_ _1155_ _3448_ net1606 VPWR VGND sg13g2_a22oi_1
X_4126_ VPWR _3502_ net493 VGND sg13g2_inv_1
XFILLER_29_617 VPWR VGND sg13g2_fill_2
X_4057_ VPWR _3433_ net579 VGND sg13g2_inv_1
XFILLER_37_683 VPWR VGND sg13g2_fill_1
XFILLER_37_672 VPWR VGND sg13g2_fill_1
XFILLER_24_311 VPWR VGND sg13g2_fill_1
X_7816_ net199 VGND VPWR net514 s0.data_out\[12\]\[1\] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_25_856 VPWR VGND sg13g2_fill_1
X_7747_ net274 VGND VPWR _0225_ s0.data_out\[18\]\[4\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_4959_ net1470 net1354 _0957_ VPWR VGND sg13g2_nor2b_1
X_7678_ net349 VGND VPWR net526 s0.data_out\[24\]\[7\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_6629_ _2463_ s0.data_out\[7\]\[3\] net1301 VPWR VGND sg13g2_nand2b_1
XFILLER_0_922 VPWR VGND sg13g2_decap_8
XFILLER_0_999 VPWR VGND sg13g2_decap_8
XFILLER_28_661 VPWR VGND sg13g2_decap_8
XFILLER_43_653 VPWR VGND sg13g2_fill_1
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_37_1017 VPWR VGND sg13g2_decap_8
XFILLER_11_550 VPWR VGND sg13g2_fill_2
Xfanout1550 net1553 net1550 VPWR VGND sg13g2_buf_1
Xfanout1583 net1584 net1583 VPWR VGND sg13g2_buf_8
Xfanout1561 net1562 net1561 VPWR VGND sg13g2_buf_1
Xfanout1572 net1574 net1572 VPWR VGND sg13g2_buf_1
Xfanout1594 net1595 net1594 VPWR VGND sg13g2_buf_1
X_6980_ _2778_ net1255 s0.data_out\[4\]\[1\] VPWR VGND sg13g2_nand2_1
X_5931_ net1194 _3483_ _1838_ VPWR VGND sg13g2_nor2_1
X_5862_ VGND VPWR s0.shift_out\[14\][0] _1772_ _1775_ _1774_ sg13g2_a21oi_1
X_7601_ VGND VPWR net1211 net1167 _3339_ _3338_ sg13g2_a21oi_1
X_4813_ net1643 net1490 _0825_ VPWR VGND sg13g2_nor2b_1
X_5793_ VGND VPWR net1402 s0.data_out\[14\]\[2\] _1715_ _1644_ sg13g2_a21oi_1
XFILLER_34_697 VPWR VGND sg13g2_fill_1
X_7532_ _3256_ _3257_ _3282_ VPWR VGND sg13g2_nor2b_1
X_4744_ VGND VPWR _0651_ _0764_ _0765_ net1512 sg13g2_a21oi_1
X_7896__113 VPWR VGND net113 sg13g2_tiehi
X_7463_ net1584 _3209_ _0085_ VPWR VGND sg13g2_nor2_1
X_4675_ net1524 VPWR _0702_ VGND _0669_ _0701_ sg13g2_o21ai_1
X_7394_ net1221 net1338 _3156_ VPWR VGND sg13g2_nor2b_1
X_6414_ _2261_ _2259_ net1682 _2272_ VPWR VGND sg13g2_a21o_1
X_6345_ VGND VPWR net1638 _3402_ _0321_ _2204_ sg13g2_a21oi_1
X_6276_ VGND VPWR _2153_ _2151_ net1673 sg13g2_or2_1
XFILLER_1_719 VPWR VGND sg13g2_decap_8
XFILLER_0_229 VPWR VGND sg13g2_fill_1
X_5227_ _1200_ net1454 net487 VPWR VGND sg13g2_nand2_1
X_5158_ VGND VPWR _1137_ _1141_ _0196_ _1142_ sg13g2_a21oi_1
XFILLER_29_436 VPWR VGND sg13g2_decap_4
XFILLER_45_907 VPWR VGND sg13g2_decap_8
X_4109_ VPWR _3485_ net757 VGND sg13g2_inv_1
X_5089_ VGND VPWR net1472 _1071_ _1074_ _1073_ sg13g2_a21oi_1
XFILLER_12_336 VPWR VGND sg13g2_decap_4
XFILLER_4_557 VPWR VGND sg13g2_fill_1
X_7812__203 VPWR VGND net203 sg13g2_tiehi
XFILLER_0_796 VPWR VGND sg13g2_decap_8
XFILLER_48_767 VPWR VGND sg13g2_decap_8
XFILLER_29_992 VPWR VGND sg13g2_decap_8
XFILLER_44_995 VPWR VGND sg13g2_decap_8
XFILLER_43_494 VPWR VGND sg13g2_fill_1
Xhold307 s0.was_valid_out\[27\][0] VPWR VGND net676 sg13g2_dlygate4sd3_1
XFILLER_7_362 VPWR VGND sg13g2_fill_1
X_4460_ _0504_ VPWR _0505_ VGND net1529 _3420_ sg13g2_o21ai_1
Xhold318 s0.data_out\[11\]\[6\] VPWR VGND net687 sg13g2_dlygate4sd3_1
X_4391_ VGND VPWR _3620_ _0447_ _0448_ net1544 sg13g2_a21oi_1
Xhold329 s0.data_out\[24\]\[4\] VPWR VGND net698 sg13g2_dlygate4sd3_1
X_6130_ VGND VPWR net1380 _2016_ _2019_ _2018_ sg13g2_a21oi_1
X_6061_ _0286_ _1954_ _1955_ _3483_ net1629 VPWR VGND sg13g2_a22oi_1
X_5012_ _1010_ net1480 s0.data_out\[20\]\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_38_244 VPWR VGND sg13g2_fill_1
Xfanout1391 net1396 net1391 VPWR VGND sg13g2_buf_8
Xfanout1380 net1381 net1380 VPWR VGND sg13g2_buf_8
XFILLER_26_406 VPWR VGND sg13g2_fill_1
X_6963_ VGND VPWR net1634 net1267 _2764_ net1258 sg13g2_a21oi_1
X_6894_ VGND VPWR _2704_ _2695_ net1660 sg13g2_or2_1
X_5914_ net1390 net577 _1825_ VPWR VGND sg13g2_and2_1
XFILLER_35_962 VPWR VGND sg13g2_decap_8
XFILLER_22_623 VPWR VGND sg13g2_fill_2
X_5845_ _1758_ net577 net1408 VPWR VGND sg13g2_nand2b_1
X_5776_ VGND VPWR _1694_ _1696_ _1701_ net1685 sg13g2_a21oi_1
X_7515_ _3265_ net1223 _3264_ VPWR VGND sg13g2_nand2b_1
X_4727_ VGND VPWR net1513 _0745_ _0748_ _0747_ sg13g2_a21oi_1
X_4658_ net1182 _3436_ _0689_ VPWR VGND sg13g2_nor2_1
X_7446_ _3200_ net1718 _3201_ VPWR VGND _3143_ sg13g2_nand3b_1
X_4589_ net1511 net1353 _0622_ VPWR VGND sg13g2_nor2b_1
X_7377_ s0.data_out\[2\]\[6\] s0.data_out\[1\]\[6\] net1224 _3139_ VPWR VGND sg13g2_mux2_1
X_6328_ net441 _2195_ _2196_ VPWR VGND sg13g2_nor2_1
XFILLER_27_1027 VPWR VGND sg13g2_fill_2
X_6259_ VGND VPWR _2136_ _2132_ net1653 sg13g2_or2_1
XFILLER_44_214 VPWR VGND sg13g2_fill_1
XFILLER_44_203 VPWR VGND sg13g2_fill_1
XFILLER_26_984 VPWR VGND sg13g2_decap_8
XFILLER_41_954 VPWR VGND sg13g2_decap_8
XFILLER_40_431 VPWR VGND sg13g2_fill_2
XFILLER_5_888 VPWR VGND sg13g2_fill_1
XFILLER_0_571 VPWR VGND sg13g2_fill_1
XFILLER_48_564 VPWR VGND sg13g2_decap_8
X_7747__274 VPWR VGND net274 sg13g2_tiehi
XFILLER_16_494 VPWR VGND sg13g2_fill_2
X_5630_ _1564_ _1565_ _1567_ VPWR VGND _1566_ sg13g2_nand3b_1
X_5561_ _1502_ net1745 _1503_ VPWR VGND _1446_ sg13g2_nand3b_1
X_7893__116 VPWR VGND net116 sg13g2_tiehi
X_4512_ net1519 net1343 _0557_ VPWR VGND sg13g2_nor2b_1
X_5492_ _1441_ net1434 s0.data_out\[16\]\[6\] VPWR VGND sg13g2_nand2_1
X_7300_ net1228 s0.data_out\[2\]\[1\] _3072_ VPWR VGND sg13g2_and2_1
Xhold115 _0343_ VPWR VGND net484 sg13g2_dlygate4sd3_1
Xhold104 _0119_ VPWR VGND net473 sg13g2_dlygate4sd3_1
X_7231_ _3004_ VPWR _3005_ VGND net1190 _3002_ sg13g2_o21ai_1
Xhold126 s0.data_out\[16\]\[1\] VPWR VGND net495 sg13g2_dlygate4sd3_1
X_4443_ net1184 VPWR _0491_ VGND s0.was_valid_out\[24\][0] net1542 sg13g2_o21ai_1
Xhold148 s0.data_out\[26\]\[4\] VPWR VGND net517 sg13g2_dlygate4sd3_1
Xhold159 _0252_ VPWR VGND net528 sg13g2_dlygate4sd3_1
Xhold137 _0055_ VPWR VGND net506 sg13g2_dlygate4sd3_1
X_4374_ _0431_ _0430_ net1647 _0423_ net1658 VPWR VGND sg13g2_a22oi_1
X_7162_ _2947_ VPWR _2948_ VGND _2899_ _2908_ sg13g2_o21ai_1
X_7093_ net1240 net1348 _2879_ VPWR VGND sg13g2_nor2b_1
X_6113_ VGND VPWR _1882_ _2001_ _2002_ net1377 sg13g2_a21oi_1
X_6044_ VPWR _0282_ _1942_ VGND sg13g2_inv_1
XFILLER_39_531 VPWR VGND sg13g2_fill_1
X_6946_ VPWR _0032_ net519 VGND sg13g2_inv_1
XFILLER_26_258 VPWR VGND sg13g2_fill_2
XFILLER_23_932 VPWR VGND sg13g2_fill_2
X_6877_ _2687_ net1688 _2683_ VPWR VGND sg13g2_nand2_1
X_5828_ _1742_ _1743_ _1744_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_998 VPWR VGND sg13g2_decap_8
X_5759_ net1404 net1341 _1684_ VPWR VGND sg13g2_nor2b_1
X_7429_ _3187_ VPWR _3188_ VGND net1719 net756 sg13g2_o21ai_1
XFILLER_2_847 VPWR VGND sg13g2_decap_8
XFILLER_49_328 VPWR VGND sg13g2_fill_1
XFILLER_18_715 VPWR VGND sg13g2_fill_1
XFILLER_1_880 VPWR VGND sg13g2_decap_8
X_4090_ VPWR _3466_ net527 VGND sg13g2_inv_1
XFILLER_36_501 VPWR VGND sg13g2_decap_8
XFILLER_36_523 VPWR VGND sg13g2_fill_1
X_6800_ _2620_ VPWR _2621_ VGND net1731 net641 sg13g2_o21ai_1
X_4992_ VGND VPWR net1483 _0987_ _0990_ _0989_ sg13g2_a21oi_1
XFILLER_23_206 VPWR VGND sg13g2_fill_1
X_7780_ net238 VGND VPWR net703 s0.data_out\[15\]\[1\] clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_17_1004 VPWR VGND sg13g2_decap_8
X_6731_ net1270 net1353 _2553_ VPWR VGND sg13g2_nor2b_1
X_6662_ VGND VPWR net1296 _2493_ _2496_ _2495_ sg13g2_a21oi_1
XFILLER_31_261 VPWR VGND sg13g2_fill_2
XFILLER_32_773 VPWR VGND sg13g2_fill_2
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
X_7760__260 VPWR VGND net260 sg13g2_tiehi
X_5613_ _1550_ net1420 net564 VPWR VGND sg13g2_nand2_1
X_6593_ _2427_ _2429_ _2430_ VPWR VGND sg13g2_nor2_1
X_5544_ VPWR _0235_ _1489_ VGND sg13g2_inv_1
X_5475_ _1423_ VPWR _1424_ VGND net1432 _3463_ sg13g2_o21ai_1
X_4426_ net1577 _0448_ _0477_ VPWR VGND sg13g2_nor2_1
X_7214_ net1718 VPWR _2991_ VGND _2988_ _2990_ sg13g2_o21ai_1
X_7145_ s0.data_out\[4\]\[7\] s0.data_out\[3\]\[7\] net1246 _2931_ VPWR VGND sg13g2_mux2_1
X_4357_ VGND VPWR net1551 _0411_ _0414_ _0413_ sg13g2_a21oi_1
X_4288_ net1560 VPWR _0355_ VGND _3574_ _0354_ sg13g2_o21ai_1
X_7076_ net1258 VPWR _2866_ VGND _2804_ _2865_ sg13g2_o21ai_1
X_6027_ VGND VPWR _1928_ _1924_ net1655 sg13g2_or2_1
XFILLER_39_350 VPWR VGND sg13g2_fill_1
XFILLER_27_578 VPWR VGND sg13g2_fill_1
X_6929_ net1261 s0.data_out\[5\]\[1\] _2737_ VPWR VGND sg13g2_and2_1
XFILLER_7_917 VPWR VGND sg13g2_fill_1
XFILLER_1_154 VPWR VGND sg13g2_fill_2
XFILLER_46_876 VPWR VGND sg13g2_decap_8
XFILLER_18_556 VPWR VGND sg13g2_fill_1
XFILLER_33_548 VPWR VGND sg13g2_fill_1
XFILLER_9_232 VPWR VGND sg13g2_fill_2
X_7744__277 VPWR VGND net277 sg13g2_tiehi
XFILLER_10_990 VPWR VGND sg13g2_decap_8
XFILLER_6_994 VPWR VGND sg13g2_decap_8
X_5260_ _1233_ net1199 _1232_ VPWR VGND sg13g2_nand2_1
X_4211_ _3573_ net1546 _3574_ _3575_ VPWR VGND sg13g2_a21o_1
X_5191_ net1617 _1112_ _1168_ VPWR VGND sg13g2_nor2_1
X_4142_ VPWR _3518_ net653 VGND sg13g2_inv_1
X_4073_ VPWR _3449_ net591 VGND sg13g2_inv_1
XFILLER_48_180 VPWR VGND sg13g2_fill_1
X_7901_ net108 VGND VPWR _0035_ s0.data_out\[6\]\[7\] clknet_leaf_12_clk sg13g2_dfrbpq_2
X_7832_ net182 VGND VPWR net640 s0.data_out\[11\]\[5\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_4975_ VPWR VGND _0972_ _0965_ _0964_ net1573 _0973_ _0956_ sg13g2_a221oi_1
X_7763_ net257 VGND VPWR _0241_ s0.was_valid_out\[16\][0] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_24_559 VPWR VGND sg13g2_decap_4
X_6714_ net1277 _2533_ _2539_ VPWR VGND sg13g2_nor2_1
X_7694_ net331 VGND VPWR _0172_ s0.shift_out\[22\][0] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_6645_ VGND VPWR _2351_ _2478_ _2479_ net1296 sg13g2_a21oi_1
Xclkload7 clknet_leaf_29_clk clkload7/X VPWR VGND sg13g2_buf_8
X_6576_ _2375_ _2415_ net1732 _2416_ VPWR VGND sg13g2_nand3_1
X_5527_ _1393_ VPWR _1476_ VGND _1448_ _1451_ sg13g2_o21ai_1
X_5458_ _1407_ net1206 _1406_ VPWR VGND sg13g2_nand2_1
Xfanout1209 net1210 net1209 VPWR VGND sg13g2_buf_8
XFILLER_8_1024 VPWR VGND sg13g2_decap_4
X_5389_ _1350_ _1349_ net1674 _1342_ net1684 VPWR VGND sg13g2_a22oi_1
X_4409_ net1551 VPWR _0464_ VGND _0395_ _0463_ sg13g2_o21ai_1
X_7128_ _2826_ VPWR _2914_ VGND net1254 _3536_ sg13g2_o21ai_1
X_7059_ net1173 _3533_ _2853_ VPWR VGND sg13g2_nor2_1
XFILLER_42_312 VPWR VGND sg13g2_fill_2
XFILLER_28_887 VPWR VGND sg13g2_fill_1
XFILLER_43_879 VPWR VGND sg13g2_decap_8
XFILLER_30_518 VPWR VGND sg13g2_fill_2
XFILLER_7_714 VPWR VGND sg13g2_fill_2
XFILLER_7_736 VPWR VGND sg13g2_fill_2
X_7698__327 VPWR VGND net327 sg13g2_tiehi
XFILLER_3_942 VPWR VGND sg13g2_decap_8
XFILLER_2_441 VPWR VGND sg13g2_decap_4
Xfanout1721 net1724 net1721 VPWR VGND sg13g2_buf_8
Xfanout1732 net1733 net1732 VPWR VGND sg13g2_buf_8
Xfanout1710 net1713 net1710 VPWR VGND sg13g2_buf_8
Xfanout1743 net1746 net1743 VPWR VGND sg13g2_buf_8
XFILLER_46_640 VPWR VGND sg13g2_fill_1
Xheichips25_top_sorter_16 VPWR VGND uio_oe[7] sg13g2_tielo
XFILLER_46_695 VPWR VGND sg13g2_decap_8
XFILLER_45_183 VPWR VGND sg13g2_fill_1
XFILLER_33_334 VPWR VGND sg13g2_fill_2
X_4760_ VGND VPWR net1494 _0780_ _0781_ _0779_ sg13g2_a21oi_1
X_4691_ net1181 VPWR _0715_ VGND s0.was_valid_out\[22\][0] net1516 sg13g2_o21ai_1
X_6430_ net1319 VPWR _2286_ VGND _2213_ _2285_ sg13g2_o21ai_1
X_6361_ VGND VPWR net1319 _2216_ _2219_ _2218_ sg13g2_a21oi_1
X_5312_ _0216_ _1275_ _1276_ _3451_ net1618 VPWR VGND sg13g2_a22oi_1
X_6292_ net1611 _2100_ _2167_ VPWR VGND sg13g2_nor2_1
X_5243_ _1216_ net1455 net805 VPWR VGND sg13g2_nand2_1
Xhold19 s0.genblk1\[10\].modules.bubble VPWR VGND net388 sg13g2_dlygate4sd3_1
X_5174_ net1606 _1096_ _1155_ VPWR VGND sg13g2_nor2_1
X_4125_ VPWR _3501_ net522 VGND sg13g2_inv_1
XFILLER_29_629 VPWR VGND sg13g2_decap_8
X_4056_ VPWR _3432_ net662 VGND sg13g2_inv_1
XFILLER_37_662 VPWR VGND sg13g2_fill_1
XFILLER_36_161 VPWR VGND sg13g2_fill_2
X_7815_ net200 VGND VPWR _0293_ s0.data_out\[12\]\[0\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_7746_ net275 VGND VPWR net488 s0.data_out\[18\]\[3\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_4958_ _0955_ VPWR _0956_ VGND net1178 _0953_ sg13g2_o21ai_1
XFILLER_24_389 VPWR VGND sg13g2_fill_2
X_7677_ net350 VGND VPWR net490 s0.data_out\[24\]\[6\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_4889_ _0898_ net1500 _0897_ VPWR VGND sg13g2_nand2b_1
X_6628_ _2460_ net1283 _2461_ _2462_ VPWR VGND sg13g2_a21o_1
X_6559_ net1608 _2332_ _2403_ VPWR VGND sg13g2_nor2_1
XFILLER_0_901 VPWR VGND sg13g2_decap_8
XFILLER_0_978 VPWR VGND sg13g2_decap_8
XFILLER_48_949 VPWR VGND sg13g2_decap_8
XFILLER_19_63 VPWR VGND sg13g2_fill_2
XFILLER_28_640 VPWR VGND sg13g2_fill_2
XFILLER_27_161 VPWR VGND sg13g2_fill_1
XFILLER_16_857 VPWR VGND sg13g2_fill_1
XFILLER_43_665 VPWR VGND sg13g2_fill_1
XFILLER_42_131 VPWR VGND sg13g2_decap_4
XFILLER_16_879 VPWR VGND sg13g2_decap_8
XFILLER_31_805 VPWR VGND sg13g2_fill_1
XFILLER_42_175 VPWR VGND sg13g2_fill_1
XFILLER_11_573 VPWR VGND sg13g2_fill_2
X_7889__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_38_404 VPWR VGND sg13g2_fill_2
Xfanout1540 net771 net1540 VPWR VGND sg13g2_buf_8
Xfanout1551 net1553 net1551 VPWR VGND sg13g2_buf_8
Xfanout1584 net1588 net1584 VPWR VGND sg13g2_buf_8
Xfanout1562 s0.shift_out\[27\][0] net1562 VPWR VGND sg13g2_buf_2
XFILLER_18_4 VPWR VGND sg13g2_decap_8
Xfanout1573 net1574 net1573 VPWR VGND sg13g2_buf_8
XFILLER_38_459 VPWR VGND sg13g2_fill_1
Xfanout1595 net1603 net1595 VPWR VGND sg13g2_buf_8
XFILLER_46_470 VPWR VGND sg13g2_fill_1
X_5930_ VPWR _0273_ _1837_ VGND sg13g2_inv_1
XFILLER_18_183 VPWR VGND sg13g2_fill_1
X_7600_ VGND VPWR net1215 net433 _3338_ net1211 sg13g2_a21oi_1
X_5861_ VGND VPWR _1652_ _1773_ _1774_ net1403 sg13g2_a21oi_1
X_4812_ net1498 VPWR _0824_ VGND net1643 net1482 sg13g2_o21ai_1
X_5792_ _0258_ _1713_ _1714_ _3475_ net1626 VPWR VGND sg13g2_a22oi_1
X_7531_ _3259_ _3280_ _3281_ VPWR VGND sg13g2_nor2b_1
X_4743_ _0764_ net552 net1516 VPWR VGND sg13g2_nand2b_1
X_7462_ _3213_ _3214_ _0084_ VPWR VGND sg13g2_nor2_1
XFILLER_30_860 VPWR VGND sg13g2_fill_1
X_6413_ _2271_ net1676 _2269_ VPWR VGND sg13g2_nand2_1
X_4674_ net1508 net610 _0701_ VPWR VGND sg13g2_and2_1
X_7393_ s0.data_out\[2\]\[5\] s0.data_out\[1\]\[5\] net1226 _3155_ VPWR VGND sg13g2_mux2_1
X_6344_ net1638 net1333 _2204_ VPWR VGND sg13g2_nor2_1
X_6275_ _2151_ net1673 _2144_ _2152_ VPWR VGND sg13g2_a21o_1
X_5226_ _1184_ VPWR _1199_ VGND net1706 _1191_ sg13g2_o21ai_1
X_5157_ VGND VPWR _1142_ net1567 net387 sg13g2_or2_1
X_5088_ VGND VPWR _0950_ _1072_ _1073_ net1472 sg13g2_a21oi_1
XFILLER_29_448 VPWR VGND sg13g2_decap_4
X_4108_ _3484_ net574 VPWR VGND sg13g2_inv_2
XFILLER_38_993 VPWR VGND sg13g2_decap_8
X_4039_ _3415_ net1701 VPWR VGND sg13g2_inv_2
XFILLER_25_676 VPWR VGND sg13g2_fill_1
XFILLER_24_186 VPWR VGND sg13g2_fill_2
X_7805__211 VPWR VGND net211 sg13g2_tiehi
XFILLER_40_657 VPWR VGND sg13g2_fill_2
X_7729_ net293 VGND VPWR _0207_ s0.genblk1\[18\].modules.bubble clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
XFILLER_48_746 VPWR VGND sg13g2_decap_8
XFILLER_0_775 VPWR VGND sg13g2_decap_8
XFILLER_29_971 VPWR VGND sg13g2_decap_8
XFILLER_28_492 VPWR VGND sg13g2_decap_8
XFILLER_44_974 VPWR VGND sg13g2_decap_8
XFILLER_15_164 VPWR VGND sg13g2_fill_2
XFILLER_16_698 VPWR VGND sg13g2_fill_2
XFILLER_31_624 VPWR VGND sg13g2_fill_2
Xhold308 _0109_ VPWR VGND net677 sg13g2_dlygate4sd3_1
Xhold319 _2183_ VPWR VGND net688 sg13g2_dlygate4sd3_1
X_4390_ _0447_ s0.data_out\[25\]\[5\] net1556 VPWR VGND sg13g2_nand2b_1
X_6060_ net1628 _1905_ _1955_ VPWR VGND sg13g2_nor2_1
X_5011_ _1009_ net1673 _1008_ VPWR VGND sg13g2_nand2_1
Xfanout1370 net1371 net1370 VPWR VGND sg13g2_buf_8
Xfanout1392 net1393 net1392 VPWR VGND sg13g2_buf_8
Xfanout1381 s0.shift_out\[12\][0] net1381 VPWR VGND sg13g2_buf_1
X_6962_ _2761_ _2762_ _2763_ VPWR VGND sg13g2_nor2_1
X_6893_ _2703_ _2702_ net1650 _2695_ net1660 VPWR VGND sg13g2_a22oi_1
X_5913_ VPWR _0269_ net658 VGND sg13g2_inv_1
X_5844_ _1755_ net1390 _1756_ _1757_ VPWR VGND sg13g2_a21o_1
X_7514_ VGND VPWR net1213 _3262_ _3264_ _3263_ sg13g2_a21oi_1
X_5775_ VPWR _1700_ _1699_ VGND sg13g2_inv_1
X_4726_ VGND VPWR _0636_ _0746_ _0747_ net1514 sg13g2_a21oi_1
X_4657_ VPWR _0149_ _0688_ VGND sg13g2_inv_1
X_7445_ net1230 VPWR _3200_ VGND _3140_ _3199_ sg13g2_o21ai_1
X_7376_ _3129_ _3137_ _3138_ VPWR VGND _3128_ sg13g2_nand3b_1
X_6327_ _2190_ VPWR _2195_ VGND net1324 _2078_ sg13g2_o21ai_1
XFILLER_1_517 VPWR VGND sg13g2_fill_1
X_4588_ s0.data_out\[24\]\[1\] s0.data_out\[23\]\[1\] net1515 _0621_ VPWR VGND sg13g2_mux2_1
X_7638__48 VPWR VGND net48 sg13g2_tiehi
XFILLER_27_1006 VPWR VGND sg13g2_decap_8
X_6258_ net1663 _2125_ _2135_ VPWR VGND sg13g2_nor2_1
X_6189_ net1380 VPWR _2071_ VGND _2008_ _2070_ sg13g2_o21ai_1
X_5209_ VGND VPWR _1068_ _1181_ _1182_ net1463 sg13g2_a21oi_1
XFILLER_45_716 VPWR VGND sg13g2_fill_1
XFILLER_29_278 VPWR VGND sg13g2_fill_2
XFILLER_44_259 VPWR VGND sg13g2_fill_1
XFILLER_41_933 VPWR VGND sg13g2_decap_8
X_7879__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_0_550 VPWR VGND sg13g2_decap_4
XFILLER_48_543 VPWR VGND sg13g2_decap_8
X_7886__124 VPWR VGND net124 sg13g2_tiehi
XFILLER_36_738 VPWR VGND sg13g2_fill_1
XFILLER_35_259 VPWR VGND sg13g2_fill_1
XFILLER_44_771 VPWR VGND sg13g2_fill_2
XFILLER_32_944 VPWR VGND sg13g2_fill_1
X_5560_ net1440 VPWR _1502_ VGND _1443_ _1501_ sg13g2_o21ai_1
X_4511_ _0553_ _0555_ net1671 _0556_ VPWR VGND sg13g2_nand3_1
X_5491_ VGND VPWR net1440 _1437_ _1440_ _1439_ sg13g2_a21oi_1
X_4442_ net1519 _0485_ _0490_ VPWR VGND sg13g2_nor2_1
X_7230_ _3004_ net1190 _3003_ VPWR VGND sg13g2_nand2_1
Xhold116 s0.data_out\[9\]\[2\] VPWR VGND net485 sg13g2_dlygate4sd3_1
Xhold105 s0.shift_out\[14\][0] VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold138 s0.was_valid_out\[0\][0] VPWR VGND net507 sg13g2_dlygate4sd3_1
Xhold149 s0.data_out\[6\]\[4\] VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold127 _0246_ VPWR VGND net496 sg13g2_dlygate4sd3_1
X_4373_ VGND VPWR net1550 _0427_ _0430_ _0429_ sg13g2_a21oi_1
X_7161_ _2947_ _2943_ _2944_ _2946_ VPWR VGND sg13g2_and3_1
X_7092_ s0.data_out\[4\]\[2\] s0.data_out\[3\]\[2\] net1246 _2878_ VPWR VGND sg13g2_mux2_1
X_6112_ _2001_ s0.data_out\[11\]\[3\] net1386 VPWR VGND sg13g2_nand2b_1
X_6043_ _1941_ VPWR _1942_ VGND net1740 net577 sg13g2_o21ai_1
XFILLER_2_1008 VPWR VGND sg13g2_decap_8
XFILLER_26_204 VPWR VGND sg13g2_decap_4
X_6945_ _2749_ VPWR _2750_ VGND net1730 net518 sg13g2_o21ai_1
XFILLER_22_421 VPWR VGND sg13g2_fill_1
X_6876_ _2667_ _2676_ _2684_ _2685_ _2686_ VPWR VGND sg13g2_nor4_1
X_5827_ net1195 VPWR _1743_ VGND net416 net1411 sg13g2_o21ai_1
XFILLER_23_977 VPWR VGND sg13g2_decap_8
X_7802__214 VPWR VGND net214 sg13g2_tiehi
X_5758_ s0.data_out\[15\]\[5\] s0.data_out\[14\]\[5\] net1410 _1683_ VPWR VGND sg13g2_mux2_1
X_4709_ _0730_ net1513 _0729_ VPWR VGND sg13g2_nand2b_1
X_7428_ _3186_ VPWR _3187_ VGND net1188 _3185_ sg13g2_o21ai_1
X_5689_ net1630 _1555_ _1618_ VPWR VGND sg13g2_nor2_1
XFILLER_2_826 VPWR VGND sg13g2_decap_8
X_7359_ net1217 net1357 _3121_ VPWR VGND sg13g2_nor2b_1
XFILLER_40_1025 VPWR VGND sg13g2_decap_4
XFILLER_27_96 VPWR VGND sg13g2_fill_2
XFILLER_32_218 VPWR VGND sg13g2_fill_2
XFILLER_43_40 VPWR VGND sg13g2_fill_2
XFILLER_41_752 VPWR VGND sg13g2_fill_2
XFILLER_43_73 VPWR VGND sg13g2_fill_2
XFILLER_14_988 VPWR VGND sg13g2_decap_8
XFILLER_0_391 VPWR VGND sg13g2_decap_4
XFILLER_49_885 VPWR VGND sg13g2_decap_8
X_4991_ VGND VPWR _0867_ _0988_ _0989_ net1483 sg13g2_a21oi_1
XFILLER_23_229 VPWR VGND sg13g2_fill_2
X_6730_ _2551_ VPWR _2552_ VGND net1278 _3514_ sg13g2_o21ai_1
X_6661_ VGND VPWR _2369_ _2494_ _2495_ net1296 sg13g2_a21oi_1
XFILLER_20_914 VPWR VGND sg13g2_fill_2
X_6592_ net471 net1292 _2429_ VPWR VGND sg13g2_nor2_1
X_5612_ VPWR VGND net1692 _1541_ _1548_ net1697 _1549_ _1524_ sg13g2_a221oi_1
XFILLER_9_981 VPWR VGND sg13g2_decap_8
X_5543_ _1488_ VPWR _1489_ VGND net1742 net705 sg13g2_o21ai_1
X_5474_ _1423_ net1432 net466 VPWR VGND sg13g2_nand2_1
X_4425_ net1545 VPWR _0476_ VGND _0445_ _0475_ sg13g2_o21ai_1
X_7213_ _2990_ _2987_ _2989_ VPWR VGND sg13g2_nand2_1
X_4356_ VGND VPWR _3590_ _0412_ _0413_ net1551 sg13g2_a21oi_1
X_7144_ _2930_ net1247 net604 VPWR VGND sg13g2_nand2_1
XFILLER_48_29 VPWR VGND sg13g2_fill_1
XFILLER_48_18 VPWR VGND sg13g2_fill_2
X_4287_ net1546 s0.data_out\[26\]\[1\] _0354_ VPWR VGND sg13g2_and2_1
X_7075_ net1173 _3531_ _2865_ VPWR VGND sg13g2_nor2_1
X_6026_ net1655 _1924_ _1927_ VPWR VGND sg13g2_nor2_1
X_6928_ VPWR _0028_ _2736_ VGND sg13g2_inv_1
X_6859_ _2668_ VPWR _2669_ VGND net1266 _3522_ sg13g2_o21ai_1
XFILLER_23_752 VPWR VGND sg13g2_fill_1
XFILLER_13_21 VPWR VGND sg13g2_fill_2
XFILLER_22_295 VPWR VGND sg13g2_fill_2
X_7737__285 VPWR VGND net285 sg13g2_tiehi
XFILLER_46_800 VPWR VGND sg13g2_fill_2
XFILLER_46_855 VPWR VGND sg13g2_decap_8
X_7883__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_14_785 VPWR VGND sg13g2_fill_1
XFILLER_6_973 VPWR VGND sg13g2_decap_8
X_4210_ net1546 net1352 _3574_ VPWR VGND sg13g2_nor2b_1
X_5190_ net1474 VPWR _1167_ VGND _1109_ _1166_ sg13g2_o21ai_1
X_4141_ VPWR _3517_ net414 VGND sg13g2_inv_1
X_4072_ VPWR _3448_ net664 VGND sg13g2_inv_1
XFILLER_49_682 VPWR VGND sg13g2_decap_8
X_7900_ net109 VGND VPWR _0034_ s0.data_out\[6\]\[6\] clknet_leaf_13_clk sg13g2_dfrbpq_2
XFILLER_37_866 VPWR VGND sg13g2_fill_2
X_7831_ net183 VGND VPWR net788 s0.data_out\[11\]\[4\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_24_505 VPWR VGND sg13g2_fill_2
XFILLER_24_516 VPWR VGND sg13g2_fill_2
X_7762_ net258 VGND VPWR _0240_ s0.data_out\[17\]\[7\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_4974_ net1570 _0971_ _0972_ VPWR VGND sg13g2_and2_1
X_6713_ net398 net1281 _2538_ VPWR VGND sg13g2_nor2_1
X_7693_ net332 VGND VPWR _0171_ s0.genblk1\[21\].modules.bubble clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_6644_ _2478_ net414 net1303 VPWR VGND sg13g2_nand2b_1
Xclkload8 VPWR clkload8/Y clknet_leaf_17_clk VGND sg13g2_inv_1
X_6575_ net1309 VPWR _2415_ VGND _2371_ _2414_ sg13g2_o21ai_1
X_5526_ VGND VPWR _1460_ _1468_ _1475_ _1452_ sg13g2_a21oi_1
X_5457_ s0.data_out\[16\]\[0\] s0.data_out\[17\]\[0\] net1443 _1406_ VPWR VGND sg13g2_mux2_1
X_4408_ net1186 _3421_ _0463_ VPWR VGND sg13g2_nor2_1
XFILLER_8_1003 VPWR VGND sg13g2_decap_8
X_5388_ VGND VPWR net1450 _1346_ _1349_ _1348_ sg13g2_a21oi_1
X_4339_ _0394_ net1536 _0395_ _0396_ VPWR VGND sg13g2_a21o_1
X_7127_ _2913_ net1249 _2912_ VPWR VGND sg13g2_nand2b_1
X_7058_ _0042_ _2851_ _2852_ _3529_ net1590 VPWR VGND sg13g2_a22oi_1
X_6009_ _1910_ net1684 _1898_ VPWR VGND sg13g2_xnor2_1
XFILLER_15_549 VPWR VGND sg13g2_fill_1
XFILLER_11_744 VPWR VGND sg13g2_decap_4
XFILLER_11_755 VPWR VGND sg13g2_fill_1
XFILLER_6_258 VPWR VGND sg13g2_fill_1
XFILLER_3_921 VPWR VGND sg13g2_decap_8
XFILLER_2_420 VPWR VGND sg13g2_fill_1
XFILLER_3_998 VPWR VGND sg13g2_decap_8
Xfanout1700 ui_in[2] net1700 VPWR VGND sg13g2_buf_8
Xfanout1722 net1723 net1722 VPWR VGND sg13g2_buf_8
Xfanout1711 net1713 net1711 VPWR VGND sg13g2_buf_8
Xfanout1733 net1751 net1733 VPWR VGND sg13g2_buf_8
Xfanout1744 net1746 net1744 VPWR VGND sg13g2_buf_8
X_7750__271 VPWR VGND net271 sg13g2_tiehi
Xheichips25_top_sorter_17 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_45_173 VPWR VGND sg13g2_fill_1
X_4690_ net1493 _0710_ _0714_ VPWR VGND sg13g2_nor2_1
X_6360_ VGND VPWR _2095_ _2217_ _2218_ net1320 sg13g2_a21oi_1
X_5311_ net1618 _1221_ _1276_ VPWR VGND sg13g2_nor2_1
X_6291_ net1365 VPWR _2166_ VGND _2097_ _2165_ sg13g2_o21ai_1
X_5242_ VGND VPWR net1461 _1212_ _1215_ _1214_ sg13g2_a21oi_1
X_5173_ net1475 VPWR _1154_ VGND _1093_ _1153_ sg13g2_o21ai_1
XFILLER_29_619 VPWR VGND sg13g2_fill_1
X_4124_ VPWR _3500_ net523 VGND sg13g2_inv_1
Xinput1 uio_in[1] net1 VPWR VGND sg13g2_buf_2
X_4055_ VPWR _3431_ net481 VGND sg13g2_inv_1
X_7814_ net201 VGND VPWR _0292_ s0.shift_out\[12\][0] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_7745_ net276 VGND VPWR _0223_ s0.data_out\[18\]\[2\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_4957_ _0955_ net1178 _0954_ VPWR VGND sg13g2_nand2_1
X_7676_ net351 VGND VPWR _0154_ s0.data_out\[24\]\[5\] clknet_leaf_43_clk sg13g2_dfrbpq_2
X_4888_ VGND VPWR net1486 _0896_ _0897_ _0894_ sg13g2_a21oi_1
X_6627_ net1283 net1347 _2461_ VPWR VGND sg13g2_nor2b_1
X_6558_ net1305 VPWR _2402_ VGND _2329_ _2401_ sg13g2_o21ai_1
X_5509_ _1343_ VPWR _1458_ VGND net1445 _3467_ sg13g2_o21ai_1
X_6489_ net1295 net1359 _2335_ VPWR VGND sg13g2_nor2b_1
XFILLER_10_66 VPWR VGND sg13g2_fill_1
XFILLER_0_957 VPWR VGND sg13g2_decap_8
XFILLER_48_928 VPWR VGND sg13g2_decap_8
X_7734__288 VPWR VGND net288 sg13g2_tiehi
Xclkbuf_leaf_39_clk clknet_3_1__leaf_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_30_349 VPWR VGND sg13g2_decap_8
XFILLER_11_585 VPWR VGND sg13g2_fill_1
XFILLER_7_578 VPWR VGND sg13g2_fill_1
XFILLER_3_784 VPWR VGND sg13g2_decap_8
XFILLER_2_283 VPWR VGND sg13g2_fill_2
XFILLER_2_294 VPWR VGND sg13g2_fill_2
Xfanout1541 s0.valid_out\[25\][0] net1541 VPWR VGND sg13g2_buf_2
Xfanout1530 net1532 net1530 VPWR VGND sg13g2_buf_2
Xfanout1563 net1564 net1563 VPWR VGND sg13g2_buf_2
Xfanout1552 net1553 net1552 VPWR VGND sg13g2_buf_1
Xfanout1574 _3414_ net1574 VPWR VGND sg13g2_buf_8
XFILLER_20_1012 VPWR VGND sg13g2_decap_8
Xfanout1585 net1586 net1585 VPWR VGND sg13g2_buf_8
Xfanout1596 net1597 net1596 VPWR VGND sg13g2_buf_8
XFILLER_47_983 VPWR VGND sg13g2_decap_8
XFILLER_19_674 VPWR VGND sg13g2_fill_1
X_5860_ _1773_ s0.data_out\[13\]\[3\] net1409 VPWR VGND sg13g2_nand2b_1
XFILLER_34_622 VPWR VGND sg13g2_fill_2
X_4811_ _0168_ _0822_ _0823_ _3432_ net1593 VPWR VGND sg13g2_a22oi_1
XFILLER_15_891 VPWR VGND sg13g2_fill_2
X_5791_ net1626 _1633_ _1714_ VPWR VGND sg13g2_nor2_1
X_7530_ _3266_ VPWR _3280_ VGND _3275_ _3277_ sg13g2_o21ai_1
X_4742_ _0761_ net1493 _0762_ _0763_ VPWR VGND sg13g2_a21o_1
X_7461_ net1720 VPWR _3214_ VGND net715 _3209_ sg13g2_o21ai_1
X_4673_ _0153_ _0699_ _0700_ _3428_ net1589 VPWR VGND sg13g2_a22oi_1
X_6412_ net1676 _2269_ _2270_ VPWR VGND sg13g2_nor2_1
X_7392_ VGND VPWR _3154_ _3150_ net1648 sg13g2_or2_1
X_6343_ VGND VPWR net1637 _3403_ _0320_ _2203_ sg13g2_a21oi_1
X_6274_ VGND VPWR net1368 _2148_ _2151_ _2150_ sg13g2_a21oi_1
X_5225_ VPWR VGND _1197_ net1712 _1195_ net1708 _1198_ _1191_ sg13g2_a221oi_1
X_5156_ _1061_ _1139_ _1140_ _1141_ VPWR VGND sg13g2_nor3_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
X_4107_ VPWR _3483_ net582 VGND sg13g2_inv_1
X_5087_ _1072_ s0.data_out\[19\]\[2\] net1479 VPWR VGND sg13g2_nand2b_1
XFILLER_44_419 VPWR VGND sg13g2_fill_1
XFILLER_38_972 VPWR VGND sg13g2_decap_8
X_7688__338 VPWR VGND net338 sg13g2_tiehi
X_4038_ VPWR _3414_ net1695 VGND sg13g2_inv_1
XFILLER_13_828 VPWR VGND sg13g2_decap_8
X_5989_ VGND VPWR _1890_ _1864_ net1574 sg13g2_or2_1
XFILLER_8_309 VPWR VGND sg13g2_fill_2
X_7728_ net294 VGND VPWR _0206_ s0.valid_out\[19\][0] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_7659_ net25 VGND VPWR net638 s0.data_out\[25\]\[0\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_7740__281 VPWR VGND net281 sg13g2_tiehi
XFILLER_43_1012 VPWR VGND sg13g2_decap_8
XFILLER_0_754 VPWR VGND sg13g2_decap_8
XFILLER_48_725 VPWR VGND sg13g2_decap_8
XFILLER_15_110 VPWR VGND sg13g2_fill_2
XFILLER_44_953 VPWR VGND sg13g2_decap_8
XFILLER_7_34 VPWR VGND sg13g2_fill_1
Xhold309 s0.data_out\[18\]\[2\] VPWR VGND net678 sg13g2_dlygate4sd3_1
X_7647__38 VPWR VGND net38 sg13g2_tiehi
X_5010_ VGND VPWR net1484 _1005_ _1008_ _1007_ sg13g2_a21oi_1
Xfanout1393 net1396 net1393 VPWR VGND sg13g2_buf_2
Xfanout1382 net1384 net1382 VPWR VGND sg13g2_buf_8
Xfanout1371 s0.shift_out\[11\][0] net1371 VPWR VGND sg13g2_buf_8
Xfanout1360 net1364 net1360 VPWR VGND sg13g2_buf_8
XFILLER_47_780 VPWR VGND sg13g2_decap_8
X_6961_ net1639 net1255 _2762_ VPWR VGND sg13g2_nor2b_1
X_6892_ VGND VPWR net1274 _2699_ _2702_ _2701_ sg13g2_a21oi_1
X_5912_ _1823_ VPWR _1824_ VGND net1747 net657 sg13g2_o21ai_1
XFILLER_22_603 VPWR VGND sg13g2_decap_4
X_5843_ net1390 net1355 _1756_ VPWR VGND sg13g2_nor2b_1
XFILLER_35_997 VPWR VGND sg13g2_decap_8
X_7513_ net1213 net1339 _3263_ VPWR VGND sg13g2_nor2b_1
X_5774_ VGND VPWR _1686_ _1688_ _1699_ net1675 sg13g2_a21oi_1
X_4725_ _0746_ net530 net1517 VPWR VGND sg13g2_nand2b_1
XFILLER_30_680 VPWR VGND sg13g2_fill_1
X_7444_ net1218 s0.data_out\[1\]\[6\] _3199_ VPWR VGND sg13g2_and2_1
X_4656_ _0687_ VPWR _0688_ VGND net1726 net626 sg13g2_o21ai_1
X_4587_ _0620_ net1517 net816 VPWR VGND sg13g2_nand2_1
X_7375_ _3137_ net1686 _3136_ VPWR VGND sg13g2_nand2_1
X_6326_ _2191_ VPWR _2194_ VGND net1323 _2193_ sg13g2_o21ai_1
X_7694__331 VPWR VGND net331 sg13g2_tiehi
X_6257_ VPWR _2134_ _2133_ VGND sg13g2_inv_1
X_6188_ net1371 s0.data_out\[11\]\[6\] _2070_ VPWR VGND sg13g2_and2_1
X_5208_ _1181_ s0.data_out\[18\]\[2\] net1467 VPWR VGND sg13g2_nand2b_1
X_5139_ VGND VPWR net1473 _1121_ _1124_ _1123_ sg13g2_a21oi_1
XFILLER_40_433 VPWR VGND sg13g2_fill_1
XFILLER_41_989 VPWR VGND sg13g2_decap_8
XFILLER_8_117 VPWR VGND sg13g2_fill_2
XFILLER_12_146 VPWR VGND sg13g2_fill_1
XFILLER_12_157 VPWR VGND sg13g2_fill_2
XFILLER_12_168 VPWR VGND sg13g2_fill_1
XFILLER_8_139 VPWR VGND sg13g2_fill_2
XFILLER_8_128 VPWR VGND sg13g2_fill_2
XFILLER_5_813 VPWR VGND sg13g2_fill_1
XFILLER_4_312 VPWR VGND sg13g2_fill_2
XFILLER_10_1011 VPWR VGND sg13g2_decap_8
XFILLER_5_879 VPWR VGND sg13g2_decap_8
XFILLER_4_389 VPWR VGND sg13g2_fill_2
XFILLER_48_599 VPWR VGND sg13g2_decap_8
XFILLER_35_238 VPWR VGND sg13g2_fill_1
XFILLER_17_997 VPWR VGND sg13g2_decap_8
XFILLER_31_433 VPWR VGND sg13g2_fill_1
XFILLER_32_989 VPWR VGND sg13g2_decap_8
XFILLER_8_651 VPWR VGND sg13g2_fill_2
X_4510_ _0555_ net1184 _0554_ VPWR VGND sg13g2_nand2_1
X_5490_ VGND VPWR _1325_ _1438_ _1439_ net1440 sg13g2_a21oi_1
X_4441_ _0487_ VPWR _0489_ VGND s0.was_valid_out\[24\][0] net1528 sg13g2_o21ai_1
XFILLER_7_161 VPWR VGND sg13g2_fill_2
Xhold106 s0.shift_out\[18\][0] VPWR VGND net475 sg13g2_dlygate4sd3_1
Xhold117 _0338_ VPWR VGND net486 sg13g2_dlygate4sd3_1
Xhold139 _0096_ VPWR VGND net508 sg13g2_dlygate4sd3_1
Xhold128 s0.data_out\[20\]\[1\] VPWR VGND net497 sg13g2_dlygate4sd3_1
X_7160_ VGND VPWR _2946_ _2936_ net1649 sg13g2_or2_1
X_4372_ VGND VPWR _3600_ _0428_ _0429_ net1550 sg13g2_a21oi_1
X_6111_ _1998_ s0.shift_out\[11\][0] _1999_ _2000_ VPWR VGND sg13g2_a21o_1
X_7091_ net1715 net381 _0050_ VPWR VGND sg13g2_and2_1
XFILLER_39_500 VPWR VGND sg13g2_decap_8
X_6042_ _1940_ VPWR _1941_ VGND net1192 _1939_ sg13g2_o21ai_1
Xfanout1190 net1191 net1190 VPWR VGND sg13g2_buf_8
X_6944_ _2748_ VPWR _2749_ VGND net1174 _2747_ sg13g2_o21ai_1
XFILLER_35_761 VPWR VGND sg13g2_fill_1
X_6875_ net1704 _2660_ _2685_ VPWR VGND sg13g2_nor2_1
X_5826_ net1394 _1737_ _1742_ VPWR VGND sg13g2_nor2_1
X_5757_ _1682_ net1411 net726 VPWR VGND sg13g2_nand2_1
X_4708_ VGND VPWR net1495 _0728_ _0729_ _0727_ sg13g2_a21oi_1
X_7427_ VGND VPWR net1188 _3109_ _3186_ net1583 sg13g2_a21oi_1
X_5688_ net1428 VPWR _1617_ VGND _1552_ _1616_ sg13g2_o21ai_1
X_4639_ VGND VPWR _0549_ _0671_ _0672_ net1524 sg13g2_a21oi_1
XFILLER_2_805 VPWR VGND sg13g2_decap_8
X_7358_ s0.data_out\[2\]\[0\] s0.data_out\[1\]\[0\] net1224 _3120_ VPWR VGND sg13g2_mux2_1
X_6309_ _0310_ _2178_ _2179_ _3496_ net1612 VPWR VGND sg13g2_a22oi_1
X_7289_ _3051_ _3059_ _3023_ _3063_ VPWR VGND _3062_ sg13g2_nand4_1
XFILLER_40_1004 VPWR VGND sg13g2_decap_8
X_7634__52 VPWR VGND net52 sg13g2_tiehi
XFILLER_41_742 VPWR VGND sg13g2_fill_1
XFILLER_49_864 VPWR VGND sg13g2_decap_8
XFILLER_1_1020 VPWR VGND sg13g2_decap_8
X_4990_ _0988_ s0.data_out\[20\]\[7\] net1489 VPWR VGND sg13g2_nand2b_1
X_6660_ _2494_ s0.data_out\[7\]\[5\] net1303 VPWR VGND sg13g2_nand2b_1
X_6591_ _2427_ VPWR _2428_ VGND net1297 _2309_ sg13g2_o21ai_1
XFILLER_20_937 VPWR VGND sg13g2_fill_2
X_5611_ VGND VPWR net1425 _1545_ _1548_ _1547_ sg13g2_a21oi_1
XFILLER_32_786 VPWR VGND sg13g2_fill_2
X_5542_ _1487_ VPWR _1488_ VGND net1207 _1486_ sg13g2_o21ai_1
X_5473_ net1706 _1405_ _1422_ VPWR VGND sg13g2_nor2_1
X_4424_ net1533 s0.data_out\[25\]\[5\] _0475_ VPWR VGND sg13g2_and2_1
X_7212_ net1190 VPWR _2989_ VGND s0.was_valid_out\[2\][0] net1247 sg13g2_o21ai_1
X_4355_ _0412_ net501 net1557 VPWR VGND sg13g2_nand2b_1
X_7143_ _2919_ _2928_ _2918_ _2929_ VPWR VGND sg13g2_nand3_1
X_7074_ _0046_ _2863_ _2864_ _3525_ net1591 VPWR VGND sg13g2_a22oi_1
X_4286_ _0113_ _0352_ _0353_ _3419_ net1578 VPWR VGND sg13g2_a22oi_1
X_7869__142 VPWR VGND net142 sg13g2_tiehi
X_6025_ VGND VPWR _1926_ _1917_ net1665 sg13g2_or2_1
XFILLER_39_396 VPWR VGND sg13g2_fill_1
X_6927_ _2735_ VPWR _2736_ VGND net1730 net643 sg13g2_o21ai_1
XFILLER_35_580 VPWR VGND sg13g2_fill_2
X_6858_ _2668_ net1266 net580 VPWR VGND sg13g2_nand2_1
X_5809_ _1727_ VPWR _1728_ VGND net1196 _1726_ sg13g2_o21ai_1
X_6789_ _2609_ _2610_ _2611_ VPWR VGND sg13g2_nor2_1
X_7876__135 VPWR VGND net135 sg13g2_tiehi
XFILLER_2_646 VPWR VGND sg13g2_fill_1
XFILLER_1_189 VPWR VGND sg13g2_fill_1
XFILLER_38_52 VPWR VGND sg13g2_fill_2
XFILLER_46_834 VPWR VGND sg13g2_decap_8
XFILLER_6_952 VPWR VGND sg13g2_decap_8
X_4140_ VPWR _3516_ net554 VGND sg13g2_inv_1
XFILLER_49_661 VPWR VGND sg13g2_decap_8
X_4071_ _3447_ net563 VPWR VGND sg13g2_inv_2
X_7830_ net184 VGND VPWR net761 s0.data_out\[11\]\[3\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_7761_ net259 VGND VPWR _0239_ s0.data_out\[17\]\[6\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_4973_ _0970_ VPWR _0971_ VGND net1179 _0968_ sg13g2_o21ai_1
X_6712_ net471 _2536_ _2537_ VPWR VGND sg13g2_nor2_1
X_7692_ net333 VGND VPWR _0170_ s0.valid_out\[22\][0] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_6643_ _2475_ net1287 _2476_ _2477_ VPWR VGND sg13g2_a21o_1
XFILLER_32_561 VPWR VGND sg13g2_fill_1
Xclkload9 clknet_leaf_26_clk clkload9/X VPWR VGND sg13g2_buf_8
X_6574_ _3394_ _3509_ _2414_ VPWR VGND sg13g2_nor2_1
XFILLER_30_1014 VPWR VGND sg13g2_decap_8
X_5525_ _1473_ VPWR _1474_ VGND _1431_ _1433_ sg13g2_o21ai_1
X_5456_ VGND VPWR net1437 _1402_ _1405_ _1404_ sg13g2_a21oi_1
X_4407_ VPWR _0125_ _0462_ VGND sg13g2_inv_1
X_5387_ VGND VPWR _1227_ _1347_ _1348_ net1450 sg13g2_a21oi_1
X_4338_ net1535 net1352 _0395_ VPWR VGND sg13g2_nor2b_1
X_7126_ VGND VPWR net1242 _2910_ _2912_ _2911_ sg13g2_a21oi_1
X_4269_ VGND VPWR net1559 _3632_ _3633_ _3628_ sg13g2_a21oi_1
X_7057_ net1591 _2775_ _2852_ VPWR VGND sg13g2_nor2_1
XFILLER_28_834 VPWR VGND sg13g2_fill_2
X_6008_ _1908_ VPWR _1909_ VGND net1693 _1888_ sg13g2_o21ai_1
XFILLER_28_867 VPWR VGND sg13g2_fill_1
X_7959_ net256 VGND VPWR _0093_ s0.data_out\[1\]\[5\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_42_314 VPWR VGND sg13g2_fill_1
XFILLER_11_701 VPWR VGND sg13g2_fill_2
XFILLER_11_767 VPWR VGND sg13g2_fill_1
XFILLER_24_87 VPWR VGND sg13g2_fill_1
XFILLER_40_75 VPWR VGND sg13g2_fill_1
XFILLER_3_900 VPWR VGND sg13g2_decap_8
XFILLER_3_977 VPWR VGND sg13g2_decap_8
Xfanout1723 net1724 net1723 VPWR VGND sg13g2_buf_8
Xfanout1701 net1704 net1701 VPWR VGND sg13g2_buf_8
Xfanout1712 net1713 net1712 VPWR VGND sg13g2_buf_8
Xfanout1745 net1746 net1745 VPWR VGND sg13g2_buf_1
Xfanout1734 net1737 net1734 VPWR VGND sg13g2_buf_8
XFILLER_1_69 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_18 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_34_837 VPWR VGND sg13g2_fill_2
XFILLER_21_509 VPWR VGND sg13g2_fill_1
XFILLER_14_1009 VPWR VGND sg13g2_decap_8
X_5310_ net1462 VPWR _1275_ VGND _1218_ _1274_ sg13g2_o21ai_1
X_6290_ net1321 net589 _2165_ VPWR VGND sg13g2_and2_1
X_5241_ VGND VPWR _1100_ _1213_ _1214_ net1461 sg13g2_a21oi_1
XFILLER_5_292 VPWR VGND sg13g2_fill_2
X_5172_ net1198 _3454_ _1153_ VPWR VGND sg13g2_nor2_1
X_4123_ VPWR _3499_ net443 VGND sg13g2_inv_1
X_4054_ VPWR _3430_ net601 VGND sg13g2_inv_1
X_7813_ net202 VGND VPWR _0291_ s0.genblk1\[11\].modules.bubble clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
XFILLER_36_174 VPWR VGND sg13g2_fill_1
X_7744_ net277 VGND VPWR _0222_ s0.data_out\[18\]\[1\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_4956_ _0834_ VPWR _0954_ VGND net1492 _3449_ sg13g2_o21ai_1
XFILLER_33_870 VPWR VGND sg13g2_fill_1
X_7727__296 VPWR VGND net296 sg13g2_tiehi
X_7675_ net352 VGND VPWR net699 s0.data_out\[24\]\[4\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_4887_ s0.data_out\[22\]\[4\] s0.data_out\[21\]\[4\] net1491 _0896_ VPWR VGND sg13g2_mux2_1
X_6626_ s0.data_out\[8\]\[3\] s0.data_out\[7\]\[3\] net1290 _2460_ VPWR VGND sg13g2_mux2_1
X_6557_ _3394_ _3513_ _2401_ VPWR VGND sg13g2_nor2_1
X_5508_ _1457_ net1442 _1456_ VPWR VGND sg13g2_nand2b_1
X_6488_ s0.data_out\[9\]\[0\] s0.data_out\[8\]\[0\] net1302 _2334_ VPWR VGND sg13g2_mux2_1
X_7873__138 VPWR VGND net138 sg13g2_tiehi
X_5439_ _1389_ _1390_ _1391_ VPWR VGND sg13g2_nor2_1
XFILLER_0_936 VPWR VGND sg13g2_decap_8
XFILLER_48_907 VPWR VGND sg13g2_decap_8
X_7109_ _2895_ net1170 _2894_ VPWR VGND sg13g2_nand2_1
XFILLER_28_642 VPWR VGND sg13g2_fill_1
XFILLER_11_542 VPWR VGND sg13g2_decap_4
XFILLER_7_524 VPWR VGND sg13g2_fill_2
XFILLER_7_502 VPWR VGND sg13g2_decap_8
X_7659__25 VPWR VGND net25 sg13g2_tiehi
XFILLER_3_763 VPWR VGND sg13g2_decap_8
Xfanout1542 net1543 net1542 VPWR VGND sg13g2_buf_8
Xfanout1520 net1527 net1520 VPWR VGND sg13g2_buf_1
Xfanout1531 net1532 net1531 VPWR VGND sg13g2_buf_1
Xfanout1575 net1576 net1575 VPWR VGND sg13g2_buf_8
Xfanout1553 net826 net1553 VPWR VGND sg13g2_buf_2
Xfanout1564 s0.valid_out\[27\][0] net1564 VPWR VGND sg13g2_buf_8
XFILLER_38_439 VPWR VGND sg13g2_fill_2
Xfanout1586 net1587 net1586 VPWR VGND sg13g2_buf_8
XFILLER_19_642 VPWR VGND sg13g2_decap_8
Xfanout1597 net1602 net1597 VPWR VGND sg13g2_buf_8
XFILLER_47_962 VPWR VGND sg13g2_decap_8
XFILLER_33_111 VPWR VGND sg13g2_fill_1
X_4810_ net1593 _0758_ _0823_ VPWR VGND sg13g2_nor2_1
X_5790_ net1414 VPWR _1713_ VGND _1630_ _1712_ sg13g2_o21ai_1
X_4741_ net1493 net1334 _0762_ VPWR VGND sg13g2_nor2b_1
X_7460_ VGND VPWR _3207_ _3210_ _3213_ _3212_ sg13g2_a21oi_1
X_4672_ net1589 _0666_ _0700_ VPWR VGND sg13g2_nor2_1
X_6411_ VGND VPWR net1324 _2266_ _2269_ _2268_ sg13g2_a21oi_1
X_7391_ net1648 _3150_ _3153_ VPWR VGND sg13g2_nor2_1
X_6342_ net1637 net1338 _2203_ VPWR VGND sg13g2_nor2_1
X_6273_ VGND VPWR _2024_ _2149_ _2150_ net1368 sg13g2_a21oi_1
X_5224_ _1197_ net1198 _1196_ VPWR VGND sg13g2_nand2_1
XFILLER_5_1007 VPWR VGND sg13g2_decap_8
X_5155_ _1114_ _1116_ _1140_ VPWR VGND sg13g2_nor2b_1
X_4106_ VPWR _3482_ net575 VGND sg13g2_inv_1
XFILLER_38_951 VPWR VGND sg13g2_decap_8
X_5086_ _1069_ net1458 _1070_ _1071_ VPWR VGND sg13g2_a21o_1
X_4037_ VPWR _3413_ net632 VGND sg13g2_inv_1
XFILLER_40_615 VPWR VGND sg13g2_fill_2
X_5988_ _1889_ net1694 _1888_ VPWR VGND sg13g2_nand2_1
X_7727_ net296 VGND VPWR net438 s0.was_valid_out\[19\][0] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_4939_ _0180_ _0938_ _0939_ _3437_ net1605 VPWR VGND sg13g2_a22oi_1
X_7658_ net26 VGND VPWR _0136_ s0.shift_out\[25\][0] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_21_873 VPWR VGND sg13g2_fill_1
X_6609_ _2443_ net1289 net802 VPWR VGND sg13g2_nand2_1
X_7589_ net1669 _3326_ _3327_ VPWR VGND sg13g2_nor2_1
X_7656__28 VPWR VGND net28 sg13g2_tiehi
XFILLER_0_733 VPWR VGND sg13g2_decap_8
XFILLER_48_704 VPWR VGND sg13g2_decap_8
XFILLER_44_932 VPWR VGND sg13g2_decap_8
X_7962__217 VPWR VGND net217 sg13g2_tiehi
XFILLER_28_483 VPWR VGND sg13g2_fill_2
XFILLER_31_615 VPWR VGND sg13g2_fill_1
XFILLER_12_862 VPWR VGND sg13g2_fill_1
Xfanout1350 net1351 net1350 VPWR VGND sg13g2_buf_8
Xfanout1383 net1384 net1383 VPWR VGND sg13g2_buf_1
Xfanout1361 net1364 net1361 VPWR VGND sg13g2_buf_1
Xfanout1372 net1373 net1372 VPWR VGND sg13g2_buf_8
Xfanout1394 net1396 net1394 VPWR VGND sg13g2_buf_8
X_6960_ net1258 VPWR _2761_ VGND net1641 net1251 sg13g2_o21ai_1
X_5911_ _1822_ VPWR _1823_ VGND net1195 _1821_ sg13g2_o21ai_1
XFILLER_35_932 VPWR VGND sg13g2_fill_1
X_6891_ VGND VPWR _2575_ _2700_ _2701_ net1274 sg13g2_a21oi_1
XFILLER_35_976 VPWR VGND sg13g2_decap_8
X_5842_ _1754_ VPWR _1755_ VGND net1397 _3481_ sg13g2_o21ai_1
X_5773_ _1698_ _1689_ _1697_ VPWR VGND sg13g2_nand2_1
X_7512_ s0.data_out\[1\]\[5\] s0.data_out\[0\]\[5\] net1215 _3262_ VPWR VGND sg13g2_mux2_1
X_4724_ _0743_ net1496 _0744_ _0745_ VPWR VGND sg13g2_a21o_1
X_7443_ VPWR _0081_ net596 VGND sg13g2_inv_1
X_7724__299 VPWR VGND net299 sg13g2_tiehi
X_4655_ _0632_ _0686_ net1725 _0687_ VPWR VGND sg13g2_nand3_1
X_7374_ VGND VPWR net1232 _3133_ _3136_ _3135_ sg13g2_a21oi_1
X_4586_ net1696 _0618_ _0619_ VPWR VGND sg13g2_nor2_1
X_6325_ s0.was_valid_out\[9\][0] net1362 _2193_ VPWR VGND sg13g2_nor2_1
X_6256_ _2133_ _2132_ net1653 _2125_ net1663 VPWR VGND sg13g2_a22oi_1
X_6187_ _0298_ _2068_ _2069_ _3488_ net1612 VPWR VGND sg13g2_a22oi_1
X_5207_ _1178_ net1447 _1179_ _1180_ VPWR VGND sg13g2_a21o_1
X_5138_ VGND VPWR _1010_ _1122_ _1123_ net1473 sg13g2_a21oi_1
XFILLER_45_707 VPWR VGND sg13g2_fill_1
XFILLER_45_729 VPWR VGND sg13g2_decap_8
X_5069_ net1736 net387 _0192_ VPWR VGND sg13g2_and2_1
XFILLER_16_11 VPWR VGND sg13g2_fill_1
XFILLER_26_998 VPWR VGND sg13g2_decap_8
XFILLER_41_968 VPWR VGND sg13g2_decap_8
XFILLER_13_659 VPWR VGND sg13g2_fill_1
XFILLER_32_87 VPWR VGND sg13g2_fill_2
XFILLER_0_563 VPWR VGND sg13g2_fill_1
XFILLER_48_578 VPWR VGND sg13g2_decap_8
XFILLER_44_751 VPWR VGND sg13g2_decap_8
XFILLER_17_976 VPWR VGND sg13g2_decap_8
XFILLER_32_968 VPWR VGND sg13g2_decap_8
XFILLER_40_990 VPWR VGND sg13g2_decap_8
X_4440_ VGND VPWR net1184 _0376_ _0488_ _0487_ sg13g2_a21oi_1
Xhold107 _1279_ VPWR VGND net476 sg13g2_dlygate4sd3_1
X_7678__349 VPWR VGND net349 sg13g2_tiehi
Xhold118 s0.data_out\[18\]\[3\] VPWR VGND net487 sg13g2_dlygate4sd3_1
Xhold129 _0198_ VPWR VGND net498 sg13g2_dlygate4sd3_1
X_4371_ _0428_ net556 net1556 VPWR VGND sg13g2_nand2b_1
X_6110_ net1367 net1169 _1999_ VPWR VGND sg13g2_nor2_1
X_7090_ net1580 _2870_ _2871_ _0049_ VPWR VGND sg13g2_nor3_1
X_6041_ VGND VPWR net1192 _1870_ _1940_ net1627 sg13g2_a21oi_1
Xfanout1180 _3391_ net1180 VPWR VGND sg13g2_buf_8
Xfanout1191 _3384_ net1191 VPWR VGND sg13g2_buf_8
XFILLER_27_718 VPWR VGND sg13g2_fill_2
X_6943_ VGND VPWR net1174 _2720_ _2748_ net1602 sg13g2_a21oi_1
X_7730__292 VPWR VGND net292 sg13g2_tiehi
X_6874_ net1688 _2683_ _2684_ VPWR VGND sg13g2_nor2_1
XFILLER_22_434 VPWR VGND sg13g2_fill_2
X_5825_ _1738_ VPWR _1741_ VGND net416 net1399 sg13g2_o21ai_1
X_5756_ _1679_ _1677_ _1681_ VPWR VGND _1678_ sg13g2_nand3b_1
XFILLER_33_1023 VPWR VGND sg13g2_decap_4
X_4707_ s0.data_out\[23\]\[0\] s0.data_out\[22\]\[0\] net1504 _0728_ VPWR VGND sg13g2_mux2_1
X_5687_ net1196 _3472_ _1616_ VPWR VGND sg13g2_nor2_1
X_7426_ VGND VPWR net1222 net659 _3185_ _3107_ sg13g2_a21oi_1
X_4638_ _0671_ s0.data_out\[23\]\[5\] net1530 VPWR VGND sg13g2_nand2b_1
X_4569_ _0605_ _0604_ _0603_ VPWR VGND sg13g2_nand2b_1
X_7357_ _3116_ _3118_ net1702 _3119_ VPWR VGND sg13g2_nand3_1
X_6308_ net1612 _2150_ _2179_ VPWR VGND sg13g2_nor2_1
X_7288_ _3049_ _3060_ _3061_ _3062_ VPWR VGND sg13g2_nor3_1
X_6239_ VGND VPWR net1366 _2113_ _2116_ _2115_ sg13g2_a21oi_1
XFILLER_27_98 VPWR VGND sg13g2_fill_1
XFILLER_49_843 VPWR VGND sg13g2_decap_8
XFILLER_1_894 VPWR VGND sg13g2_decap_8
X_7684__342 VPWR VGND net342 sg13g2_tiehi
XFILLER_17_784 VPWR VGND sg13g2_fill_1
XFILLER_17_1018 VPWR VGND sg13g2_decap_8
X_6590_ VGND VPWR _2427_ _2426_ _2425_ sg13g2_or2_1
X_5610_ VGND VPWR _1423_ _1546_ _1547_ net1425 sg13g2_a21oi_1
XFILLER_31_275 VPWR VGND sg13g2_fill_2
X_5541_ VGND VPWR net1206 _1417_ _1487_ net1620 sg13g2_a21oi_1
XFILLER_8_471 VPWR VGND sg13g2_fill_2
X_5472_ _1421_ net1573 _1419_ VPWR VGND sg13g2_xnor2_1
X_7211_ net1229 _2983_ _2988_ VPWR VGND sg13g2_nor2_1
X_4423_ _0129_ _0473_ _0474_ _3407_ net1579 VPWR VGND sg13g2_a22oi_1
X_4354_ _0409_ net1535 _0410_ _0411_ VPWR VGND sg13g2_a21o_1
X_7142_ _2928_ net1677 _2926_ VPWR VGND sg13g2_xnor2_1
X_7691__335 VPWR VGND net335 sg13g2_tiehi
X_7073_ net1591 _2814_ _2864_ VPWR VGND sg13g2_nor2_1
X_6024_ _1925_ _1924_ net1655 _1917_ net1665 VPWR VGND sg13g2_a22oi_1
X_4285_ net1578 _3579_ _0353_ VPWR VGND sg13g2_nor2_1
XFILLER_27_515 VPWR VGND sg13g2_decap_4
X_7631__56 VPWR VGND net56 sg13g2_tiehi
X_6926_ _2662_ _2734_ net1730 _2735_ VPWR VGND sg13g2_nand3_1
X_6857_ VPWR VGND _2666_ net1713 _2662_ net1703 _2667_ _2660_ sg13g2_a221oi_1
X_6788_ VGND VPWR _2605_ _2607_ _2610_ net1670 sg13g2_a21oi_1
XFILLER_13_23 VPWR VGND sg13g2_fill_1
XFILLER_22_264 VPWR VGND sg13g2_fill_1
X_5808_ VGND VPWR _3380_ _1687_ _1727_ net1630 sg13g2_a21oi_1
X_5739_ s0.data_out\[15\]\[7\] s0.data_out\[14\]\[7\] net1410 _1664_ VPWR VGND sg13g2_mux2_1
X_7409_ _3170_ VPWR _3171_ VGND _3403_ _3160_ sg13g2_o21ai_1
Xhold460 s0.data_new_delayed\[4\] VPWR VGND net829 sg13g2_dlygate4sd3_1
XFILLER_46_802 VPWR VGND sg13g2_fill_1
XFILLER_46_813 VPWR VGND sg13g2_decap_8
X_7668__359 VPWR VGND net359 sg13g2_tiehi
XFILLER_6_931 VPWR VGND sg13g2_decap_8
XFILLER_6_920 VPWR VGND sg13g2_decap_8
XFILLER_9_279 VPWR VGND sg13g2_fill_2
XFILLER_49_640 VPWR VGND sg13g2_decap_8
X_4070_ VPWR _3446_ net509 VGND sg13g2_inv_1
XFILLER_37_868 VPWR VGND sg13g2_fill_1
XFILLER_36_323 VPWR VGND sg13g2_fill_2
XFILLER_24_518 VPWR VGND sg13g2_fill_1
X_7760_ net260 VGND VPWR _0238_ s0.data_out\[17\]\[5\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_4972_ _0970_ net1179 _0969_ VPWR VGND sg13g2_nand2_1
XFILLER_24_529 VPWR VGND sg13g2_fill_2
X_6711_ _2535_ VPWR _2536_ VGND net1285 _2426_ sg13g2_o21ai_1
X_7691_ net335 VGND VPWR _0169_ s0.was_valid_out\[22\][0] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_6642_ net1286 net1332 _2476_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_724 VPWR VGND sg13g2_fill_2
X_6573_ VPWR _0340_ _2413_ VGND sg13g2_inv_1
X_5524_ _1452_ _1469_ _1470_ _1472_ _1473_ VPWR VGND sg13g2_nor4_1
X_5455_ VGND VPWR _1292_ _1403_ _1404_ net1436 sg13g2_a21oi_1
X_4406_ _0461_ VPWR _0462_ VGND net1715 net798 sg13g2_o21ai_1
X_5386_ _1347_ s0.data_out\[17\]\[5\] net1455 VPWR VGND sg13g2_nand2b_1
X_7125_ net1242 net1338 _2911_ VPWR VGND sg13g2_nor2b_1
X_4337_ _0393_ VPWR _0394_ VGND net1540 _3416_ sg13g2_o21ai_1
X_4268_ _3630_ net1545 _3631_ _3632_ VPWR VGND sg13g2_a21o_1
X_7056_ net1260 VPWR _2851_ VGND _2772_ _2850_ sg13g2_o21ai_1
X_6007_ _1908_ net1675 _1906_ VPWR VGND sg13g2_nand2_1
X_4199_ VGND VPWR net1564 _3413_ _3563_ _3562_ sg13g2_a21oi_1
X_7958_ net269 VGND VPWR _0092_ s0.data_out\[1\]\[4\] clknet_leaf_12_clk sg13g2_dfrbpq_2
X_7889_ net121 VGND VPWR _0023_ s0.data_out\[7\]\[7\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_6909_ _2719_ net1275 _2718_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_562 VPWR VGND sg13g2_decap_8
XFILLER_11_735 VPWR VGND sg13g2_decap_4
XFILLER_6_227 VPWR VGND sg13g2_fill_1
XFILLER_3_956 VPWR VGND sg13g2_decap_8
Xhold290 s0.data_out\[1\]\[2\] VPWR VGND net659 sg13g2_dlygate4sd3_1
Xfanout1724 net1733 net1724 VPWR VGND sg13g2_buf_8
Xfanout1713 ui_in[0] net1713 VPWR VGND sg13g2_buf_8
Xfanout1702 net1704 net1702 VPWR VGND sg13g2_buf_1
Xfanout1746 net1750 net1746 VPWR VGND sg13g2_buf_8
Xfanout1735 net1737 net1735 VPWR VGND sg13g2_buf_1
XFILLER_46_610 VPWR VGND sg13g2_fill_1
Xheichips25_top_sorter_19 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_46_676 VPWR VGND sg13g2_fill_1
X_7681__345 VPWR VGND net345 sg13g2_tiehi
X_7859__153 VPWR VGND net153 sg13g2_tiehi
X_5240_ _1213_ s0.data_out\[18\]\[6\] net1466 VPWR VGND sg13g2_nand2b_1
X_5171_ _0199_ _1151_ _1152_ _3449_ net1607 VPWR VGND sg13g2_a22oi_1
X_4122_ VPWR _3498_ net589 VGND sg13g2_inv_1
X_4053_ VPWR _3429_ net478 VGND sg13g2_inv_1
X_7866__146 VPWR VGND net146 sg13g2_tiehi
X_7812_ net203 VGND VPWR _0290_ s0.valid_out\[12\][0] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_4955_ VGND VPWR net1470 _0951_ _0953_ _0952_ sg13g2_a21oi_1
X_7743_ net278 VGND VPWR _0221_ s0.data_out\[18\]\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_4886_ _0895_ net1489 s0.data_out\[21\]\[4\] VPWR VGND sg13g2_nand2_1
X_7674_ net353 VGND VPWR net479 s0.data_out\[24\]\[3\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_6625_ _2459_ net1290 net593 VPWR VGND sg13g2_nand2_1
X_6556_ VPWR _0336_ _2400_ VGND sg13g2_inv_1
XFILLER_4_709 VPWR VGND sg13g2_fill_1
X_5507_ VGND VPWR net1426 _1454_ _1456_ _1455_ sg13g2_a21oi_1
X_6487_ VGND VPWR net1305 _2330_ _2333_ _2332_ sg13g2_a21oi_1
X_5438_ net1644 _3376_ _1390_ VPWR VGND sg13g2_nor2_1
X_5369_ VGND VPWR _1216_ _1329_ _1330_ net1451 sg13g2_a21oi_1
XFILLER_0_915 VPWR VGND sg13g2_decap_8
X_7108_ s0.data_out\[3\]\[0\] s0.data_out\[4\]\[0\] net1253 _2894_ VPWR VGND sg13g2_mux2_1
X_7039_ _2819_ _2834_ _2835_ _2836_ _2837_ VPWR VGND sg13g2_nor4_1
XFILLER_28_621 VPWR VGND sg13g2_fill_1
XFILLER_43_602 VPWR VGND sg13g2_fill_1
XFILLER_24_860 VPWR VGND sg13g2_fill_2
XFILLER_2_296 VPWR VGND sg13g2_fill_1
Xfanout1532 s0.valid_out\[24\][0] net1532 VPWR VGND sg13g2_buf_1
Xfanout1521 net1522 net1521 VPWR VGND sg13g2_buf_2
Xfanout1510 net1511 net1510 VPWR VGND sg13g2_buf_2
Xfanout1554 s0.valid_out\[26\][0] net1554 VPWR VGND sg13g2_buf_8
Xfanout1543 s0.valid_out\[25\][0] net1543 VPWR VGND sg13g2_buf_8
Xfanout1565 net1569 net1565 VPWR VGND sg13g2_buf_8
XFILLER_47_941 VPWR VGND sg13g2_decap_8
Xfanout1587 net1588 net1587 VPWR VGND sg13g2_buf_8
Xfanout1576 net1577 net1576 VPWR VGND sg13g2_buf_8
Xfanout1598 net1602 net1598 VPWR VGND sg13g2_buf_8
XFILLER_33_101 VPWR VGND sg13g2_fill_2
XFILLER_33_123 VPWR VGND sg13g2_fill_2
XFILLER_22_819 VPWR VGND sg13g2_decap_4
X_4740_ s0.data_out\[23\]\[6\] s0.data_out\[22\]\[6\] net1503 _0761_ VPWR VGND sg13g2_mux2_1
XFILLER_15_893 VPWR VGND sg13g2_fill_1
XFILLER_30_841 VPWR VGND sg13g2_fill_1
X_4671_ net1524 VPWR _0699_ VGND _0663_ _0698_ sg13g2_o21ai_1
X_6410_ VGND VPWR _2145_ _2267_ _2268_ net1324 sg13g2_a21oi_1
XFILLER_30_885 VPWR VGND sg13g2_fill_2
XFILLER_30_896 VPWR VGND sg13g2_fill_1
X_7390_ net1659 _3144_ _3152_ VPWR VGND sg13g2_nor2_1
X_6341_ VGND VPWR net1637 _3406_ _0319_ _2202_ sg13g2_a21oi_1
XFILLER_6_580 VPWR VGND sg13g2_decap_4
X_6272_ _2149_ net493 net1374 VPWR VGND sg13g2_nand2b_1
XFILLER_6_591 VPWR VGND sg13g2_fill_1
X_5223_ s0.data_out\[18\]\[0\] s0.data_out\[19\]\[0\] net1465 _1196_ VPWR VGND sg13g2_mux2_1
X_5154_ VGND VPWR _1133_ _1138_ _1139_ _1117_ sg13g2_a21oi_1
X_4105_ VPWR _3481_ net603 VGND sg13g2_inv_1
X_5085_ net1458 net1350 _1070_ VPWR VGND sg13g2_nor2b_1
X_4036_ VPWR _3412_ net464 VGND sg13g2_inv_1
XFILLER_37_484 VPWR VGND sg13g2_fill_2
XFILLER_24_134 VPWR VGND sg13g2_fill_2
XFILLER_40_627 VPWR VGND sg13g2_fill_1
XFILLER_36_1021 VPWR VGND sg13g2_decap_8
X_5987_ VGND VPWR net1391 _1885_ _1888_ _1887_ sg13g2_a21oi_1
X_7726_ net297 VGND VPWR net628 s0.data_out\[20\]\[7\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_4938_ net1604 _0872_ _0939_ VPWR VGND sg13g2_nor2_1
X_4869_ _0878_ s0.data_out\[21\]\[6\] net1505 VPWR VGND sg13g2_nand2b_1
X_7657_ net27 VGND VPWR _0135_ s0.genblk1\[24\].modules.bubble clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_21_12 VPWR VGND sg13g2_decap_8
X_6608_ net1699 _2441_ _2442_ VPWR VGND sg13g2_nor2_1
X_7588_ _3325_ VPWR _3326_ VGND _3393_ net1338 sg13g2_o21ai_1
X_6539_ _2382_ _2384_ net1685 _2385_ VPWR VGND sg13g2_nand3_1
XFILLER_0_712 VPWR VGND sg13g2_decap_8
XFILLER_0_789 VPWR VGND sg13g2_decap_8
XFILLER_44_911 VPWR VGND sg13g2_decap_8
XFILLER_16_613 VPWR VGND sg13g2_fill_2
XFILLER_29_985 VPWR VGND sg13g2_decap_8
XFILLER_44_988 VPWR VGND sg13g2_decap_8
XFILLER_30_115 VPWR VGND sg13g2_fill_2
XFILLER_7_311 VPWR VGND sg13g2_fill_2
XFILLER_7_355 VPWR VGND sg13g2_decap_8
XFILLER_7_377 VPWR VGND sg13g2_decap_8
X_7856__156 VPWR VGND net156 sg13g2_tiehi
XFILLER_3_594 VPWR VGND sg13g2_decap_8
Xfanout1340 net1342 net1340 VPWR VGND sg13g2_buf_8
Xfanout1362 net1364 net1362 VPWR VGND sg13g2_buf_8
Xfanout1384 net1385 net1384 VPWR VGND sg13g2_buf_1
XFILLER_16_4 VPWR VGND sg13g2_fill_1
Xfanout1351 s0.data_new_delayed\[2\] net1351 VPWR VGND sg13g2_buf_8
Xfanout1373 s0.valid_out\[11\][0] net1373 VPWR VGND sg13g2_buf_8
Xfanout1395 net1396 net1395 VPWR VGND sg13g2_buf_1
X_5910_ VGND VPWR net1195 _1765_ _1822_ net1626 sg13g2_a21oi_1
X_6890_ _2700_ net566 net1280 VPWR VGND sg13g2_nand2b_1
XFILLER_35_944 VPWR VGND sg13g2_fill_2
XFILLER_35_955 VPWR VGND sg13g2_decap_8
X_7863__149 VPWR VGND net149 sg13g2_tiehi
X_5841_ _1754_ net1397 s0.data_out\[13\]\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_22_638 VPWR VGND sg13g2_fill_1
X_5772_ _1694_ _1696_ net1684 _1697_ VPWR VGND sg13g2_nand3_1
X_7511_ _3261_ net1201 _3260_ VPWR VGND sg13g2_nand2_1
X_4723_ net1496 net1169 _0744_ VPWR VGND sg13g2_nor2_1
X_7442_ _3197_ VPWR _3198_ VGND net1719 net595 sg13g2_o21ai_1
X_4654_ net1525 VPWR _0686_ VGND _0628_ _0685_ sg13g2_o21ai_1
X_7373_ VGND VPWR _3015_ _3134_ _3135_ net1232 sg13g2_a21oi_1
X_4585_ VGND VPWR net1525 _0615_ _0618_ _0617_ sg13g2_a21oi_1
X_6324_ net1311 _2187_ _2192_ VPWR VGND sg13g2_nor2_1
X_6255_ VGND VPWR net1368 _2129_ _2132_ _2131_ sg13g2_a21oi_1
X_5206_ net1448 net1350 _1179_ VPWR VGND sg13g2_nor2b_1
X_6186_ net1612 _2029_ _2069_ VPWR VGND sg13g2_nor2_1
X_5137_ _1122_ _3392_ net435 VPWR VGND sg13g2_nand2_1
X_5068_ _0191_ _1056_ _1057_ _3441_ net1604 VPWR VGND sg13g2_a22oi_1
X_4019_ VPWR _3395_ net1284 VGND sg13g2_inv_1
XFILLER_38_793 VPWR VGND sg13g2_fill_1
XFILLER_40_402 VPWR VGND sg13g2_fill_2
XFILLER_16_45 VPWR VGND sg13g2_fill_2
XFILLER_41_947 VPWR VGND sg13g2_decap_8
XFILLER_12_159 VPWR VGND sg13g2_fill_1
X_7709_ net315 VGND VPWR net535 s0.data_out\[21\]\[3\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_32_44 VPWR VGND sg13g2_fill_2
XFILLER_4_369 VPWR VGND sg13g2_fill_1
XFILLER_48_557 VPWR VGND sg13g2_decap_8
XFILLER_31_413 VPWR VGND sg13g2_fill_2
XFILLER_8_653 VPWR VGND sg13g2_fill_1
Xhold108 s0.shift_out\[21\][0] VPWR VGND net477 sg13g2_dlygate4sd3_1
X_4370_ _0425_ net1534 _0426_ _0427_ VPWR VGND sg13g2_a21o_1
Xhold119 _0224_ VPWR VGND net488 sg13g2_dlygate4sd3_1
XFILLER_4_892 VPWR VGND sg13g2_decap_8
X_6040_ VGND VPWR net1378 net513 _1939_ _1867_ sg13g2_a21oi_1
XFILLER_39_524 VPWR VGND sg13g2_fill_2
Xfanout1181 net1183 net1181 VPWR VGND sg13g2_buf_8
X_7643__43 VPWR VGND net43 sg13g2_tiehi
Xfanout1170 net1172 net1170 VPWR VGND sg13g2_buf_8
Xfanout1192 net1193 net1192 VPWR VGND sg13g2_buf_8
X_6942_ VGND VPWR net1265 s0.data_out\[5\]\[4\] _2747_ _2715_ sg13g2_a21oi_1
X_6873_ VGND VPWR net1273 _2680_ _2683_ _2682_ sg13g2_a21oi_1
X_5824_ _1739_ VPWR _1740_ VGND net1407 _1620_ sg13g2_o21ai_1
XFILLER_33_1002 VPWR VGND sg13g2_decap_8
X_5755_ VPWR _1680_ _1679_ VGND sg13g2_inv_1
X_4706_ net1495 net1359 _0727_ VPWR VGND sg13g2_nor2b_1
X_5686_ VPWR _0251_ net743 VGND sg13g2_inv_1
X_4637_ _0668_ net1508 _0669_ _0670_ VPWR VGND sg13g2_a21o_1
X_7425_ VPWR _0077_ net751 VGND sg13g2_inv_1
X_4568_ _0604_ net1634 net1516 VPWR VGND sg13g2_nand2_1
X_7356_ _3118_ net1187 _3117_ VPWR VGND sg13g2_nand2_1
X_6307_ net1368 VPWR _2178_ VGND _2147_ _2177_ sg13g2_o21ai_1
X_4499_ _0544_ _0543_ net1658 _0536_ net1647 VPWR VGND sg13g2_a22oi_1
X_7287_ net1678 _3058_ _3061_ VPWR VGND sg13g2_nor2_1
X_6238_ VGND VPWR _1997_ _2114_ _2115_ net1366 sg13g2_a21oi_1
X_6169_ net1614 _1987_ _2056_ VPWR VGND sg13g2_nor2_1
XFILLER_26_763 VPWR VGND sg13g2_fill_2
XFILLER_13_413 VPWR VGND sg13g2_fill_2
XFILLER_14_936 VPWR VGND sg13g2_fill_2
XFILLER_43_65 VPWR VGND sg13g2_fill_2
XFILLER_41_788 VPWR VGND sg13g2_fill_1
XFILLER_22_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_20_clk clknet_3_6__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_5_656 VPWR VGND sg13g2_fill_2
XFILLER_4_122 VPWR VGND sg13g2_fill_1
XFILLER_4_155 VPWR VGND sg13g2_decap_4
X_7677__350 VPWR VGND net350 sg13g2_tiehi
XFILLER_49_822 VPWR VGND sg13g2_decap_8
XFILLER_1_873 VPWR VGND sg13g2_decap_8
XFILLER_49_899 VPWR VGND sg13g2_decap_8
X_7640__46 VPWR VGND net46 sg13g2_tiehi
Xclkbuf_leaf_11_clk clknet_3_2__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
XFILLER_13_991 VPWR VGND sg13g2_decap_8
X_5540_ VGND VPWR net1423 net655 _1486_ _1415_ sg13g2_a21oi_1
XFILLER_9_995 VPWR VGND sg13g2_decap_8
X_5471_ VGND VPWR _1420_ _1419_ net1573 sg13g2_or2_1
X_4422_ net1579 _0441_ _0474_ VPWR VGND sg13g2_nor2_1
X_7210_ _2985_ VPWR _2987_ VGND s0.was_valid_out\[2\][0] net1235 sg13g2_o21ai_1
X_4353_ net1535 net1167 _0410_ VPWR VGND sg13g2_nor2_1
X_7141_ _3406_ _2926_ _2927_ VPWR VGND sg13g2_nor2_1
X_4284_ net1560 VPWR _0352_ VGND _3580_ _0351_ sg13g2_o21ai_1
X_7072_ net1258 VPWR _2863_ VGND _2811_ _2862_ sg13g2_o21ai_1
X_6023_ VGND VPWR net1393 _1921_ _1924_ _1923_ sg13g2_a21oi_1
X_6925_ net1270 VPWR _2734_ VGND _2663_ _2733_ sg13g2_o21ai_1
XFILLER_23_711 VPWR VGND sg13g2_fill_2
XFILLER_35_582 VPWR VGND sg13g2_fill_1
X_7919__88 VPWR VGND net88 sg13g2_tiehi
X_6856_ _2666_ net1270 _2665_ VPWR VGND sg13g2_nand2b_1
XFILLER_11_917 VPWR VGND sg13g2_fill_1
X_3999_ _3375_ net1440 VPWR VGND sg13g2_inv_2
XFILLER_23_777 VPWR VGND sg13g2_fill_2
X_5807_ VGND VPWR net1404 net726 _1726_ _1684_ sg13g2_a21oi_1
X_6787_ net1689 _2572_ _2609_ VPWR VGND sg13g2_nor2_1
X_5738_ _1663_ net1410 net819 VPWR VGND sg13g2_nand2_1
X_5669_ _0247_ _1601_ _1602_ _3470_ net1620 VPWR VGND sg13g2_a22oi_1
XFILLER_2_604 VPWR VGND sg13g2_fill_1
X_7408_ _3170_ net1678 _3169_ VPWR VGND sg13g2_nand2_1
X_7339_ _3104_ _3101_ _3103_ VPWR VGND sg13g2_nand2_1
Xhold461 s0.data_new_delayed\[0\] VPWR VGND net830 sg13g2_dlygate4sd3_1
Xhold450 s0.data_out\[14\]\[7\] VPWR VGND net819 sg13g2_dlygate4sd3_1
XFILLER_18_516 VPWR VGND sg13g2_fill_2
XFILLER_46_869 VPWR VGND sg13g2_decap_8
XFILLER_33_519 VPWR VGND sg13g2_decap_4
XFILLER_14_733 VPWR VGND sg13g2_fill_2
XFILLER_26_593 VPWR VGND sg13g2_fill_1
XFILLER_10_983 VPWR VGND sg13g2_decap_8
XFILLER_6_987 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_1_681 VPWR VGND sg13g2_decap_8
XFILLER_23_1012 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_49_696 VPWR VGND sg13g2_decap_8
XFILLER_36_368 VPWR VGND sg13g2_fill_2
XFILLER_17_560 VPWR VGND sg13g2_fill_2
X_4971_ s0.data_out\[20\]\[0\] s0.data_out\[21\]\[0\] net1492 _0969_ VPWR VGND sg13g2_mux2_1
X_6710_ _2535_ _2534_ _2533_ VPWR VGND sg13g2_nand2b_1
X_7690_ net336 VGND VPWR _0168_ s0.data_out\[23\]\[7\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_6641_ s0.data_out\[8\]\[7\] s0.data_out\[7\]\[7\] net1292 _2475_ VPWR VGND sg13g2_mux2_1
XFILLER_20_714 VPWR VGND sg13g2_fill_2
XFILLER_20_747 VPWR VGND sg13g2_fill_2
X_6572_ _2412_ VPWR _2413_ VGND net1731 net446 sg13g2_o21ai_1
X_5523_ VGND VPWR _1465_ _1467_ _1472_ net1683 sg13g2_a21oi_1
X_5454_ _1403_ net495 net1443 VPWR VGND sg13g2_nand2b_1
X_7953__334 VPWR VGND net334 sg13g2_tiehi
X_5385_ _1344_ net1439 _1345_ _1346_ VPWR VGND sg13g2_a21o_1
X_4405_ _0405_ _0460_ net1717 _0461_ VPWR VGND sg13g2_nand3_1
X_4336_ _0393_ net1541 net707 VPWR VGND sg13g2_nand2_1
X_7124_ s0.data_out\[4\]\[5\] s0.data_out\[3\]\[5\] net1245 _2910_ VPWR VGND sg13g2_mux2_1
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_1017 VPWR VGND sg13g2_decap_8
X_4267_ net1549 net1343 _3631_ VPWR VGND sg13g2_nor2b_1
X_7055_ net1250 s0.data_out\[4\]\[2\] _2850_ VPWR VGND sg13g2_and2_1
X_6006_ net1675 _1906_ _1907_ VPWR VGND sg13g2_nor2_1
X_4198_ _3386_ VPWR _3562_ VGND net1564 net464 sg13g2_o21ai_1
XFILLER_15_508 VPWR VGND sg13g2_fill_1
XFILLER_27_346 VPWR VGND sg13g2_decap_4
XFILLER_27_368 VPWR VGND sg13g2_fill_2
X_7957_ net282 VGND VPWR _0091_ s0.data_out\[1\]\[3\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_36_891 VPWR VGND sg13g2_fill_1
X_7888_ net122 VGND VPWR _0022_ s0.data_out\[7\]\[6\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_6908_ VGND VPWR net1265 _2717_ _2718_ _2715_ sg13g2_a21oi_1
X_6839_ _2652_ _2649_ _2651_ VPWR VGND sg13g2_nand2_1
XFILLER_24_45 VPWR VGND sg13g2_decap_4
XFILLER_6_206 VPWR VGND sg13g2_fill_1
XFILLER_40_44 VPWR VGND sg13g2_fill_2
XFILLER_3_935 VPWR VGND sg13g2_decap_8
XFILLER_46_1023 VPWR VGND sg13g2_decap_4
XFILLER_2_434 VPWR VGND sg13g2_decap_8
XFILLER_2_445 VPWR VGND sg13g2_fill_1
Xhold280 s0.data_out\[8\]\[1\] VPWR VGND net649 sg13g2_dlygate4sd3_1
Xhold291 _3295_ VPWR VGND net660 sg13g2_dlygate4sd3_1
X_7674__353 VPWR VGND net353 sg13g2_tiehi
Xfanout1714 net1717 net1714 VPWR VGND sg13g2_buf_8
Xfanout1703 net1704 net1703 VPWR VGND sg13g2_buf_8
Xfanout1725 net1728 net1725 VPWR VGND sg13g2_buf_8
Xfanout1736 net1737 net1736 VPWR VGND sg13g2_buf_8
Xfanout1747 net1750 net1747 VPWR VGND sg13g2_buf_8
XFILLER_46_688 VPWR VGND sg13g2_decap_8
XFILLER_34_839 VPWR VGND sg13g2_fill_1
XFILLER_5_294 VPWR VGND sg13g2_fill_1
X_5170_ net1607 _1073_ _1152_ VPWR VGND sg13g2_nor2_1
X_4121_ VPWR _3497_ net787 VGND sg13g2_inv_1
X_4052_ VPWR _3428_ net698 VGND sg13g2_inv_1
XFILLER_36_121 VPWR VGND sg13g2_fill_2
XFILLER_25_806 VPWR VGND sg13g2_fill_2
X_7811_ net205 VGND VPWR net451 s0.was_valid_out\[12\][0] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_7742_ net279 VGND VPWR _0220_ s0.shift_out\[18\][0] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_4954_ net1470 net1351 _0952_ VPWR VGND sg13g2_nor2b_1
XFILLER_17_390 VPWR VGND sg13g2_fill_2
X_4885_ net1486 net1346 _0894_ VPWR VGND sg13g2_nor2b_1
X_7673_ net354 VGND VPWR net602 s0.data_out\[24\]\[2\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_20_566 VPWR VGND sg13g2_fill_1
X_6624_ _2442_ _2456_ _2457_ _2458_ VPWR VGND sg13g2_nor3_1
X_6555_ _2399_ VPWR _2400_ VGND net1738 net661 sg13g2_o21ai_1
XFILLER_3_209 VPWR VGND sg13g2_fill_1
X_5506_ net1426 net1340 _1455_ VPWR VGND sg13g2_nor2b_1
X_6486_ VGND VPWR _2214_ _2331_ _2332_ net1307 sg13g2_a21oi_1
X_5437_ net1440 VPWR _1389_ VGND net1644 net1429 sg13g2_o21ai_1
X_5368_ _1329_ net585 net1456 VPWR VGND sg13g2_nand2b_1
X_4319_ _0377_ _0378_ _0379_ VPWR VGND sg13g2_nor2_1
X_5299_ _0213_ _1265_ _1266_ _3453_ net1617 VPWR VGND sg13g2_a22oi_1
X_7107_ VGND VPWR net1241 _2891_ _2893_ _2892_ sg13g2_a21oi_1
X_7038_ _2833_ VPWR _2836_ VGND net1680 _2825_ sg13g2_o21ai_1
XFILLER_28_699 VPWR VGND sg13g2_fill_2
XFILLER_42_124 VPWR VGND sg13g2_decap_8
XFILLER_42_168 VPWR VGND sg13g2_fill_2
XFILLER_35_99 VPWR VGND sg13g2_fill_2
XFILLER_7_526 VPWR VGND sg13g2_fill_1
XFILLER_4_0 VPWR VGND sg13g2_fill_1
XFILLER_3_798 VPWR VGND sg13g2_decap_8
XFILLER_2_253 VPWR VGND sg13g2_fill_1
XFILLER_2_264 VPWR VGND sg13g2_fill_2
Xfanout1533 net1536 net1533 VPWR VGND sg13g2_buf_8
Xfanout1500 net1502 net1500 VPWR VGND sg13g2_buf_8
Xfanout1522 net1527 net1522 VPWR VGND sg13g2_buf_1
Xfanout1511 net1514 net1511 VPWR VGND sg13g2_buf_1
Xfanout1555 s0.valid_out\[26\][0] net1555 VPWR VGND sg13g2_buf_1
Xfanout1544 net1548 net1544 VPWR VGND sg13g2_buf_8
Xfanout1566 net1569 net1566 VPWR VGND sg13g2_buf_8
XFILLER_47_920 VPWR VGND sg13g2_decap_8
Xfanout1577 net1578 net1577 VPWR VGND sg13g2_buf_8
Xfanout1588 net1603 net1588 VPWR VGND sg13g2_buf_8
XFILLER_19_633 VPWR VGND sg13g2_fill_2
Xfanout1599 net1602 net1599 VPWR VGND sg13g2_buf_1
XFILLER_20_1026 VPWR VGND sg13g2_fill_2
XFILLER_47_997 VPWR VGND sg13g2_decap_8
XFILLER_46_485 VPWR VGND sg13g2_fill_2
X_4670_ net1508 s0.data_out\[23\]\[4\] _0698_ VPWR VGND sg13g2_and2_1
X_6340_ net1637 net1343 _2202_ VPWR VGND sg13g2_nor2_1
X_6271_ _2146_ net1325 _2147_ _2148_ VPWR VGND sg13g2_a21o_1
X_5222_ _1195_ net1459 _1194_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_0 VPWR VGND sg13g2_decap_4
X_5153_ _1124_ net1683 _1138_ VPWR VGND _1132_ sg13g2_nand3b_1
X_4104_ VPWR _3480_ net730 VGND sg13g2_inv_1
X_5084_ s0.data_out\[20\]\[2\] s0.data_out\[19\]\[2\] net1464 _1069_ VPWR VGND sg13g2_mux2_1
X_4035_ VPWR _3411_ net1347 VGND sg13g2_inv_1
XFILLER_38_986 VPWR VGND sg13g2_decap_8
XFILLER_40_617 VPWR VGND sg13g2_fill_1
XFILLER_36_1000 VPWR VGND sg13g2_decap_8
X_5986_ VGND VPWR _1769_ _1886_ _1887_ net1391 sg13g2_a21oi_1
X_4937_ net1498 VPWR _0938_ VGND _0869_ _0937_ sg13g2_o21ai_1
X_7725_ net298 VGND VPWR _0203_ s0.data_out\[20\]\[6\] clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_21_831 VPWR VGND sg13g2_fill_1
X_7656_ net28 VGND VPWR _0134_ s0.valid_out\[25\][0] clknet_leaf_43_clk sg13g2_dfrbpq_2
X_4868_ _0875_ net1482 _0876_ _0877_ VPWR VGND sg13g2_a21o_1
XFILLER_21_842 VPWR VGND sg13g2_fill_1
X_6607_ VGND VPWR net1293 _2438_ _2441_ _2440_ sg13g2_a21oi_1
X_7587_ net439 net1216 net1212 _3325_ VPWR VGND sg13g2_a21o_1
X_4799_ VGND VPWR net1494 net755 _0814_ _0773_ sg13g2_a21oi_1
XFILLER_4_507 VPWR VGND sg13g2_fill_1
X_6538_ _2384_ _2383_ net1306 VPWR VGND sg13g2_nand2b_1
X_6469_ net1741 VPWR _2318_ VGND _2315_ _2317_ sg13g2_o21ai_1
XFILLER_43_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_768 VPWR VGND sg13g2_decap_8
X_7671__356 VPWR VGND net356 sg13g2_tiehi
XFILLER_48_739 VPWR VGND sg13g2_decap_8
XFILLER_29_931 VPWR VGND sg13g2_fill_2
XFILLER_46_32 VPWR VGND sg13g2_fill_2
XFILLER_28_452 VPWR VGND sg13g2_fill_1
XFILLER_28_463 VPWR VGND sg13g2_fill_1
X_7849__164 VPWR VGND net164 sg13g2_tiehi
XFILLER_44_967 VPWR VGND sg13g2_decap_8
XFILLER_12_820 VPWR VGND sg13g2_fill_2
XFILLER_30_127 VPWR VGND sg13g2_fill_2
XFILLER_8_868 VPWR VGND sg13g2_fill_2
X_7655__30 VPWR VGND net30 sg13g2_tiehi
Xfanout1330 net1332 net1330 VPWR VGND sg13g2_buf_8
Xfanout1341 net1342 net1341 VPWR VGND sg13g2_buf_8
Xfanout1374 s0.valid_out\[11\][0] net1374 VPWR VGND sg13g2_buf_8
Xfanout1363 net1364 net1363 VPWR VGND sg13g2_buf_2
Xfanout1352 net1353 net1352 VPWR VGND sg13g2_buf_8
Xfanout1396 net729 net1396 VPWR VGND sg13g2_buf_2
XFILLER_38_249 VPWR VGND sg13g2_fill_2
Xfanout1385 s0.shift_out\[12\][0] net1385 VPWR VGND sg13g2_buf_1
XFILLER_47_794 VPWR VGND sg13g2_decap_8
X_5840_ VGND VPWR _1753_ _1752_ net1698 sg13g2_or2_1
XFILLER_21_127 VPWR VGND sg13g2_fill_2
X_5771_ _1696_ net1196 _1695_ VPWR VGND sg13g2_nand2_1
X_7510_ s0.data_out\[0\]\[5\] s0.data_out\[1\]\[5\] net1227 _3260_ VPWR VGND sg13g2_mux2_1
X_4722_ _0742_ VPWR _0743_ VGND net1504 _3434_ sg13g2_o21ai_1
X_7441_ _3196_ VPWR _3197_ VGND net1188 _3195_ sg13g2_o21ai_1
X_4653_ net1510 s0.data_out\[23\]\[0\] _0685_ VPWR VGND sg13g2_and2_1
X_7372_ _3134_ net614 net1237 VPWR VGND sg13g2_nand2b_1
X_4584_ VGND VPWR _0510_ _0616_ _0617_ net1525 sg13g2_a21oi_1
X_6323_ _2189_ VPWR _2191_ VGND s0.was_valid_out\[9\][0] net1317 sg13g2_o21ai_1
X_6254_ VGND VPWR _2013_ _2130_ _2131_ net1368 sg13g2_a21oi_1
X_5205_ s0.data_out\[19\]\[2\] s0.data_out\[18\]\[2\] net1453 _1178_ VPWR VGND sg13g2_mux2_1
X_6185_ net1379 VPWR _2068_ VGND _2026_ _2067_ sg13g2_o21ai_1
X_5136_ _1119_ net1457 _1120_ _1121_ VPWR VGND sg13g2_a21o_1
X_5067_ net1604 _0989_ _1057_ VPWR VGND sg13g2_nor2_1
X_4018_ net1294 _3394_ VPWR VGND sg13g2_inv_4
X_7961__230 VPWR VGND net230 sg13g2_tiehi
XFILLER_41_926 VPWR VGND sg13g2_decap_8
XFILLER_25_455 VPWR VGND sg13g2_fill_2
X_5969_ _1754_ VPWR _1870_ VGND net1397 _3491_ sg13g2_o21ai_1
X_7708_ net316 VGND VPWR _0186_ s0.data_out\[21\]\[2\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_7639_ net47 VGND VPWR net470 s0.data_out\[27\]\[4\] clknet_leaf_44_clk sg13g2_dfrbpq_2
XFILLER_10_1025 VPWR VGND sg13g2_decap_4
XFILLER_4_359 VPWR VGND sg13g2_fill_1
XFILLER_0_554 VPWR VGND sg13g2_fill_2
XFILLER_48_536 VPWR VGND sg13g2_fill_2
X_7652__33 VPWR VGND net33 sg13g2_tiehi
XFILLER_36_709 VPWR VGND sg13g2_fill_2
XFILLER_28_271 VPWR VGND sg13g2_fill_2
X_7862__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_31_447 VPWR VGND sg13g2_fill_1
Xhold109 s0.data_out\[24\]\[3\] VPWR VGND net478 sg13g2_dlygate4sd3_1
X_7719__304 VPWR VGND net304 sg13g2_tiehi
XFILLER_4_871 VPWR VGND sg13g2_decap_8
Xfanout1182 net1183 net1182 VPWR VGND sg13g2_buf_8
Xfanout1171 net1172 net1171 VPWR VGND sg13g2_buf_1
XFILLER_26_208 VPWR VGND sg13g2_fill_2
Xfanout1193 net1194 net1193 VPWR VGND sg13g2_buf_1
XFILLER_47_591 VPWR VGND sg13g2_fill_2
XFILLER_19_260 VPWR VGND sg13g2_fill_2
X_6941_ _0031_ _2745_ _2746_ _3521_ net1597 VPWR VGND sg13g2_a22oi_1
X_6872_ VGND VPWR _2566_ _2681_ _2682_ net1273 sg13g2_a21oi_1
X_5823_ VPWR _1739_ _1738_ VGND sg13g2_inv_1
XFILLER_22_436 VPWR VGND sg13g2_fill_1
X_5754_ VGND VPWR _1679_ _1669_ net1655 sg13g2_or2_1
X_4705_ _0726_ net1182 _0725_ VPWR VGND sg13g2_nand2_1
X_5685_ _1614_ VPWR _1615_ VGND net1744 net742 sg13g2_o21ai_1
XFILLER_31_992 VPWR VGND sg13g2_decap_8
X_4636_ net1508 net1339 _0669_ VPWR VGND sg13g2_nor2b_1
X_7424_ _3183_ VPWR _3184_ VGND net1718 net750 sg13g2_o21ai_1
X_7355_ _2992_ VPWR _3117_ VGND net1235 _3542_ sg13g2_o21ai_1
X_6306_ net1325 net493 _2177_ VPWR VGND sg13g2_and2_1
X_4567_ net1524 VPWR _0603_ VGND net1641 net1509 sg13g2_o21ai_1
XFILLER_2_819 VPWR VGND sg13g2_decap_8
X_7839__174 VPWR VGND net174 sg13g2_tiehi
X_4498_ VGND VPWR net1537 _0540_ _0543_ _0542_ sg13g2_a21oi_1
X_7286_ net1686 _3021_ _3060_ VPWR VGND sg13g2_nor2_1
X_6237_ _2114_ net443 net1373 VPWR VGND sg13g2_nand2b_1
X_6168_ net1376 VPWR _2055_ VGND _1982_ _2054_ sg13g2_o21ai_1
XFILLER_40_1018 VPWR VGND sg13g2_decap_8
X_5119_ _1104_ net645 net1480 VPWR VGND sg13g2_nand2b_1
X_6099_ VGND VPWR net1376 _1985_ _1988_ _1987_ sg13g2_a21oi_1
XFILLER_45_539 VPWR VGND sg13g2_fill_1
XFILLER_27_78 VPWR VGND sg13g2_fill_2
XFILLER_40_200 VPWR VGND sg13g2_fill_2
X_7846__167 VPWR VGND net167 sg13g2_tiehi
XFILLER_41_767 VPWR VGND sg13g2_fill_1
XFILLER_40_299 VPWR VGND sg13g2_fill_2
XFILLER_49_801 VPWR VGND sg13g2_decap_8
XFILLER_1_852 VPWR VGND sg13g2_decap_8
XFILLER_0_384 VPWR VGND sg13g2_decap_8
XFILLER_0_395 VPWR VGND sg13g2_fill_1
XFILLER_49_878 VPWR VGND sg13g2_decap_8
XFILLER_16_230 VPWR VGND sg13g2_fill_1
X_7928__78 VPWR VGND net78 sg13g2_tiehi
XFILLER_9_974 VPWR VGND sg13g2_decap_8
X_5470_ _1418_ VPWR _1419_ VGND net1206 _1416_ sg13g2_o21ai_1
X_4421_ net1550 VPWR _0473_ VGND _0438_ _0472_ sg13g2_o21ai_1
X_4352_ _0408_ VPWR _0409_ VGND net1541 _3409_ sg13g2_o21ai_1
X_7140_ _2925_ VPWR _2926_ VGND net1173 _2923_ sg13g2_o21ai_1
X_4283_ net1546 s0.data_out\[26\]\[0\] _0351_ VPWR VGND sg13g2_and2_1
X_7071_ net1173 _3532_ _2862_ VPWR VGND sg13g2_nor2_1
X_6022_ VGND VPWR _1778_ _1922_ _1923_ net1392 sg13g2_a21oi_1
XFILLER_39_366 VPWR VGND sg13g2_fill_1
XFILLER_27_506 VPWR VGND sg13g2_decap_4
X_7973_ net29 VGND VPWR _0107_ s0.data_out\[0\]\[7\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_6924_ net1262 s0.data_out\[5\]\[0\] _2733_ VPWR VGND sg13g2_and2_1
X_6855_ VGND VPWR net1262 _2664_ _2665_ _2663_ sg13g2_a21oi_1
X_6786_ _2605_ _2607_ net1670 _2608_ VPWR VGND sg13g2_nand3_1
XFILLER_13_14 VPWR VGND sg13g2_decap_8
X_3998_ VPWR _3374_ net1735 VGND sg13g2_inv_1
X_5806_ VPWR _0261_ _1725_ VGND sg13g2_inv_1
X_5737_ _1661_ VPWR _1662_ VGND _1649_ _1659_ sg13g2_o21ai_1
X_7407_ VGND VPWR net1233 _3166_ _3169_ _3168_ sg13g2_a21oi_1
X_5668_ net1620 _1523_ _1602_ VPWR VGND sg13g2_nor2_1
X_4619_ s0.data_out\[24\]\[6\] s0.data_out\[23\]\[6\] net1515 _0652_ VPWR VGND sg13g2_mux2_1
X_5599_ VGND VPWR net1412 _1534_ _1536_ _1535_ sg13g2_a21oi_1
Xhold462 s0.valid_out\[13\][0] VPWR VGND net831 sg13g2_dlygate4sd3_1
Xhold451 s0.valid_out\[18\][0] VPWR VGND net820 sg13g2_dlygate4sd3_1
Xhold440 _1368_ VPWR VGND net809 sg13g2_dlygate4sd3_1
X_7338_ net1187 VPWR _3103_ VGND s0.was_valid_out\[1\][0] net1235 sg13g2_o21ai_1
X_7269_ _3042_ VPWR _3043_ VGND net1237 _3536_ sg13g2_o21ai_1
XFILLER_46_848 VPWR VGND sg13g2_decap_8
XFILLER_13_200 VPWR VGND sg13g2_fill_1
XFILLER_41_531 VPWR VGND sg13g2_fill_1
XFILLER_9_204 VPWR VGND sg13g2_fill_2
XFILLER_6_966 VPWR VGND sg13g2_decap_8
XFILLER_5_465 VPWR VGND sg13g2_fill_2
X_7716__307 VPWR VGND net307 sg13g2_tiehi
XFILLER_1_660 VPWR VGND sg13g2_fill_2
XFILLER_0_170 VPWR VGND sg13g2_fill_2
XFILLER_49_675 VPWR VGND sg13g2_decap_8
XFILLER_36_325 VPWR VGND sg13g2_fill_1
X_4970_ VGND VPWR net1470 _0966_ _0968_ _0967_ sg13g2_a21oi_1
X_6640_ _2474_ net1291 net414 VPWR VGND sg13g2_nand2_1
X_6571_ _2384_ _2411_ net1731 _2412_ VPWR VGND sg13g2_nand3_1
X_5522_ VPWR _1471_ _1470_ VGND sg13g2_inv_1
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
X_5453_ _1400_ net1423 _1401_ _1402_ VPWR VGND sg13g2_a21o_1
X_5384_ net1439 net1341 _1345_ VPWR VGND sg13g2_nor2b_1
X_4404_ net1551 VPWR _0460_ VGND _0401_ _0459_ sg13g2_o21ai_1
X_7836__177 VPWR VGND net177 sg13g2_tiehi
XFILLER_5_81 VPWR VGND sg13g2_fill_2
X_4335_ VGND VPWR _0392_ _0391_ net1695 sg13g2_or2_1
X_7123_ _2909_ net1245 net503 VPWR VGND sg13g2_nand2_1
X_4266_ s0.data_out\[27\]\[4\] s0.data_out\[26\]\[4\] net1554 _3630_ VPWR VGND sg13g2_mux2_1
X_7054_ _0041_ _2848_ _2849_ _3530_ net1590 VPWR VGND sg13g2_a22oi_1
XFILLER_39_130 VPWR VGND sg13g2_fill_2
X_6005_ VGND VPWR net1392 _1903_ _1906_ _1905_ sg13g2_a21oi_1
X_4197_ net1714 net370 _0111_ VPWR VGND sg13g2_and2_1
XFILLER_39_185 VPWR VGND sg13g2_fill_1
XFILLER_39_174 VPWR VGND sg13g2_fill_2
XFILLER_27_314 VPWR VGND sg13g2_fill_2
XFILLER_27_325 VPWR VGND sg13g2_fill_2
X_7956_ net295 VGND VPWR _0090_ s0.data_out\[1\]\[2\] clknet_leaf_11_clk sg13g2_dfrbpq_2
XFILLER_39_1020 VPWR VGND sg13g2_decap_8
X_7887_ net123 VGND VPWR _0021_ s0.data_out\[7\]\[5\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_6907_ s0.data_out\[6\]\[4\] s0.data_out\[5\]\[4\] net1269 _2717_ VPWR VGND sg13g2_mux2_1
X_7667__361 VPWR VGND net361 sg13g2_tiehi
XFILLER_35_391 VPWR VGND sg13g2_fill_2
X_6838_ net1174 VPWR _2651_ VGND s0.was_valid_out\[5\][0] net1280 sg13g2_o21ai_1
X_6769_ VGND VPWR _2591_ _2588_ net1661 sg13g2_or2_1
X_7915__92 VPWR VGND net92 sg13g2_tiehi
XFILLER_3_914 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_46_1002 VPWR VGND sg13g2_decap_8
Xhold270 s0.data_out\[11\]\[5\] VPWR VGND net639 sg13g2_dlygate4sd3_1
XFILLER_6_4 VPWR VGND sg13g2_fill_1
Xfanout1715 net1717 net1715 VPWR VGND sg13g2_buf_1
Xfanout1704 ui_in[1] net1704 VPWR VGND sg13g2_buf_8
Xhold292 s0.data_out\[9\]\[0\] VPWR VGND net661 sg13g2_dlygate4sd3_1
Xhold281 _0005_ VPWR VGND net650 sg13g2_dlygate4sd3_1
Xfanout1726 net1728 net1726 VPWR VGND sg13g2_buf_1
Xfanout1737 net1751 net1737 VPWR VGND sg13g2_buf_8
Xfanout1748 net1749 net1748 VPWR VGND sg13g2_buf_8
XFILLER_14_575 VPWR VGND sg13g2_fill_1
XFILLER_41_394 VPWR VGND sg13g2_fill_1
XFILLER_5_240 VPWR VGND sg13g2_fill_1
X_4120_ VPWR _3496_ net639 VGND sg13g2_inv_1
XFILLER_2_980 VPWR VGND sg13g2_decap_8
X_4051_ VPWR _3427_ net407 VGND sg13g2_inv_1
X_7810_ net206 VGND VPWR net576 s0.data_out\[13\]\[7\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_7907__101 VPWR VGND net101 sg13g2_tiehi
XFILLER_24_306 VPWR VGND sg13g2_fill_1
X_7741_ net280 VGND VPWR _0219_ s0.genblk1\[17\].modules.bubble clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
X_4953_ _0950_ VPWR _0951_ VGND net1478 _3444_ sg13g2_o21ai_1
XFILLER_24_328 VPWR VGND sg13g2_fill_2
X_7672_ net355 VGND VPWR net482 s0.data_out\[24\]\[1\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_4884_ _0890_ _0892_ net1673 _0893_ VPWR VGND sg13g2_nand3_1
X_6623_ VPWR VGND _2455_ net1711 _2453_ net1709 _2457_ _2449_ sg13g2_a221oi_1
X_6554_ _2339_ _2398_ net1738 _2399_ VPWR VGND sg13g2_nand3_1
XFILLER_9_590 VPWR VGND sg13g2_fill_2
X_5505_ s0.data_out\[17\]\[5\] s0.data_out\[16\]\[5\] net1433 _1454_ VPWR VGND sg13g2_mux2_1
X_6485_ _2331_ s0.data_out\[8\]\[1\] net1314 VPWR VGND sg13g2_nand2b_1
X_5436_ _0228_ _1387_ _1388_ _3457_ net1624 VPWR VGND sg13g2_a22oi_1
XFILLER_10_48 VPWR VGND sg13g2_fill_1
X_5367_ _1326_ net1441 _1327_ _1328_ VPWR VGND sg13g2_a21o_1
X_5298_ net1617 _1240_ _1266_ VPWR VGND sg13g2_nor2_1
X_4318_ VGND VPWR net1633 net1556 _0378_ net1549 sg13g2_a21oi_1
XFILLER_19_13 VPWR VGND sg13g2_decap_8
X_7106_ net1240 net1356 _2892_ VPWR VGND sg13g2_nor2b_1
X_4249_ _3613_ _3612_ net1658 _3604_ net1647 VPWR VGND sg13g2_a22oi_1
X_7037_ net1670 _2832_ _2835_ VPWR VGND sg13g2_nor2_1
X_7939_ net66 VGND VPWR _0073_ s0.valid_out\[2\][0] clknet_leaf_8_clk sg13g2_dfrbpq_2
XFILLER_24_862 VPWR VGND sg13g2_fill_1
XFILLER_11_523 VPWR VGND sg13g2_fill_2
XFILLER_13_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_777 VPWR VGND sg13g2_decap_8
Xfanout1512 net1513 net1512 VPWR VGND sg13g2_buf_8
Xfanout1523 net1524 net1523 VPWR VGND sg13g2_buf_8
Xfanout1501 net1502 net1501 VPWR VGND sg13g2_buf_1
Xfanout1556 net1557 net1556 VPWR VGND sg13g2_buf_2
Xfanout1534 net1536 net1534 VPWR VGND sg13g2_buf_1
Xfanout1545 net1548 net1545 VPWR VGND sg13g2_buf_1
Xfanout1589 net1592 net1589 VPWR VGND sg13g2_buf_8
Xfanout1578 net1588 net1578 VPWR VGND sg13g2_buf_8
Xfanout1567 net1569 net1567 VPWR VGND sg13g2_buf_8
XFILLER_47_976 VPWR VGND sg13g2_decap_8
XFILLER_46_420 VPWR VGND sg13g2_fill_2
XFILLER_20_1005 VPWR VGND sg13g2_decap_8
XFILLER_33_103 VPWR VGND sg13g2_fill_1
XFILLER_34_637 VPWR VGND sg13g2_fill_2
XFILLER_42_670 VPWR VGND sg13g2_fill_2
XFILLER_14_361 VPWR VGND sg13g2_fill_1
X_6270_ net1325 net1340 _2147_ VPWR VGND sg13g2_nor2b_1
X_5221_ VGND VPWR net1447 _1192_ _1194_ _1193_ sg13g2_a21oi_1
X_5152_ _1137_ _1099_ _1136_ VPWR VGND sg13g2_nand2_1
X_4103_ VPWR _3479_ net612 VGND sg13g2_inv_1
X_5083_ _1068_ net1467 net634 VPWR VGND sg13g2_nand2_1
XFILLER_38_965 VPWR VGND sg13g2_decap_8
X_4034_ _3410_ net448 VPWR VGND sg13g2_inv_2
XFILLER_37_486 VPWR VGND sg13g2_fill_1
X_7724_ net299 VGND VPWR net510 s0.data_out\[20\]\[5\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_5985_ _1886_ net597 net1397 VPWR VGND sg13g2_nand2b_1
X_4936_ net1180 _3441_ _0937_ VPWR VGND sg13g2_nor2_1
X_7655_ net30 VGND VPWR net420 s0.was_valid_out\[25\][0] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_7664__364 VPWR VGND net364 sg13g2_tiehi
X_4867_ net1482 net1335 _0876_ VPWR VGND sg13g2_nor2b_1
X_7586_ _3402_ _3319_ _3324_ VPWR VGND sg13g2_nor2_1
X_6606_ VGND VPWR _2319_ _2439_ _2440_ net1293 sg13g2_a21oi_1
X_4798_ VPWR _0165_ _0813_ VGND sg13g2_inv_1
X_6537_ _2255_ VPWR _2383_ VGND net1314 _3510_ sg13g2_o21ai_1
X_6468_ _2314_ VPWR _2317_ VGND net1310 _2316_ sg13g2_o21ai_1
X_5419_ _0224_ _1374_ _1375_ _3460_ net1618 VPWR VGND sg13g2_a22oi_1
X_6399_ net1312 net1346 _2257_ VPWR VGND sg13g2_nor2b_1
XFILLER_43_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_747 VPWR VGND sg13g2_decap_8
XFILLER_48_718 VPWR VGND sg13g2_decap_8
XFILLER_16_615 VPWR VGND sg13g2_fill_1
XFILLER_44_946 VPWR VGND sg13g2_decap_8
XFILLER_7_324 VPWR VGND sg13g2_decap_4
XFILLER_7_313 VPWR VGND sg13g2_fill_1
XFILLER_7_27 VPWR VGND sg13g2_fill_2
Xfanout1331 net1332 net1331 VPWR VGND sg13g2_buf_8
Xfanout1320 net1327 net1320 VPWR VGND sg13g2_buf_8
Xfanout1364 s0.valid_out\[10\][0] net1364 VPWR VGND sg13g2_buf_2
Xfanout1375 s0.valid_out\[11\][0] net1375 VPWR VGND sg13g2_buf_2
Xfanout1353 s0.data_new_delayed\[1\] net1353 VPWR VGND sg13g2_buf_8
Xfanout1342 s0.data_new_delayed\[5\] net1342 VPWR VGND sg13g2_buf_8
Xfanout1386 net1388 net1386 VPWR VGND sg13g2_buf_8
Xfanout1397 net1398 net1397 VPWR VGND sg13g2_buf_8
XFILLER_47_773 VPWR VGND sg13g2_decap_8
XFILLER_22_607 VPWR VGND sg13g2_fill_1
X_7904__104 VPWR VGND net104 sg13g2_tiehi
X_5770_ _1568_ VPWR _1695_ VGND net1420 _3478_ sg13g2_o21ai_1
X_4721_ _0742_ net1504 net530 VPWR VGND sg13g2_nand2_1
X_7440_ VGND VPWR net1189 _3158_ _3196_ net1586 sg13g2_a21oi_1
X_4652_ VGND VPWR _0680_ _0683_ _0148_ _0684_ sg13g2_a21oi_1
X_7371_ _3131_ net1221 _3132_ _3133_ VPWR VGND sg13g2_a21o_1
X_4583_ _0616_ s0.data_out\[23\]\[2\] net1531 VPWR VGND sg13g2_nand2b_1
X_6322_ VPWR _2190_ _2189_ VGND sg13g2_inv_1
X_6253_ _2130_ net522 net1374 VPWR VGND sg13g2_nand2b_1
X_5204_ _1177_ net1454 s0.data_out\[18\]\[2\] VPWR VGND sg13g2_nand2_1
X_6184_ _3383_ _3496_ _2067_ VPWR VGND sg13g2_nor2_1
X_5135_ net1457 net1345 _1120_ VPWR VGND sg13g2_nor2b_1
X_5066_ net1483 VPWR _1056_ VGND _0986_ _1055_ sg13g2_o21ai_1
X_4017_ net1210 _3393_ VPWR VGND sg13g2_inv_4
XFILLER_16_47 VPWR VGND sg13g2_fill_1
X_5968_ _1869_ net1390 _1868_ VPWR VGND sg13g2_nand2b_1
X_4919_ net1500 VPWR _0924_ VGND _0858_ _0923_ sg13g2_o21ai_1
X_7707_ net317 VGND VPWR _0185_ s0.data_out\[21\]\[1\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_5899_ net1675 _1810_ _1812_ VPWR VGND sg13g2_nor2_1
XFILLER_32_46 VPWR VGND sg13g2_fill_1
X_7638_ net48 VGND VPWR _0116_ s0.data_out\[27\]\[3\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_7569_ VPWR _0094_ _3311_ VGND sg13g2_inv_1
XFILLER_10_1004 VPWR VGND sg13g2_decap_8
XFILLER_17_913 VPWR VGND sg13g2_fill_1
XFILLER_16_445 VPWR VGND sg13g2_decap_4
XFILLER_43_253 VPWR VGND sg13g2_fill_2
XFILLER_31_415 VPWR VGND sg13g2_fill_1
XFILLER_32_949 VPWR VGND sg13g2_fill_2
XFILLER_8_644 VPWR VGND sg13g2_fill_2
XFILLER_8_633 VPWR VGND sg13g2_fill_2
XFILLER_11_161 VPWR VGND sg13g2_fill_2
XFILLER_39_526 VPWR VGND sg13g2_fill_1
Xfanout1183 _3390_ net1183 VPWR VGND sg13g2_buf_8
Xfanout1172 net1173 net1172 VPWR VGND sg13g2_buf_2
Xfanout1194 _3382_ net1194 VPWR VGND sg13g2_buf_8
X_6940_ net1596 _2682_ _2746_ VPWR VGND sg13g2_nor2_1
XFILLER_47_581 VPWR VGND sg13g2_fill_1
XFILLER_23_916 VPWR VGND sg13g2_fill_2
X_6871_ _2681_ net693 net1279 VPWR VGND sg13g2_nand2b_1
X_5822_ VGND VPWR net1635 net1399 _1738_ _1737_ sg13g2_a21oi_1
X_5753_ net1665 _1676_ _1678_ VPWR VGND sg13g2_nor2_1
X_4704_ s0.data_out\[22\]\[0\] s0.data_out\[23\]\[0\] net1517 _0725_ VPWR VGND sg13g2_mux2_1
XFILLER_31_971 VPWR VGND sg13g2_decap_8
X_7661__367 VPWR VGND net367 sg13g2_tiehi
X_5684_ _1613_ net1744 _1614_ VPWR VGND _1562_ sg13g2_nand3b_1
X_4635_ s0.data_out\[24\]\[5\] s0.data_out\[23\]\[5\] net1515 _0668_ VPWR VGND sg13g2_mux2_1
X_7423_ _3182_ VPWR _3183_ VGND net1187 _3181_ sg13g2_o21ai_1
X_4566_ _0144_ _0601_ _0602_ _3424_ net1579 VPWR VGND sg13g2_a22oi_1
X_7354_ _3116_ net1230 _3115_ VPWR VGND sg13g2_nand2b_1
X_6305_ _0309_ _2175_ _2176_ _3497_ net1612 VPWR VGND sg13g2_a22oi_1
X_4497_ VGND VPWR _0417_ _0541_ _0542_ net1537 sg13g2_a21oi_1
X_7285_ _3059_ _3058_ net1678 _3048_ net1669 VPWR VGND sg13g2_a22oi_1
X_6236_ _2111_ net1322 _2112_ _2113_ VPWR VGND sg13g2_a21o_1
X_6167_ _3383_ _3492_ _2054_ VPWR VGND sg13g2_nor2_1
X_5118_ _1101_ net1457 _1102_ _1103_ VPWR VGND sg13g2_a21o_1
X_6098_ VGND VPWR _1865_ _1986_ _1987_ net1376 sg13g2_a21oi_1
X_5049_ net1605 _0979_ _1043_ VPWR VGND sg13g2_nor2_1
XFILLER_26_710 VPWR VGND sg13g2_decap_4
XFILLER_13_415 VPWR VGND sg13g2_fill_1
XFILLER_43_67 VPWR VGND sg13g2_fill_1
XFILLER_49_1011 VPWR VGND sg13g2_decap_8
XFILLER_1_831 VPWR VGND sg13g2_decap_8
XFILLER_49_857 VPWR VGND sg13g2_decap_8
XFILLER_1_1013 VPWR VGND sg13g2_decap_8
XFILLER_29_570 VPWR VGND sg13g2_decap_4
XFILLER_16_220 VPWR VGND sg13g2_fill_1
XFILLER_44_595 VPWR VGND sg13g2_fill_2
XFILLER_32_779 VPWR VGND sg13g2_decap_8
X_4420_ net1534 net431 _0472_ VPWR VGND sg13g2_and2_1
X_4351_ _0408_ net1541 net501 VPWR VGND sg13g2_nand2_1
X_7070_ _0045_ _2860_ _2861_ _3526_ net1596 VPWR VGND sg13g2_a22oi_1
X_4282_ VGND VPWR _0344_ _0348_ _0112_ _0350_ sg13g2_a21oi_1
X_6021_ _1922_ net540 net1399 VPWR VGND sg13g2_nand2b_1
XFILLER_12_0 VPWR VGND sg13g2_fill_1
X_7972_ net67 VGND VPWR _0106_ s0.data_out\[0\]\[6\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_6923_ VGND VPWR _2728_ _2731_ _0027_ _2732_ sg13g2_a21oi_1
XFILLER_23_713 VPWR VGND sg13g2_fill_1
XFILLER_35_573 VPWR VGND sg13g2_decap_8
XFILLER_22_212 VPWR VGND sg13g2_fill_2
X_6854_ s0.data_out\[6\]\[0\] s0.data_out\[5\]\[0\] net1269 _2664_ VPWR VGND sg13g2_mux2_1
X_6785_ _2607_ _3395_ _2606_ VPWR VGND sg13g2_nand2_1
X_3997_ VPWR _3373_ net1644 VGND sg13g2_inv_1
X_5805_ _1724_ VPWR _1725_ VGND net1748 net777 sg13g2_o21ai_1
X_5736_ _1661_ net1693 _1658_ VPWR VGND sg13g2_nand2_1
X_5667_ net1424 VPWR _1601_ VGND _1520_ _1600_ sg13g2_o21ai_1
X_7406_ VGND VPWR _3052_ _3167_ _3168_ net1232 sg13g2_a21oi_1
X_4618_ _0651_ net1516 net579 VPWR VGND sg13g2_nand2_1
X_5598_ net1412 net1358 _1535_ VPWR VGND sg13g2_nor2b_1
Xhold463 s0.data_out\[9\]\[6\] VPWR VGND net832 sg13g2_dlygate4sd3_1
Xhold430 s0.data_out\[1\]\[0\] VPWR VGND net799 sg13g2_dlygate4sd3_1
Xhold452 s0.was_valid_out\[18\][0] VPWR VGND net821 sg13g2_dlygate4sd3_1
X_4549_ VGND VPWR net1184 _0562_ _0589_ net1589 sg13g2_a21oi_1
Xhold441 s0.data_out\[23\]\[3\] VPWR VGND net810 sg13g2_dlygate4sd3_1
X_7337_ net1218 _3096_ _3102_ VPWR VGND sg13g2_nor2_1
X_7268_ _3042_ net1238 s0.data_out\[2\]\[5\] VPWR VGND sg13g2_nand2_1
X_7852__161 VPWR VGND net161 sg13g2_tiehi
X_6219_ _2095_ VPWR _2096_ VGND net1361 _3492_ sg13g2_o21ai_1
X_7199_ net1248 VPWR _2978_ VGND _2938_ _2977_ sg13g2_o21ai_1
XFILLER_18_507 VPWR VGND sg13g2_fill_1
XFILLER_46_827 VPWR VGND sg13g2_decap_8
X_7709__315 VPWR VGND net315 sg13g2_tiehi
XFILLER_26_562 VPWR VGND sg13g2_fill_2
XFILLER_41_598 VPWR VGND sg13g2_fill_2
XFILLER_9_238 VPWR VGND sg13g2_fill_2
XFILLER_6_945 VPWR VGND sg13g2_decap_8
XFILLER_5_422 VPWR VGND sg13g2_fill_2
XFILLER_49_654 VPWR VGND sg13g2_decap_8
XFILLER_45_893 VPWR VGND sg13g2_decap_8
X_7829__185 VPWR VGND net185 sg13g2_tiehi
XFILLER_20_749 VPWR VGND sg13g2_fill_1
X_6570_ net1306 VPWR _2411_ VGND _2378_ _2410_ sg13g2_o21ai_1
X_5521_ VGND VPWR _1457_ _1459_ _1470_ net1674 sg13g2_a21oi_1
XFILLER_30_1007 VPWR VGND sg13g2_decap_8
X_5452_ net1423 net1354 _1401_ VPWR VGND sg13g2_nor2b_1
X_5383_ s0.data_out\[18\]\[5\] s0.data_out\[17\]\[5\] net1445 _1344_ VPWR VGND sg13g2_mux2_1
X_4403_ net1186 _3420_ _0459_ VPWR VGND sg13g2_nor2_1
X_4334_ VGND VPWR net1551 _0388_ _0391_ _0390_ sg13g2_a21oi_1
X_7122_ _2907_ VPWR _2908_ VGND net1571 _2883_ sg13g2_o21ai_1
X_7053_ net1590 _2783_ _2849_ VPWR VGND sg13g2_nor2_1
X_6004_ VGND VPWR _1804_ _1904_ _1905_ net1392 sg13g2_a21oi_1
X_4265_ _3629_ net1556 net517 VPWR VGND sg13g2_nand2_1
X_4196_ net1575 _3556_ _0110_ VPWR VGND sg13g2_nor2_1
X_7955_ net308 VGND VPWR _0089_ s0.data_out\[1\]\[1\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_6906_ _2716_ net1269 net668 VPWR VGND sg13g2_nand2_1
X_7886_ net124 VGND VPWR _0020_ s0.data_out\[7\]\[4\] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_6837_ net1264 _2646_ _2650_ VPWR VGND sg13g2_nor2_1
X_6768_ VGND VPWR _2590_ _2581_ net1651 sg13g2_or2_1
X_7958__269 VPWR VGND net269 sg13g2_tiehi
X_6699_ _0009_ _2525_ _2526_ _3509_ net1600 VPWR VGND sg13g2_a22oi_1
X_5719_ net1401 net1350 _1644_ VPWR VGND sg13g2_nor2b_1
Xhold271 _0310_ VPWR VGND net640 sg13g2_dlygate4sd3_1
Xhold260 s0.data_out\[21\]\[1\] VPWR VGND net629 sg13g2_dlygate4sd3_1
Xhold282 s0.was_valid_out\[20\][0] VPWR VGND net651 sg13g2_dlygate4sd3_1
Xhold293 s0.data_out\[23\]\[7\] VPWR VGND net662 sg13g2_dlygate4sd3_1
Xfanout1705 net1709 net1705 VPWR VGND sg13g2_buf_8
Xfanout1738 net1741 net1738 VPWR VGND sg13g2_buf_8
Xfanout1716 net1717 net1716 VPWR VGND sg13g2_buf_8
Xfanout1727 net1728 net1727 VPWR VGND sg13g2_buf_8
Xfanout1749 net1750 net1749 VPWR VGND sg13g2_buf_8
XFILLER_19_805 VPWR VGND sg13g2_fill_2
XFILLER_19_816 VPWR VGND sg13g2_fill_2
XFILLER_45_189 VPWR VGND sg13g2_fill_2
XFILLER_14_532 VPWR VGND sg13g2_fill_1
XFILLER_26_370 VPWR VGND sg13g2_fill_1
X_7722__301 VPWR VGND net301 sg13g2_tiehi
X_4050_ VPWR _3426_ net489 VGND sg13g2_inv_1
XFILLER_37_613 VPWR VGND sg13g2_fill_2
XFILLER_36_123 VPWR VGND sg13g2_fill_1
X_7740_ net281 VGND VPWR _0218_ s0.valid_out\[18\][0] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_4952_ _0950_ net1479 net591 VPWR VGND sg13g2_nand2_1
XFILLER_18_882 VPWR VGND sg13g2_fill_1
X_4883_ _0892_ _0891_ net1498 VPWR VGND sg13g2_nand2b_1
X_7671_ net356 VGND VPWR _0149_ s0.data_out\[24\]\[0\] clknet_leaf_4_clk sg13g2_dfrbpq_2
XFILLER_17_392 VPWR VGND sg13g2_fill_1
XFILLER_32_340 VPWR VGND sg13g2_fill_1
X_6622_ net1709 _2449_ _2456_ VPWR VGND sg13g2_nor2_1
X_7842__171 VPWR VGND net171 sg13g2_tiehi
XFILLER_9_580 VPWR VGND sg13g2_fill_1
X_6553_ net1305 VPWR _2398_ VGND _2335_ _2397_ sg13g2_o21ai_1
X_5504_ _1453_ net1433 net457 VPWR VGND sg13g2_nand2_1
X_6484_ _2328_ net1295 _2329_ _2330_ VPWR VGND sg13g2_a21o_1
X_5435_ net1624 _1330_ _1388_ VPWR VGND sg13g2_nor2_1
X_7912__96 VPWR VGND net96 sg13g2_tiehi
XFILLER_0_929 VPWR VGND sg13g2_decap_8
X_5366_ net1441 net1331 _1327_ VPWR VGND sg13g2_nor2b_1
X_4317_ VGND VPWR net1633 net1540 _0377_ _0375_ sg13g2_a21oi_1
X_5297_ net1462 VPWR _1265_ VGND _1235_ _1264_ sg13g2_o21ai_1
X_7105_ s0.data_out\[4\]\[0\] s0.data_out\[3\]\[0\] net1246 _2891_ VPWR VGND sg13g2_mux2_1
X_4248_ VGND VPWR net1558 _3611_ _3612_ _3607_ sg13g2_a21oi_1
X_7036_ net1688 _2799_ _2834_ VPWR VGND sg13g2_nor2_1
XFILLER_16_808 VPWR VGND sg13g2_fill_1
X_4179_ s0.data_out\[27\]\[5\] net1166 _3550_ VPWR VGND sg13g2_nor2_1
XFILLER_27_112 VPWR VGND sg13g2_fill_2
X_7938_ net68 VGND VPWR net422 s0.was_valid_out\[2\][0] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_7869_ net142 VGND VPWR _0003_ s0.shift_out\[8\][0] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_7706__318 VPWR VGND net318 sg13g2_tiehi
XFILLER_24_896 VPWR VGND sg13g2_fill_1
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_3_756 VPWR VGND sg13g2_decap_8
Xfanout1524 net1527 net1524 VPWR VGND sg13g2_buf_8
Xfanout1502 net424 net1502 VPWR VGND sg13g2_buf_1
Xfanout1513 net1514 net1513 VPWR VGND sg13g2_buf_8
Xfanout1557 s0.valid_out\[26\][0] net1557 VPWR VGND sg13g2_buf_8
Xfanout1546 net1548 net1546 VPWR VGND sg13g2_buf_8
Xfanout1535 net1536 net1535 VPWR VGND sg13g2_buf_8
Xfanout1579 net1580 net1579 VPWR VGND sg13g2_buf_8
Xfanout1568 net1569 net1568 VPWR VGND sg13g2_buf_8
XFILLER_47_955 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_487 VPWR VGND sg13g2_fill_1
XFILLER_33_159 VPWR VGND sg13g2_fill_2
X_7826__188 VPWR VGND net188 sg13g2_tiehi
XFILLER_14_351 VPWR VGND sg13g2_fill_2
XFILLER_41_192 VPWR VGND sg13g2_decap_4
X_7796__221 VPWR VGND net221 sg13g2_tiehi
XFILLER_6_561 VPWR VGND sg13g2_fill_1
X_5220_ net1447 net1358 _1193_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_1020 VPWR VGND sg13g2_decap_8
X_5151_ _1117_ _1132_ _1134_ _1135_ _1136_ VPWR VGND sg13g2_nor4_1
X_5082_ net1723 net397 _0195_ VPWR VGND sg13g2_and2_1
X_4102_ VPWR _3478_ s0.data_out\[14\]\[4\] VGND sg13g2_inv_1
X_4033_ _3409_ net452 VPWR VGND sg13g2_inv_2
X_7723_ net300 VGND VPWR _0201_ s0.data_out\[20\]\[4\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_5984_ _1883_ net1385 _1884_ _1885_ VPWR VGND sg13g2_a21o_1
X_4935_ _0179_ _0935_ _0936_ _3438_ net1604 VPWR VGND sg13g2_a22oi_1
X_7654_ net31 VGND VPWR _0132_ s0.data_out\[26\]\[7\] clknet_leaf_44_clk sg13g2_dfrbpq_2
X_4866_ s0.data_out\[22\]\[6\] s0.data_out\[21\]\[6\] net1490 _0875_ VPWR VGND sg13g2_mux2_1
X_7585_ VGND VPWR _3402_ _3319_ _3323_ _3322_ sg13g2_a21oi_1
X_4797_ _0812_ VPWR _0813_ VGND net1727 net764 sg13g2_o21ai_1
X_6605_ _2439_ net554 net1301 VPWR VGND sg13g2_nand2b_1
X_6536_ _2382_ net1309 _2381_ VPWR VGND sg13g2_nand2b_1
XFILLER_21_59 VPWR VGND sg13g2_fill_1
X_6467_ s0.was_valid_out\[8\][0] net1316 _2316_ VPWR VGND sg13g2_nor2_1
X_5418_ net1618 _1314_ _1375_ VPWR VGND sg13g2_nor2_1
X_6398_ s0.data_out\[10\]\[4\] s0.data_out\[9\]\[4\] net1314 _2256_ VPWR VGND sg13g2_mux2_1
XFILLER_0_726 VPWR VGND sg13g2_decap_8
X_5349_ s0.data_out\[18\]\[3\] s0.data_out\[17\]\[3\] net1446 _1310_ VPWR VGND sg13g2_mux2_1
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_34 VPWR VGND sg13g2_fill_1
X_7019_ VGND VPWR _2817_ _2815_ net1660 sg13g2_or2_1
XFILLER_29_933 VPWR VGND sg13g2_fill_1
XFILLER_44_925 VPWR VGND sg13g2_decap_8
XFILLER_29_999 VPWR VGND sg13g2_decap_8
XFILLER_15_115 VPWR VGND sg13g2_decap_4
XFILLER_43_468 VPWR VGND sg13g2_fill_1
XFILLER_12_822 VPWR VGND sg13g2_fill_1
XFILLER_8_848 VPWR VGND sg13g2_fill_2
Xfanout1332 s0.data_new_delayed\[7\] net1332 VPWR VGND sg13g2_buf_8
Xfanout1310 net1313 net1310 VPWR VGND sg13g2_buf_1
Xfanout1321 net1322 net1321 VPWR VGND sg13g2_buf_2
Xfanout1343 net1344 net1343 VPWR VGND sg13g2_buf_8
Xfanout1354 net1355 net1354 VPWR VGND sg13g2_buf_8
Xfanout1365 net1366 net1365 VPWR VGND sg13g2_buf_8
Xfanout1398 net825 net1398 VPWR VGND sg13g2_buf_8
XFILLER_4_1011 VPWR VGND sg13g2_decap_8
Xfanout1376 net1377 net1376 VPWR VGND sg13g2_buf_2
Xfanout1387 net1388 net1387 VPWR VGND sg13g2_buf_8
XFILLER_47_752 VPWR VGND sg13g2_decap_8
XFILLER_35_936 VPWR VGND sg13g2_fill_1
XFILLER_35_969 VPWR VGND sg13g2_decap_8
XFILLER_43_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_41_clk clknet_3_1__leaf_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
X_4720_ net1705 _0724_ _0741_ VPWR VGND sg13g2_nor2_1
X_4651_ VGND VPWR _0684_ net1566 net374 sg13g2_or2_1
XFILLER_30_696 VPWR VGND sg13g2_fill_2
X_7370_ net1221 net1167 _3132_ VPWR VGND sg13g2_nor2_1
X_4582_ _0613_ net1510 _0614_ _0615_ VPWR VGND sg13g2_a21o_1
X_6321_ _2187_ _2188_ _2189_ VPWR VGND sg13g2_nor2_1
X_6252_ _2127_ net1326 _2128_ _2129_ VPWR VGND sg13g2_a21o_1
X_6183_ VPWR _0297_ _2066_ VGND sg13g2_inv_1
X_5203_ net1744 net392 _0207_ VPWR VGND sg13g2_and2_1
X_5134_ _1118_ VPWR _1119_ VGND net1464 _3447_ sg13g2_o21ai_1
X_5065_ net1468 s0.data_out\[20\]\[7\] _1055_ VPWR VGND sg13g2_and2_1
XFILLER_38_752 VPWR VGND sg13g2_fill_2
X_4016_ _3392_ net1480 VPWR VGND sg13g2_inv_2
X_7949__55 VPWR VGND net55 sg13g2_tiehi
X_5967_ VGND VPWR net1378 _1866_ _1868_ _1867_ sg13g2_a21oi_1
Xclkbuf_leaf_32_clk clknet_3_5__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
X_4918_ _3391_ _3443_ _0923_ VPWR VGND sg13g2_nor2_1
X_7706_ net318 VGND VPWR _0184_ s0.data_out\[21\]\[0\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_34_991 VPWR VGND sg13g2_decap_8
X_5898_ _1811_ net1675 _1810_ VPWR VGND sg13g2_nand2_1
X_7637_ net49 VGND VPWR net633 s0.data_out\[27\]\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_4849_ net1486 net1168 _0858_ VPWR VGND sg13g2_nor2_1
XFILLER_20_151 VPWR VGND sg13g2_fill_1
XFILLER_20_184 VPWR VGND sg13g2_decap_4
X_7568_ _3310_ VPWR _3311_ VGND net1720 net737 sg13g2_o21ai_1
X_7499_ _3247_ net1223 _3248_ _3249_ VPWR VGND sg13g2_a21o_1
X_6519_ _2365_ _2364_ net1667 _2357_ net1657 VPWR VGND sg13g2_a22oi_1
XFILLER_0_534 VPWR VGND sg13g2_fill_2
XFILLER_48_538 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_23_clk clknet_3_7__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_8_612 VPWR VGND sg13g2_fill_2
XFILLER_40_983 VPWR VGND sg13g2_decap_8
X_7793__224 VPWR VGND net224 sg13g2_tiehi
XFILLER_26_1012 VPWR VGND sg13g2_decap_8
XFILLER_39_549 VPWR VGND sg13g2_fill_1
Xfanout1173 _3397_ net1173 VPWR VGND sg13g2_buf_8
Xfanout1184 net1186 net1184 VPWR VGND sg13g2_buf_8
Xfanout1195 _3381_ net1195 VPWR VGND sg13g2_buf_8
XFILLER_19_262 VPWR VGND sg13g2_fill_1
X_6870_ _2678_ net1262 _2679_ _2680_ VPWR VGND sg13g2_a21o_1
XFILLER_35_755 VPWR VGND sg13g2_fill_1
X_5821_ net1406 VPWR _1737_ VGND net1645 net1394 sg13g2_o21ai_1
X_5752_ _1677_ _1676_ net1665 _1669_ net1655 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_14_clk clknet_3_3__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_4703_ VGND VPWR net1513 _0721_ _0724_ _0723_ sg13g2_a21oi_1
XFILLER_33_1016 VPWR VGND sg13g2_decap_8
X_5683_ net1430 VPWR _1613_ VGND _1559_ _1612_ sg13g2_o21ai_1
XFILLER_33_1027 VPWR VGND sg13g2_fill_2
X_4634_ VGND VPWR net1524 _0664_ _0667_ _0666_ sg13g2_a21oi_1
X_7422_ VGND VPWR net1187 _3117_ _3182_ net1582 sg13g2_a21oi_1
X_4565_ net1580 _0535_ _0602_ VPWR VGND sg13g2_nor2_1
X_7353_ VGND VPWR net1217 _3113_ _3115_ _3114_ sg13g2_a21oi_1
X_6304_ net1612 _2142_ _2176_ VPWR VGND sg13g2_nor2_1
X_4496_ _0541_ net489 net1542 VPWR VGND sg13g2_nand2b_1
X_7284_ VGND VPWR net1243 _3055_ _3058_ _3057_ sg13g2_a21oi_1
X_6235_ net1322 net1168 _2112_ VPWR VGND sg13g2_nor2_1
X_6166_ VPWR _0293_ _2053_ VGND sg13g2_inv_1
X_5117_ net1460 net1336 _1102_ VPWR VGND sg13g2_nor2b_1
X_6097_ _1986_ s0.data_out\[11\]\[1\] net1386 VPWR VGND sg13g2_nand2b_1
XFILLER_45_519 VPWR VGND sg13g2_fill_2
X_5048_ net1488 VPWR _1042_ VGND _0976_ _1041_ sg13g2_o21ai_1
XFILLER_26_700 VPWR VGND sg13g2_decap_4
XFILLER_41_714 VPWR VGND sg13g2_fill_1
X_7937__69 VPWR VGND net69 sg13g2_tiehi
XFILLER_13_427 VPWR VGND sg13g2_fill_1
X_6999_ _2797_ net505 net1267 VPWR VGND sg13g2_nand2b_1
XFILLER_40_279 VPWR VGND sg13g2_fill_2
XFILLER_22_994 VPWR VGND sg13g2_decap_8
XFILLER_4_29 VPWR VGND sg13g2_fill_2
XFILLER_1_810 VPWR VGND sg13g2_decap_8
XFILLER_1_887 VPWR VGND sg13g2_decap_8
XFILLER_49_836 VPWR VGND sg13g2_decap_8
XFILLER_16_287 VPWR VGND sg13g2_fill_1
X_7901__108 VPWR VGND net108 sg13g2_tiehi
X_4350_ _0392_ VPWR _0407_ VGND net1701 _0399_ sg13g2_o21ai_1
X_4281_ VGND VPWR _0350_ net1565 net380 sg13g2_or2_1
X_6020_ _1919_ net1383 _1920_ _1921_ VPWR VGND sg13g2_a21o_1
Xclkbuf_leaf_3_clk clknet_3_0__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_7971_ net80 VGND VPWR _0105_ s0.data_out\[0\]\[5\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_6922_ VGND VPWR _2732_ net1566 net386 sg13g2_or2_1
X_6853_ net1262 net1357 _2663_ VPWR VGND sg13g2_nor2b_1
X_5804_ _1723_ VPWR _1724_ VGND net1196 _1722_ sg13g2_o21ai_1
X_6784_ s0.data_out\[6\]\[5\] s0.data_out\[7\]\[5\] net1291 _2606_ VPWR VGND sg13g2_mux2_1
X_3996_ VPWR _3372_ net524 VGND sg13g2_inv_1
X_5735_ _1641_ _1650_ _1651_ _1659_ _1660_ VPWR VGND sg13g2_nor4_1
X_5666_ net1197 _3474_ _1600_ VPWR VGND sg13g2_nor2_1
XFILLER_30_290 VPWR VGND sg13g2_fill_2
X_7405_ _3167_ s0.data_out\[1\]\[4\] net1238 VPWR VGND sg13g2_nand2b_1
X_4617_ VGND VPWR net1523 _0647_ _0650_ _0649_ sg13g2_a21oi_1
X_5597_ s0.data_out\[16\]\[0\] s0.data_out\[15\]\[0\] net1419 _1534_ VPWR VGND sg13g2_mux2_1
Xhold420 s0.data_out\[12\]\[2\] VPWR VGND net789 sg13g2_dlygate4sd3_1
Xhold431 _3288_ VPWR VGND net800 sg13g2_dlygate4sd3_1
X_4548_ VGND VPWR net1520 net698 _0588_ _0557_ sg13g2_a21oi_1
Xhold442 _0164_ VPWR VGND net811 sg13g2_dlygate4sd3_1
Xhold453 s0.data_new_delayed\[2\] VPWR VGND net822 sg13g2_dlygate4sd3_1
X_7336_ _3098_ VPWR _3101_ VGND s0.was_valid_out\[1\][0] net1224 sg13g2_o21ai_1
Xhold464 _2303_ VPWR VGND net833 sg13g2_dlygate4sd3_1
X_4479_ VGND VPWR _0408_ _0523_ _0524_ net1535 sg13g2_a21oi_1
X_7267_ VGND VPWR _3028_ _3030_ _3041_ net1659 sg13g2_a21oi_1
X_6218_ _2095_ net1360 net589 VPWR VGND sg13g2_nand2_1
X_7198_ net1244 s0.data_out\[3\]\[6\] _2977_ VPWR VGND sg13g2_and2_1
XFILLER_46_806 VPWR VGND sg13g2_decap_8
X_6149_ _1892_ VPWR _2038_ VGND net1388 _3497_ sg13g2_o21ai_1
XFILLER_9_206 VPWR VGND sg13g2_fill_1
XFILLER_6_913 VPWR VGND sg13g2_decap_8
XFILLER_10_997 VPWR VGND sg13g2_decap_8
X_7790__227 VPWR VGND net227 sg13g2_tiehi
XFILLER_49_633 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_fill_2
XFILLER_0_150 VPWR VGND sg13g2_decap_4
XFILLER_1_695 VPWR VGND sg13g2_decap_8
XFILLER_23_1026 VPWR VGND sg13g2_fill_2
XFILLER_45_872 VPWR VGND sg13g2_decap_8
X_5520_ _1469_ _1460_ _1468_ VPWR VGND sg13g2_nand2_1
X_7924__83 VPWR VGND net83 sg13g2_tiehi
XFILLER_8_283 VPWR VGND sg13g2_decap_4
X_5451_ _1399_ VPWR _1400_ VGND net1432 _3465_ sg13g2_o21ai_1
X_4402_ net370 net1565 _0458_ _0124_ VPWR VGND sg13g2_nor3_1
X_5382_ _1343_ net1445 s0.data_out\[17\]\[5\] VPWR VGND sg13g2_nand2_1
X_4333_ VGND VPWR _3564_ _0389_ _0390_ net1547 sg13g2_a21oi_1
X_7121_ _2907_ net1686 _2906_ VPWR VGND sg13g2_nand2_1
X_4264_ net1559 _3626_ _3627_ _3628_ VPWR VGND sg13g2_nor3_1
X_7052_ net1260 VPWR _2848_ VGND _2780_ _2847_ sg13g2_o21ai_1
X_6003_ _1904_ s0.data_out\[12\]\[5\] net1399 VPWR VGND sg13g2_nand2b_1
XFILLER_39_132 VPWR VGND sg13g2_fill_1
X_4195_ VGND VPWR _3557_ _3560_ _0109_ _3561_ sg13g2_a21oi_1
XFILLER_28_828 VPWR VGND sg13g2_fill_1
X_7954_ net321 VGND VPWR _0088_ s0.data_out\[1\]\[0\] clknet_leaf_9_clk sg13g2_dfrbpq_2
XFILLER_27_327 VPWR VGND sg13g2_fill_1
X_6905_ net1265 net1344 _2715_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_533 VPWR VGND sg13g2_fill_1
X_7885_ net125 VGND VPWR net594 s0.data_out\[7\]\[3\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_35_360 VPWR VGND sg13g2_fill_2
X_6836_ _2647_ VPWR _2649_ VGND s0.was_valid_out\[5\][0] net1268 sg13g2_o21ai_1
XFILLER_35_393 VPWR VGND sg13g2_fill_1
X_6767_ _2589_ _2588_ net1661 _2581_ net1651 VPWR VGND sg13g2_a22oi_1
XFILLER_11_739 VPWR VGND sg13g2_fill_1
X_5718_ _1642_ VPWR _1643_ VGND net1408 _3474_ sg13g2_o21ai_1
X_6698_ net1600 net427 _2526_ VPWR VGND sg13g2_nor2_1
X_5649_ _1583_ _1584_ _1585_ _1586_ VPWR VGND sg13g2_nor3_1
Xhold261 s0.data_out\[6\]\[7\] VPWR VGND net630 sg13g2_dlygate4sd3_1
XFILLER_3_949 VPWR VGND sg13g2_decap_8
Xhold250 s0.data_out\[23\]\[2\] VPWR VGND net619 sg13g2_dlygate4sd3_1
X_7319_ net1243 VPWR _3087_ VGND _3044_ _3086_ sg13g2_o21ai_1
Xhold294 s0.was_valid_out\[14\][0] VPWR VGND net663 sg13g2_dlygate4sd3_1
Xhold283 _0193_ VPWR VGND net652 sg13g2_dlygate4sd3_1
XFILLER_2_459 VPWR VGND sg13g2_decap_4
Xfanout1706 net1708 net1706 VPWR VGND sg13g2_buf_8
Xhold272 s0.data_out\[7\]\[0\] VPWR VGND net641 sg13g2_dlygate4sd3_1
Xfanout1739 net1740 net1739 VPWR VGND sg13g2_buf_8
Xfanout1717 net1733 net1717 VPWR VGND sg13g2_buf_2
Xfanout1728 net1733 net1728 VPWR VGND sg13g2_buf_8
XFILLER_18_327 VPWR VGND sg13g2_fill_1
XFILLER_14_555 VPWR VGND sg13g2_fill_1
X_7921__86 VPWR VGND net86 sg13g2_tiehi
XFILLER_1_492 VPWR VGND sg13g2_fill_2
XFILLER_36_146 VPWR VGND sg13g2_fill_2
X_4951_ net1606 _0942_ _0943_ _0182_ VPWR VGND sg13g2_nor3_1
X_4882_ _0771_ VPWR _0891_ VGND net1505 _3442_ sg13g2_o21ai_1
X_7670_ net357 VGND VPWR _0148_ s0.shift_out\[24\][0] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_6621_ _2455_ _2454_ net1293 VPWR VGND sg13g2_nand2b_1
X_6552_ net1295 s0.data_out\[8\]\[0\] _2397_ VPWR VGND sg13g2_and2_1
X_5503_ _1450_ _1448_ _1452_ VPWR VGND _1449_ sg13g2_nand3b_1
X_6483_ net1295 net1355 _2329_ VPWR VGND sg13g2_nor2b_1
X_5434_ net1451 VPWR _1387_ VGND _1327_ _1386_ sg13g2_o21ai_1
XFILLER_0_908 VPWR VGND sg13g2_decap_8
X_5365_ s0.data_out\[18\]\[7\] s0.data_out\[17\]\[7\] net1444 _1326_ VPWR VGND sg13g2_mux2_1
X_7104_ _2887_ _2889_ net1701 _2890_ VPWR VGND sg13g2_nand3_1
X_4316_ _0376_ net1633 net1542 VPWR VGND sg13g2_nand2_1
X_5296_ net1204 _3459_ _1264_ VPWR VGND sg13g2_nor2_1
X_4247_ _3609_ net1544 _3610_ _3611_ VPWR VGND sg13g2_a21o_1
X_7035_ _2833_ _2832_ net1670 _2825_ net1680 VPWR VGND sg13g2_a22oi_1
X_7630__204 VPWR VGND net204 sg13g2_tiehi
X_4178_ VGND VPWR _3406_ net1166 net7 _3549_ sg13g2_a21oi_1
XFILLER_19_48 VPWR VGND sg13g2_fill_2
XFILLER_42_105 VPWR VGND sg13g2_fill_2
XFILLER_15_319 VPWR VGND sg13g2_fill_2
X_7937_ net69 VGND VPWR net605 s0.data_out\[3\]\[7\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_7868_ net143 VGND VPWR _0002_ s0.genblk1\[7\].modules.bubble clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
XFILLER_23_330 VPWR VGND sg13g2_fill_2
X_6819_ VGND VPWR net1276 s0.data_out\[6\]\[5\] _2635_ _2603_ sg13g2_a21oi_1
X_7799_ net218 VGND VPWR net417 s0.was_valid_out\[13\][0] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_7819__196 VPWR VGND net196 sg13g2_tiehi
Xfanout1514 s0.shift_out\[23\][0] net1514 VPWR VGND sg13g2_buf_1
Xfanout1503 net1507 net1503 VPWR VGND sg13g2_buf_8
Xfanout1536 net1539 net1536 VPWR VGND sg13g2_buf_2
Xfanout1525 net1527 net1525 VPWR VGND sg13g2_buf_8
Xfanout1547 net1548 net1547 VPWR VGND sg13g2_buf_1
Xfanout1558 net1562 net1558 VPWR VGND sg13g2_buf_8
Xfanout1569 _0349_ net1569 VPWR VGND sg13g2_buf_8
XFILLER_47_934 VPWR VGND sg13g2_decap_8
XFILLER_46_422 VPWR VGND sg13g2_fill_1
XFILLER_18_146 VPWR VGND sg13g2_fill_2
XFILLER_18_168 VPWR VGND sg13g2_fill_2
XFILLER_33_116 VPWR VGND sg13g2_decap_8
XFILLER_34_639 VPWR VGND sg13g2_fill_1
XFILLER_42_672 VPWR VGND sg13g2_fill_1
XFILLER_10_591 VPWR VGND sg13g2_fill_1
XFILLER_6_584 VPWR VGND sg13g2_fill_1
X_5150_ _1135_ net1683 _1124_ VPWR VGND sg13g2_xnor2_1
X_5081_ net1606 _1061_ _0194_ VPWR VGND sg13g2_nor2_1
X_4101_ VPWR _3477_ net726 VGND sg13g2_inv_1
X_4032_ VPWR _3408_ net469 VGND sg13g2_inv_1
XFILLER_24_105 VPWR VGND sg13g2_fill_1
X_5983_ net1385 net1169 _1884_ VPWR VGND sg13g2_nor2_1
X_4934_ net1604 _0879_ _0936_ VPWR VGND sg13g2_nor2_1
X_7722_ net301 VGND VPWR net665 s0.data_out\[20\]\[3\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_36_1014 VPWR VGND sg13g2_decap_8
X_4865_ _0874_ net1489 net718 VPWR VGND sg13g2_nand2_1
X_7653_ net32 VGND VPWR _0131_ s0.data_out\[26\]\[6\] clknet_leaf_44_clk sg13g2_dfrbpq_2
X_7584_ net1649 _3321_ _3322_ VPWR VGND sg13g2_nor2_1
X_4796_ _0811_ VPWR _0812_ VGND net1181 _0810_ sg13g2_o21ai_1
X_6604_ _2436_ net1282 _2437_ _2438_ VPWR VGND sg13g2_a21o_1
X_6535_ VGND VPWR net1298 _2380_ _2381_ _2378_ sg13g2_a21oi_1
X_6466_ net1299 _2308_ _2315_ VPWR VGND sg13g2_nor2_1
XFILLER_0_705 VPWR VGND sg13g2_decap_8
X_5417_ net1449 VPWR _1374_ VGND _1311_ _1373_ sg13g2_o21ai_1
X_6397_ _2255_ net1314 s0.data_out\[9\]\[4\] VPWR VGND sg13g2_nand2_1
X_5348_ _1309_ net1446 net542 VPWR VGND sg13g2_nand2_1
X_7712__312 VPWR VGND net312 sg13g2_tiehi
X_5279_ VGND VPWR net1447 s0.data_out\[18\]\[0\] _1251_ _1193_ sg13g2_a21oi_1
X_7018_ _2816_ _2815_ net1660 _2808_ net1650 VPWR VGND sg13g2_a22oi_1
XFILLER_29_912 VPWR VGND sg13g2_fill_1
XFILLER_44_904 VPWR VGND sg13g2_decap_8
XFILLER_29_978 VPWR VGND sg13g2_decap_8
XFILLER_28_499 VPWR VGND sg13g2_fill_2
XFILLER_12_812 VPWR VGND sg13g2_fill_2
XFILLER_23_193 VPWR VGND sg13g2_fill_1
XFILLER_3_510 VPWR VGND sg13g2_fill_1
Xfanout1300 s0.shift_out\[8\][0] net1300 VPWR VGND sg13g2_buf_2
Xfanout1311 net1312 net1311 VPWR VGND sg13g2_buf_2
Xfanout1322 net1327 net1322 VPWR VGND sg13g2_buf_1
Xfanout1344 net829 net1344 VPWR VGND sg13g2_buf_8
Xfanout1333 net1334 net1333 VPWR VGND sg13g2_buf_8
Xfanout1355 s0.data_new_delayed\[1\] net1355 VPWR VGND sg13g2_buf_8
Xfanout1366 net1367 net1366 VPWR VGND sg13g2_buf_8
XFILLER_47_731 VPWR VGND sg13g2_decap_8
Xfanout1399 net1400 net1399 VPWR VGND sg13g2_buf_8
X_7832__182 VPWR VGND net182 sg13g2_tiehi
Xfanout1377 net1381 net1377 VPWR VGND sg13g2_buf_1
Xfanout1388 net1389 net1388 VPWR VGND sg13g2_buf_8
XFILLER_34_414 VPWR VGND sg13g2_fill_2
XFILLER_43_970 VPWR VGND sg13g2_decap_8
X_4650_ _0606_ _0681_ _0682_ _0683_ VPWR VGND sg13g2_nor3_1
X_6320_ net1646 net1316 _2188_ VPWR VGND sg13g2_nor2b_1
X_4581_ net1510 net1349 _0614_ VPWR VGND sg13g2_nor2b_1
X_6251_ net1326 net1330 _2128_ VPWR VGND sg13g2_nor2b_1
X_6182_ _2065_ VPWR _2066_ VGND net1739 net418 sg13g2_o21ai_1
X_5202_ net1742 _1175_ _0206_ VPWR VGND sg13g2_and2_1
X_5133_ _1118_ net1464 net435 VPWR VGND sg13g2_nand2_1
XFILLER_35_0 VPWR VGND sg13g2_fill_2
XFILLER_38_731 VPWR VGND sg13g2_decap_8
X_5064_ VPWR _0190_ _1054_ VGND sg13g2_inv_1
X_4015_ VPWR _3391_ net1488 VGND sg13g2_inv_1
XFILLER_16_38 VPWR VGND sg13g2_fill_2
X_5966_ net1378 net1355 _1867_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_970 VPWR VGND sg13g2_decap_8
X_5897_ VGND VPWR net1406 _1807_ _1810_ _1809_ sg13g2_a21oi_1
X_7705_ net319 VGND VPWR _0183_ s0.shift_out\[21\][0] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_4917_ VPWR _0175_ _0922_ VGND sg13g2_inv_1
XFILLER_33_480 VPWR VGND sg13g2_fill_1
XFILLER_33_491 VPWR VGND sg13g2_fill_2
X_4848_ _0842_ VPWR _0857_ VGND net1705 _0849_ sg13g2_o21ai_1
X_7636_ net50 VGND VPWR net560 s0.data_out\[27\]\[1\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_7567_ _3309_ VPWR _3310_ VGND net1202 _3308_ sg13g2_o21ai_1
X_4779_ _0798_ VPWR _0799_ VGND net1728 net740 sg13g2_o21ai_1
X_7498_ net1223 _3244_ _3248_ VPWR VGND sg13g2_nor2_1
X_6518_ VGND VPWR net1310 _2361_ _2364_ _2363_ sg13g2_a21oi_1
X_6449_ _0329_ _2299_ _2300_ _3502_ net1610 VPWR VGND sg13g2_a22oi_1
X_7816__199 VPWR VGND net199 sg13g2_tiehi
XFILLER_28_241 VPWR VGND sg13g2_fill_1
X_7786__232 VPWR VGND net232 sg13g2_tiehi
XFILLER_44_767 VPWR VGND sg13g2_decap_4
XFILLER_44_734 VPWR VGND sg13g2_decap_4
XFILLER_25_981 VPWR VGND sg13g2_decap_8
XFILLER_40_962 VPWR VGND sg13g2_decap_8
XFILLER_8_646 VPWR VGND sg13g2_fill_1
XFILLER_22_70 VPWR VGND sg13g2_fill_2
XFILLER_4_830 VPWR VGND sg13g2_decap_4
XFILLER_4_885 VPWR VGND sg13g2_decap_8
Xfanout1174 _3396_ net1174 VPWR VGND sg13g2_buf_8
Xfanout1185 net1186 net1185 VPWR VGND sg13g2_buf_1
Xfanout1196 _3380_ net1196 VPWR VGND sg13g2_buf_8
XFILLER_47_572 VPWR VGND sg13g2_fill_2
X_7946__59 VPWR VGND net59 sg13g2_tiehi
X_5820_ _0264_ _1735_ _1736_ _3472_ net1630 VPWR VGND sg13g2_a22oi_1
XFILLER_35_778 VPWR VGND sg13g2_fill_1
XFILLER_16_981 VPWR VGND sg13g2_decap_8
X_5751_ VGND VPWR net1418 _1673_ _1676_ _1675_ sg13g2_a21oi_1
X_4702_ VGND VPWR _0620_ _0722_ _0723_ net1513 sg13g2_a21oi_1
X_5682_ net1416 s0.data_out\[15\]\[6\] _1612_ VPWR VGND sg13g2_and2_1
XFILLER_30_450 VPWR VGND sg13g2_fill_1
X_7421_ VGND VPWR net1217 s0.data_out\[1\]\[1\] _3181_ _3114_ sg13g2_a21oi_1
X_4633_ VGND VPWR _0558_ _0665_ _0666_ net1524 sg13g2_a21oi_1
X_4564_ net1537 VPWR _0601_ VGND _0532_ _0600_ sg13g2_o21ai_1
X_7352_ net1217 net1352 _3114_ VPWR VGND sg13g2_nor2b_1
X_6303_ net1366 VPWR _2175_ VGND _2139_ _2174_ sg13g2_o21ai_1
X_7283_ VGND VPWR _2921_ _3056_ _3057_ net1243 sg13g2_a21oi_1
X_4495_ _0538_ net1520 _0539_ _0540_ VPWR VGND sg13g2_a21o_1
X_6234_ _2110_ VPWR _2111_ VGND net1361 _3493_ sg13g2_o21ai_1
X_6165_ _2052_ VPWR _2053_ VGND net1740 net692 sg13g2_o21ai_1
X_5116_ s0.data_out\[20\]\[6\] s0.data_out\[19\]\[6\] net1464 _1101_ VPWR VGND sg13g2_mux2_1
X_6096_ _1984_ net1367 _1982_ _1985_ VPWR VGND sg13g2_a21o_1
X_5047_ net1471 s0.data_out\[20\]\[3\] _1041_ VPWR VGND sg13g2_and2_1
XFILLER_14_918 VPWR VGND sg13g2_fill_2
X_6998_ _2794_ net1252 _2795_ _2796_ VPWR VGND sg13g2_a21o_1
X_5949_ _1850_ VPWR _1853_ VGND s0.was_valid_out\[12\][0] net1389 sg13g2_o21ai_1
XFILLER_41_759 VPWR VGND sg13g2_fill_2
XFILLER_22_973 VPWR VGND sg13g2_decap_8
X_7619_ net1721 net459 _3354_ VPWR VGND sg13g2_nor2_1
XFILLER_4_159 VPWR VGND sg13g2_fill_1
XFILLER_49_815 VPWR VGND sg13g2_decap_8
XFILLER_1_866 VPWR VGND sg13g2_decap_8
XFILLER_17_712 VPWR VGND sg13g2_fill_2
XFILLER_16_200 VPWR VGND sg13g2_fill_1
XFILLER_17_734 VPWR VGND sg13g2_fill_1
XFILLER_44_597 VPWR VGND sg13g2_fill_1
X_7936__70 VPWR VGND net70 sg13g2_tiehi
XFILLER_8_410 VPWR VGND sg13g2_fill_2
XFILLER_12_472 VPWR VGND sg13g2_fill_2
XFILLER_13_984 VPWR VGND sg13g2_decap_8
XFILLER_9_988 VPWR VGND sg13g2_decap_8
X_4280_ _0349_ net1638 net1718 VPWR VGND sg13g2_nand2_1
X_7970_ net93 VGND VPWR _0104_ s0.data_out\[0\]\[4\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_6921_ VGND VPWR _2726_ _2729_ _2731_ _2730_ sg13g2_a21oi_1
X_6852_ _2662_ net1175 _2661_ VPWR VGND sg13g2_nand2_1
XFILLER_22_214 VPWR VGND sg13g2_fill_1
X_5803_ VGND VPWR net1196 _1695_ _1723_ net1630 sg13g2_a21oi_1
X_6783_ _2605_ net1285 _2604_ VPWR VGND sg13g2_nand2b_1
X_3995_ VPWR _3371_ net419 VGND sg13g2_inv_1
X_5734_ net1693 _1658_ _1659_ VPWR VGND sg13g2_nor2_1
X_5665_ _0246_ _1598_ _1599_ _3471_ net1620 VPWR VGND sg13g2_a22oi_1
X_7404_ _3164_ net1221 _3165_ _3166_ VPWR VGND sg13g2_a21o_1
X_4616_ VGND VPWR _0530_ _0648_ _0649_ net1523 sg13g2_a21oi_1
Xhold410 s0.data_out\[18\]\[0\] VPWR VGND net779 sg13g2_dlygate4sd3_1
X_5596_ net1706 _1532_ _1533_ VPWR VGND sg13g2_nor2_1
X_7776__242 VPWR VGND net242 sg13g2_tiehi
X_7335_ _3098_ _3099_ _3100_ VPWR VGND sg13g2_nor2_1
Xhold432 s0.data_out\[7\]\[6\] VPWR VGND net801 sg13g2_dlygate4sd3_1
X_4547_ _0140_ _0586_ _0587_ _3422_ net1579 VPWR VGND sg13g2_a22oi_1
Xhold454 s0.valid_out\[17\][0] VPWR VGND net823 sg13g2_dlygate4sd3_1
Xhold443 s0.data_out\[3\]\[6\] VPWR VGND net812 sg13g2_dlygate4sd3_1
Xhold421 _0295_ VPWR VGND net790 sg13g2_dlygate4sd3_1
Xhold465 s0.data_out\[25\]\[6\] VPWR VGND net834 sg13g2_dlygate4sd3_1
X_4478_ _0523_ net478 net1540 VPWR VGND sg13g2_nand2b_1
X_7266_ net1648 _3038_ _3040_ VPWR VGND sg13g2_nor2_1
X_6217_ VGND VPWR _2094_ _2093_ net1697 sg13g2_or2_1
X_7197_ VPWR _0057_ _2976_ VGND sg13g2_inv_1
X_6148_ _2037_ net1379 _2036_ VPWR VGND sg13g2_nand2b_1
X_6079_ s0.was_valid_out\[11\][0] net1387 _1971_ VPWR VGND sg13g2_nor2_1
X_7783__235 VPWR VGND net235 sg13g2_tiehi
XFILLER_16_1023 VPWR VGND sg13g2_decap_4
X_7933__73 VPWR VGND net73 sg13g2_tiehi
XFILLER_10_976 VPWR VGND sg13g2_decap_8
XFILLER_1_641 VPWR VGND sg13g2_decap_8
XFILLER_49_612 VPWR VGND sg13g2_decap_8
XFILLER_1_674 VPWR VGND sg13g2_decap_8
XFILLER_23_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_689 VPWR VGND sg13g2_decap_8
XFILLER_17_520 VPWR VGND sg13g2_decap_4
XFILLER_45_851 VPWR VGND sg13g2_decap_8
XFILLER_9_741 VPWR VGND sg13g2_fill_2
XFILLER_8_251 VPWR VGND sg13g2_decap_8
X_5450_ _1399_ net1432 net495 VPWR VGND sg13g2_nand2_1
X_4401_ VPWR VGND _0453_ _0457_ _0456_ _0416_ _0458_ _0455_ sg13g2_a221oi_1
X_5381_ VGND VPWR net1451 _1339_ _1342_ _1341_ sg13g2_a21oi_1
X_4332_ _0389_ s0.data_out\[25\]\[2\] net1557 VPWR VGND sg13g2_nand2b_1
X_7120_ VGND VPWR net1249 _2903_ _2906_ _2905_ sg13g2_a21oi_1
X_4263_ net1563 s0.data_out\[26\]\[4\] _3627_ VPWR VGND sg13g2_nor2_1
X_7051_ net1250 net716 _2847_ VPWR VGND sg13g2_and2_1
XFILLER_39_100 VPWR VGND sg13g2_decap_4
X_6002_ _1901_ net1382 _1902_ _1903_ VPWR VGND sg13g2_a21o_1
X_4194_ net1714 VPWR _3561_ VGND net676 _3556_ sg13g2_o21ai_1
XFILLER_28_818 VPWR VGND sg13g2_fill_1
X_7953_ net334 VGND VPWR _0087_ s0.shift_out\[1\][0] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_6904_ _2711_ _2713_ net1670 _2714_ VPWR VGND sg13g2_nand3_1
XFILLER_36_884 VPWR VGND sg13g2_fill_2
X_7884_ net126 VGND VPWR net555 s0.data_out\[7\]\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_6835_ VGND VPWR _3396_ _2534_ _2648_ _2647_ sg13g2_a21oi_1
X_6766_ VGND VPWR net1285 _2585_ _2588_ _2587_ sg13g2_a21oi_1
X_5717_ _1642_ net1408 net730 VPWR VGND sg13g2_nand2_1
X_6697_ net1296 VPWR _2525_ VGND _2492_ _2524_ sg13g2_o21ai_1
X_5648_ net1674 _1581_ _1585_ VPWR VGND sg13g2_nor2_1
X_7930__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_3_928 VPWR VGND sg13g2_decap_8
X_5579_ net1622 _1511_ _0242_ VPWR VGND sg13g2_nor2_1
Xhold240 _0010_ VPWR VGND net609 sg13g2_dlygate4sd3_1
Xhold262 _2644_ VPWR VGND net631 sg13g2_dlygate4sd3_1
Xhold251 _0806_ VPWR VGND net620 sg13g2_dlygate4sd3_1
X_7318_ net1233 s0.data_out\[2\]\[5\] _3086_ VPWR VGND sg13g2_and2_1
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_1016 VPWR VGND sg13g2_decap_8
Xhold284 s0.data_out\[7\]\[4\] VPWR VGND net653 sg13g2_dlygate4sd3_1
Xhold295 s0.data_out\[20\]\[3\] VPWR VGND net664 sg13g2_dlygate4sd3_1
Xhold273 _2621_ VPWR VGND net642 sg13g2_dlygate4sd3_1
X_7249_ _3022_ VPWR _3023_ VGND _3012_ _3014_ sg13g2_o21ai_1
Xfanout1729 net1730 net1729 VPWR VGND sg13g2_buf_8
Xfanout1718 net1719 net1718 VPWR VGND sg13g2_buf_8
Xfanout1707 net1708 net1707 VPWR VGND sg13g2_buf_8
XFILLER_42_865 VPWR VGND sg13g2_fill_2
XFILLER_6_788 VPWR VGND sg13g2_fill_2
XFILLER_2_994 VPWR VGND sg13g2_decap_8
XFILLER_49_464 VPWR VGND sg13g2_decap_4
XFILLER_37_648 VPWR VGND sg13g2_fill_1
X_4950_ VGND VPWR _3368_ _0944_ _0181_ _0949_ sg13g2_a21oi_1
X_4881_ _0890_ net1498 _0889_ VPWR VGND sg13g2_nand2b_1
X_6620_ s0.data_out\[7\]\[0\] s0.data_out\[8\]\[0\] net1301 _2454_ VPWR VGND sg13g2_mux2_1
XFILLER_32_375 VPWR VGND sg13g2_fill_1
X_6551_ VGND VPWR _2391_ _2395_ _0335_ _2396_ sg13g2_a21oi_1
X_5502_ VPWR _1451_ _1450_ VGND sg13g2_inv_1
X_6482_ s0.data_out\[9\]\[1\] s0.data_out\[8\]\[1\] net1302 _2328_ VPWR VGND sg13g2_mux2_1
X_7957__282 VPWR VGND net282 sg13g2_tiehi
X_5433_ net1207 _3462_ _1386_ VPWR VGND sg13g2_nor2_1
X_5364_ _1325_ net1444 net585 VPWR VGND sg13g2_nand2_1
X_4315_ net1549 VPWR _0375_ VGND net1639 net1533 sg13g2_o21ai_1
X_7103_ _2889_ net1170 _2888_ VPWR VGND sg13g2_nand2_1
X_5295_ _0212_ _1262_ _1263_ _3454_ net1617 VPWR VGND sg13g2_a22oi_1
X_4246_ net1544 net1333 _3610_ VPWR VGND sg13g2_nor2b_1
X_7034_ VGND VPWR net1263 _2829_ _2832_ _2831_ sg13g2_a21oi_1
X_4177_ s0.data_out\[27\]\[4\] net1166 _3549_ VPWR VGND sg13g2_nor2_1
XFILLER_42_117 VPWR VGND sg13g2_decap_8
X_7936_ net70 VGND VPWR _0070_ s0.data_out\[3\]\[6\] clknet_leaf_2_clk sg13g2_dfrbpq_2
X_7867_ net144 VGND VPWR _0001_ s0.valid_out\[8\][0] clknet_leaf_15_clk sg13g2_dfrbpq_2
XFILLER_11_504 VPWR VGND sg13g2_decap_4
XFILLER_23_353 VPWR VGND sg13g2_fill_1
X_7780__238 VPWR VGND net238 sg13g2_tiehi
X_6818_ VPWR _0020_ net654 VGND sg13g2_inv_1
X_7798_ net219 VGND VPWR _0276_ s0.data_out\[14\]\[7\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_6749_ VGND VPWR _2459_ _2570_ _2571_ net1284 sg13g2_a21oi_1
XFILLER_13_1026 VPWR VGND sg13g2_fill_2
XFILLER_3_714 VPWR VGND sg13g2_fill_1
Xfanout1515 net1518 net1515 VPWR VGND sg13g2_buf_8
Xfanout1504 net1507 net1504 VPWR VGND sg13g2_buf_1
Xfanout1537 net1538 net1537 VPWR VGND sg13g2_buf_8
Xfanout1548 s0.shift_out\[26\][0] net1548 VPWR VGND sg13g2_buf_2
Xfanout1526 net1527 net1526 VPWR VGND sg13g2_buf_1
XFILLER_47_913 VPWR VGND sg13g2_decap_8
Xfanout1559 net1562 net1559 VPWR VGND sg13g2_buf_1
XFILLER_19_604 VPWR VGND sg13g2_fill_2
XFILLER_18_114 VPWR VGND sg13g2_fill_2
XFILLER_20_1019 VPWR VGND sg13g2_decap_8
XFILLER_46_478 VPWR VGND sg13g2_fill_2
XFILLER_27_670 VPWR VGND sg13g2_fill_2
XFILLER_14_375 VPWR VGND sg13g2_fill_2
XFILLER_37_4 VPWR VGND sg13g2_fill_2
X_5080_ VGND VPWR _1063_ _1066_ _0193_ _1067_ sg13g2_a21oi_1
XFILLER_2_791 VPWR VGND sg13g2_decap_8
X_4100_ VPWR _3476_ net819 VGND sg13g2_inv_1
X_4031_ VPWR _3407_ net517 VGND sg13g2_inv_1
XFILLER_38_979 VPWR VGND sg13g2_decap_8
X_5982_ _1882_ VPWR _1883_ VGND net1389 _3485_ sg13g2_o21ai_1
X_4933_ net1499 VPWR _0935_ VGND _0876_ _0934_ sg13g2_o21ai_1
X_7721_ net302 VGND VPWR net592 s0.data_out\[20\]\[2\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_7652_ net33 VGND VPWR net492 s0.data_out\[26\]\[5\] clknet_leaf_0_clk sg13g2_dfrbpq_2
X_4864_ VGND VPWR net1498 _0870_ _0873_ _0872_ sg13g2_a21oi_1
X_7583_ _3320_ VPWR _3321_ VGND _3393_ net1329 sg13g2_o21ai_1
X_4795_ VGND VPWR net1181 _0783_ _0811_ net1594 sg13g2_a21oi_1
X_6603_ net1282 net1349 _2437_ VPWR VGND sg13g2_nor2b_1
X_6534_ s0.data_out\[9\]\[4\] s0.data_out\[8\]\[4\] net1302 _2380_ VPWR VGND sg13g2_mux2_1
X_6465_ _2310_ VPWR _2314_ VGND s0.was_valid_out\[8\][0] net1304 sg13g2_o21ai_1
X_5416_ net1206 _3463_ _1373_ VPWR VGND sg13g2_nor2_1
X_6396_ _2253_ _2251_ _2254_ VPWR VGND _2252_ sg13g2_nand3b_1
X_5347_ VPWR VGND _1306_ _1307_ _1299_ net1573 _1308_ _1291_ sg13g2_a221oi_1
XFILLER_43_1019 VPWR VGND sg13g2_decap_8
X_5278_ net372 net1568 _1250_ _0208_ VPWR VGND sg13g2_nor3_1
X_4229_ _3591_ net1547 _3592_ _3593_ VPWR VGND sg13g2_a21o_1
X_7017_ VGND VPWR net1258 _2812_ _2815_ _2814_ sg13g2_a21oi_1
XFILLER_28_445 VPWR VGND sg13g2_decap_8
XFILLER_43_448 VPWR VGND sg13g2_fill_1
X_7919_ net88 VGND VPWR _0053_ s0.data_out\[4\]\[1\] clknet_leaf_4_clk sg13g2_dfrbpq_2
XFILLER_24_673 VPWR VGND sg13g2_fill_1
XFILLER_12_835 VPWR VGND sg13g2_fill_2
XFILLER_7_338 VPWR VGND sg13g2_decap_4
Xfanout1323 net1324 net1323 VPWR VGND sg13g2_buf_8
Xfanout1312 net1313 net1312 VPWR VGND sg13g2_buf_2
Xfanout1301 s0.valid_out\[8\][0] net1301 VPWR VGND sg13g2_buf_8
Xfanout1334 net1337 net1334 VPWR VGND sg13g2_buf_8
Xfanout1356 net1357 net1356 VPWR VGND sg13g2_buf_8
Xfanout1345 net1346 net1345 VPWR VGND sg13g2_buf_8
XFILLER_47_710 VPWR VGND sg13g2_decap_8
Xfanout1389 s0.valid_out\[12\][0] net1389 VPWR VGND sg13g2_buf_8
XFILLER_16_9 VPWR VGND sg13g2_fill_2
Xfanout1378 net1381 net1378 VPWR VGND sg13g2_buf_2
Xfanout1367 s0.shift_out\[11\][0] net1367 VPWR VGND sg13g2_buf_8
XFILLER_47_787 VPWR VGND sg13g2_decap_8
XFILLER_42_492 VPWR VGND sg13g2_fill_2
X_4580_ s0.data_out\[24\]\[2\] s0.data_out\[23\]\[2\] net1515 _0613_ VPWR VGND sg13g2_mux2_1
XFILLER_7_872 VPWR VGND sg13g2_decap_4
X_6250_ s0.data_out\[11\]\[7\] s0.data_out\[10\]\[7\] net1363 _2127_ VPWR VGND sg13g2_mux2_1
X_6181_ _2039_ _2064_ net1739 _2065_ VPWR VGND sg13g2_nand3_1
X_5201_ VGND VPWR _3367_ _1175_ _0205_ _1176_ sg13g2_a21oi_1
X_5132_ _1116_ _1114_ _1117_ VPWR VGND _1115_ sg13g2_nand3b_1
X_5063_ _1053_ VPWR _1054_ VGND net1736 net718 sg13g2_o21ai_1
X_4014_ VPWR _3390_ net1513 VGND sg13g2_inv_1
XFILLER_26_905 VPWR VGND sg13g2_fill_1
X_5965_ s0.data_out\[13\]\[1\] s0.data_out\[12\]\[1\] net1386 _1866_ VPWR VGND sg13g2_mux2_1
X_5896_ VGND VPWR _1682_ _1808_ _1809_ net1406 sg13g2_a21oi_1
X_7704_ net320 VGND VPWR _0182_ s0.valid_out\[21\][0] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_4916_ _0921_ VPWR _0922_ VGND net1735 net711 sg13g2_o21ai_1
X_7635_ net51 VGND VPWR net573 s0.data_out\[27\]\[0\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_4847_ VPWR VGND _0855_ net1711 _0853_ net1705 _0856_ _0849_ sg13g2_a221oi_1
X_7566_ VGND VPWR net1202 _3250_ _3309_ net1583 sg13g2_a21oi_1
X_4778_ _0797_ VPWR _0798_ VGND net1182 _0796_ sg13g2_o21ai_1
X_7497_ VGND VPWR net1212 _3245_ _3247_ _3246_ sg13g2_a21oi_1
X_6517_ VGND VPWR _2244_ _2362_ _2363_ net1309 sg13g2_a21oi_1
XFILLER_10_1018 VPWR VGND sg13g2_decap_8
X_6448_ net1610 _2268_ _2300_ VPWR VGND sg13g2_nor2_1
X_6379_ _2237_ net1316 net483 VPWR VGND sg13g2_nand2_1
XFILLER_0_536 VPWR VGND sg13g2_fill_1
XFILLER_0_569 VPWR VGND sg13g2_fill_2
XFILLER_48_529 VPWR VGND sg13g2_decap_8
X_7966__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_29_732 VPWR VGND sg13g2_decap_4
XFILLER_19_1021 VPWR VGND sg13g2_decap_8
XFILLER_40_941 VPWR VGND sg13g2_decap_8
XFILLER_4_820 VPWR VGND sg13g2_decap_4
XFILLER_39_507 VPWR VGND sg13g2_decap_4
Xfanout1175 _3396_ net1175 VPWR VGND sg13g2_buf_8
Xfanout1186 _3388_ net1186 VPWR VGND sg13g2_buf_8
Xfanout1197 _3380_ net1197 VPWR VGND sg13g2_buf_8
XFILLER_47_551 VPWR VGND sg13g2_fill_2
XFILLER_34_267 VPWR VGND sg13g2_fill_1
XFILLER_15_481 VPWR VGND sg13g2_fill_2
X_5750_ VGND VPWR _1557_ _1674_ _1675_ net1417 sg13g2_a21oi_1
X_4701_ _0722_ net599 net1517 VPWR VGND sg13g2_nand2b_1
X_5681_ _0250_ _1610_ _1611_ _3467_ net1623 VPWR VGND sg13g2_a22oi_1
X_4632_ _0665_ s0.data_out\[23\]\[4\] net1530 VPWR VGND sg13g2_nand2b_1
X_7420_ VPWR _0076_ net722 VGND sg13g2_inv_1
XFILLER_31_985 VPWR VGND sg13g2_decap_8
X_7702__323 VPWR VGND net323 sg13g2_tiehi
X_4563_ net1520 net525 _0600_ VPWR VGND sg13g2_and2_1
X_7351_ s0.data_out\[2\]\[1\] s0.data_out\[1\]\[1\] net1224 _3113_ VPWR VGND sg13g2_mux2_1
X_4494_ net1520 net1333 _0539_ VPWR VGND sg13g2_nor2b_1
X_7282_ _3056_ net520 s0.valid_out\[3\][0] VPWR VGND sg13g2_nand2b_1
X_6302_ net1322 net747 _2174_ VPWR VGND sg13g2_and2_1
X_6233_ _2110_ net1361 net443 VPWR VGND sg13g2_nand2_1
X_6164_ _1994_ _2051_ net1740 _2052_ VPWR VGND sg13g2_nand3_1
X_5115_ _1100_ net1466 net645 VPWR VGND sg13g2_nand2_1
X_6095_ _1983_ VPWR _1984_ VGND net1373 _3491_ sg13g2_o21ai_1
X_5046_ VPWR _0186_ net512 VGND sg13g2_inv_1
X_6997_ net1252 net1167 _2795_ VPWR VGND sg13g2_nor2_1
X_5948_ _1850_ _1851_ _1852_ VPWR VGND sg13g2_nor2_1
X_7945__60 VPWR VGND net60 sg13g2_tiehi
X_5879_ _1792_ _1791_ net1665 _1784_ net1656 VPWR VGND sg13g2_a22oi_1
X_7618_ VGND VPWR net1720 _3329_ _0101_ _3353_ sg13g2_a21oi_1
X_7549_ VPWR _0090_ net660 VGND sg13g2_inv_1
X_7822__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_49_1025 VPWR VGND sg13g2_decap_4
XFILLER_0_311 VPWR VGND sg13g2_fill_1
XFILLER_1_845 VPWR VGND sg13g2_decap_8
XFILLER_1_1027 VPWR VGND sg13g2_fill_2
XFILLER_9_967 VPWR VGND sg13g2_decap_8
XFILLER_8_488 VPWR VGND sg13g2_fill_1
XFILLER_48_893 VPWR VGND sg13g2_decap_8
X_6920_ _2648_ VPWR _2730_ VGND _2703_ _2705_ sg13g2_o21ai_1
X_7769__250 VPWR VGND net250 sg13g2_tiehi
X_6851_ s0.data_out\[5\]\[0\] s0.data_out\[6\]\[0\] net1278 _2661_ VPWR VGND sg13g2_mux2_1
X_5802_ VGND VPWR net1404 net588 _1722_ _1690_ sg13g2_a21oi_1
X_6782_ VGND VPWR net1276 _2602_ _2604_ _2603_ sg13g2_a21oi_1
X_3994_ VPWR _3370_ net409 VGND sg13g2_inv_1
X_5733_ VGND VPWR net1414 _1655_ _1658_ _1657_ sg13g2_a21oi_1
X_5664_ net1620 _1531_ _1599_ VPWR VGND sg13g2_nor2_1
X_7942__63 VPWR VGND net63 sg13g2_tiehi
X_7403_ net1221 net1344 _3165_ VPWR VGND sg13g2_nor2b_1
X_4615_ _0648_ s0.data_out\[23\]\[7\] net1530 VPWR VGND sg13g2_nand2b_1
X_5595_ VGND VPWR net1425 _1529_ _1532_ _1531_ sg13g2_a21oi_1
XFILLER_30_292 VPWR VGND sg13g2_fill_1
X_4546_ net1579 _0524_ _0587_ VPWR VGND sg13g2_nor2_1
X_7334_ net1229 _2984_ _3099_ VPWR VGND sg13g2_nor2_1
Xhold411 s0.data_out\[4\]\[7\] VPWR VGND net780 sg13g2_dlygate4sd3_1
Xhold400 s0.data_out\[1\]\[1\] VPWR VGND net769 sg13g2_dlygate4sd3_1
Xhold422 s0.data_out\[16\]\[4\] VPWR VGND net791 sg13g2_dlygate4sd3_1
Xhold444 s0.data_out\[17\]\[1\] VPWR VGND net813 sg13g2_dlygate4sd3_1
Xhold433 s0.data_out\[7\]\[1\] VPWR VGND net802 sg13g2_dlygate4sd3_1
Xhold466 s0.data_out\[20\]\[6\] VPWR VGND net835 sg13g2_dlygate4sd3_1
X_4477_ _0520_ net1521 _0521_ _0522_ VPWR VGND sg13g2_a21o_1
Xhold455 s0.valid_out\[3\][0] VPWR VGND net824 sg13g2_dlygate4sd3_1
X_7265_ _3039_ _3038_ net1648 _3031_ net1659 VPWR VGND sg13g2_a22oi_1
X_6216_ VGND VPWR net1365 _2090_ _2093_ _2092_ sg13g2_a21oi_1
X_7196_ _2975_ VPWR _2976_ VGND net1723 net793 sg13g2_o21ai_1
X_6147_ VGND VPWR net1370 _2034_ _2036_ _2035_ sg13g2_a21oi_1
XFILLER_38_59 VPWR VGND sg13g2_fill_1
X_6078_ net1370 _1963_ _1970_ VPWR VGND sg13g2_nor2_1
X_5029_ _0942_ _0943_ _1025_ _1026_ _1027_ VPWR VGND sg13g2_nor4_1
XFILLER_41_524 VPWR VGND sg13g2_decap_8
XFILLER_13_226 VPWR VGND sg13g2_fill_2
XFILLER_16_1002 VPWR VGND sg13g2_decap_8
XFILLER_22_760 VPWR VGND sg13g2_fill_1
XFILLER_6_959 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_668 VPWR VGND sg13g2_decap_8
XFILLER_45_830 VPWR VGND sg13g2_decap_8
XFILLER_44_340 VPWR VGND sg13g2_fill_1
XFILLER_32_535 VPWR VGND sg13g2_fill_2
XFILLER_9_731 VPWR VGND sg13g2_decap_4
XFILLER_9_775 VPWR VGND sg13g2_fill_2
XFILLER_8_296 VPWR VGND sg13g2_fill_2
X_4400_ _0379_ VPWR _0457_ VGND _0431_ _0433_ sg13g2_o21ai_1
X_5380_ VGND VPWR _1236_ _1340_ _1341_ net1450 sg13g2_a21oi_1
X_4331_ _0386_ net1535 _0387_ _0388_ VPWR VGND sg13g2_a21o_1
XFILLER_4_480 VPWR VGND sg13g2_fill_2
X_4262_ net469 net1563 _3626_ VPWR VGND sg13g2_nor2b_1
X_7050_ VPWR _0040_ _2846_ VGND sg13g2_inv_1
X_6001_ net1382 net1341 _1902_ VPWR VGND sg13g2_nor2b_1
X_4193_ _3558_ _3559_ _3560_ VPWR VGND sg13g2_nor2_1
XFILLER_48_690 VPWR VGND sg13g2_decap_8
X_7952_ net347 VGND VPWR _0086_ s0.genblk1\[19\].modules.bubble clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_6903_ _2713_ net1174 _2712_ VPWR VGND sg13g2_nand2_1
XFILLER_39_1013 VPWR VGND sg13g2_decap_8
XFILLER_23_524 VPWR VGND sg13g2_fill_1
X_7883_ net127 VGND VPWR net803 s0.data_out\[7\]\[1\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_6834_ VGND VPWR net1634 net1268 _2647_ _2646_ sg13g2_a21oi_1
X_6765_ VGND VPWR _2467_ _2586_ _2587_ net1285 sg13g2_a21oi_1
XFILLER_10_207 VPWR VGND sg13g2_fill_1
X_5716_ VPWR VGND _1640_ net1712 _1636_ net1707 _1641_ _1634_ sg13g2_a221oi_1
X_6696_ net1286 net712 _2524_ VPWR VGND sg13g2_and2_1
X_5647_ net1683 _1574_ _1584_ VPWR VGND sg13g2_nor2_1
XFILLER_3_907 VPWR VGND sg13g2_decap_8
X_5578_ VGND VPWR _1513_ _1516_ _0241_ _1517_ sg13g2_a21oi_1
X_7317_ _0068_ _3084_ _3085_ _3537_ net1585 VPWR VGND sg13g2_a22oi_1
Xhold241 s0.data_out\[23\]\[5\] VPWR VGND net610 sg13g2_dlygate4sd3_1
XFILLER_2_428 VPWR VGND sg13g2_fill_2
X_4529_ VGND VPWR _0574_ net1565 net379 sg13g2_or2_1
Xhold230 s0.data_out\[22\]\[1\] VPWR VGND net599 sg13g2_dlygate4sd3_1
Xhold252 s0.data_out\[26\]\[1\] VPWR VGND net621 sg13g2_dlygate4sd3_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
Xhold285 _2634_ VPWR VGND net654 sg13g2_dlygate4sd3_1
Xhold296 _0200_ VPWR VGND net665 sg13g2_dlygate4sd3_1
Xhold263 s0.data_out\[27\]\[2\] VPWR VGND net632 sg13g2_dlygate4sd3_1
X_7248_ _3022_ _3021_ net1686 _3011_ net1696 VPWR VGND sg13g2_a22oi_1
Xhold274 s0.data_out\[6\]\[0\] VPWR VGND net643 sg13g2_dlygate4sd3_1
Xfanout1719 net1724 net1719 VPWR VGND sg13g2_buf_2
Xfanout1708 net1709 net1708 VPWR VGND sg13g2_buf_8
X_7179_ VGND VPWR net1240 s0.data_out\[3\]\[2\] _2962_ _2879_ sg13g2_a21oi_1
XFILLER_46_638 VPWR VGND sg13g2_fill_2
XFILLER_27_852 VPWR VGND sg13g2_fill_2
XFILLER_26_351 VPWR VGND sg13g2_fill_1
XFILLER_42_844 VPWR VGND sg13g2_fill_2
XFILLER_41_343 VPWR VGND sg13g2_decap_4
XFILLER_2_973 VPWR VGND sg13g2_decap_8
XFILLER_49_432 VPWR VGND sg13g2_fill_2
XFILLER_7_1011 VPWR VGND sg13g2_decap_8
XFILLER_1_494 VPWR VGND sg13g2_fill_1
X_7766__253 VPWR VGND net253 sg13g2_tiehi
X_4880_ VGND VPWR net1485 _0887_ _0889_ _0888_ sg13g2_a21oi_1
XFILLER_33_899 VPWR VGND sg13g2_fill_2
X_6550_ VGND VPWR _2396_ net1567 net394 sg13g2_or2_1
X_5501_ VGND VPWR _1450_ _1440_ net1654 sg13g2_or2_1
X_6481_ _2327_ net1301 net649 VPWR VGND sg13g2_nand2_1
X_5432_ VPWR _0227_ net768 VGND sg13g2_inv_1
X_5363_ VGND VPWR net1451 _1321_ _1324_ _1323_ sg13g2_a21oi_1
X_4314_ _0120_ _0373_ _0374_ _3399_ net1575 VPWR VGND sg13g2_a22oi_1
X_7102_ s0.data_out\[3\]\[1\] s0.data_out\[4\]\[1\] net1253 _2888_ VPWR VGND sg13g2_mux2_1
X_7773__246 VPWR VGND net246 sg13g2_tiehi
X_5294_ net1617 _1205_ _1263_ VPWR VGND sg13g2_nor2_1
X_4245_ s0.data_out\[27\]\[6\] s0.data_out\[26\]\[6\] net1554 _3609_ VPWR VGND sg13g2_mux2_1
X_7033_ VGND VPWR _2707_ _2830_ _2831_ net1263 sg13g2_a21oi_1
X_4176_ _3548_ VPWR net6 VGND _3410_ net1165 sg13g2_o21ai_1
XFILLER_28_627 VPWR VGND sg13g2_fill_2
XFILLER_42_107 VPWR VGND sg13g2_fill_1
X_7935_ net71 VGND VPWR net504 s0.data_out\[3\]\[5\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_7866_ net146 VGND VPWR net749 s0.was_valid_out\[8\][0] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_24_833 VPWR VGND sg13g2_fill_1
XFILLER_35_192 VPWR VGND sg13g2_fill_1
X_6817_ _2633_ VPWR _2634_ VGND net1731 net653 sg13g2_o21ai_1
X_7797_ net220 VGND VPWR _0275_ s0.data_out\[14\]\[6\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_7_509 VPWR VGND sg13g2_decap_8
XFILLER_13_1005 VPWR VGND sg13g2_decap_8
X_6748_ _2570_ s0.data_out\[6\]\[3\] net1290 VPWR VGND sg13g2_nand2b_1
X_6679_ VPWR _0004_ _2511_ VGND sg13g2_inv_1
XFILLER_2_247 VPWR VGND sg13g2_fill_1
Xfanout1505 net1507 net1505 VPWR VGND sg13g2_buf_2
Xfanout1516 net1518 net1516 VPWR VGND sg13g2_buf_8
Xfanout1538 net1539 net1538 VPWR VGND sg13g2_buf_8
Xfanout1527 s0.shift_out\[24\][0] net1527 VPWR VGND sg13g2_buf_8
Xfanout1549 net1553 net1549 VPWR VGND sg13g2_buf_8
XFILLER_19_649 VPWR VGND sg13g2_fill_1
XFILLER_47_969 VPWR VGND sg13g2_decap_8
XFILLER_18_148 VPWR VGND sg13g2_fill_1
XFILLER_2_770 VPWR VGND sg13g2_decap_8
X_4030_ _3406_ net1677 VPWR VGND sg13g2_inv_8
XFILLER_38_958 VPWR VGND sg13g2_decap_8
X_5981_ _1882_ net1388 net597 VPWR VGND sg13g2_nand2_1
X_4932_ net1482 s0.data_out\[21\]\[6\] _0934_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_44_clk clknet_3_0__leaf_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
X_7720_ net303 VGND VPWR net498 s0.data_out\[20\]\[1\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_7651_ net34 VGND VPWR _0129_ s0.data_out\[26\]\[4\] clknet_leaf_44_clk sg13g2_dfrbpq_2
X_4863_ VGND VPWR _0753_ _0871_ _0872_ net1498 sg13g2_a21oi_1
X_6602_ s0.data_out\[8\]\[2\] s0.data_out\[7\]\[2\] net1289 _2436_ VPWR VGND sg13g2_mux2_1
X_7582_ net447 net1215 net1210 _3320_ VPWR VGND sg13g2_a21o_1
X_4794_ VGND VPWR net1494 net411 _0810_ _0779_ sg13g2_a21oi_1
X_6533_ _2379_ net1301 net818 VPWR VGND sg13g2_nand2_1
X_6464_ net455 _2312_ _2313_ VPWR VGND sg13g2_nor2_1
X_5415_ VPWR _0223_ _1372_ VGND sg13g2_inv_1
X_6395_ VGND VPWR _2253_ _2243_ net1653 sg13g2_or2_1
X_5346_ VGND VPWR _1296_ _1298_ _1307_ net1708 sg13g2_a21oi_1
X_5277_ VPWR VGND _1245_ _1249_ _1248_ _1208_ _1250_ _1247_ sg13g2_a221oi_1
X_4228_ net1551 net1167 _3592_ VPWR VGND sg13g2_nor2_1
X_7016_ VGND VPWR _2689_ _2813_ _2814_ net1258 sg13g2_a21oi_1
X_4159_ VPWR _3535_ net604 VGND sg13g2_inv_1
XFILLER_44_939 VPWR VGND sg13g2_decap_8
X_7918_ net89 VGND VPWR _0052_ s0.data_out\[4\]\[0\] clknet_leaf_3_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_35_clk clknet_3_4__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
X_7849_ net164 VGND VPWR net546 s0.data_out\[10\]\[3\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_7_328 VPWR VGND sg13g2_fill_2
XFILLER_11_368 VPWR VGND sg13g2_fill_2
XFILLER_20_880 VPWR VGND sg13g2_fill_1
Xfanout1313 net704 net1313 VPWR VGND sg13g2_buf_8
Xfanout1302 s0.valid_out\[8\][0] net1302 VPWR VGND sg13g2_buf_2
Xfanout1335 net1337 net1335 VPWR VGND sg13g2_buf_8
Xfanout1324 net1327 net1324 VPWR VGND sg13g2_buf_2
Xfanout1346 s0.data_new_delayed\[4\] net1346 VPWR VGND sg13g2_buf_8
Xfanout1357 net830 net1357 VPWR VGND sg13g2_buf_8
Xfanout1368 net1371 net1368 VPWR VGND sg13g2_buf_8
Xfanout1379 net1380 net1379 VPWR VGND sg13g2_buf_8
XFILLER_4_1025 VPWR VGND sg13g2_decap_4
XFILLER_47_766 VPWR VGND sg13g2_decap_8
XFILLER_19_479 VPWR VGND sg13g2_fill_1
XFILLER_34_416 VPWR VGND sg13g2_fill_1
XFILLER_15_630 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_26_clk clknet_3_6__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_30_600 VPWR VGND sg13g2_fill_1
XFILLER_7_884 VPWR VGND sg13g2_fill_2
X_6180_ net1379 VPWR _2064_ VGND _2035_ _2063_ sg13g2_o21ai_1
X_5200_ net1742 VPWR _1176_ VGND _1172_ _1174_ sg13g2_o21ai_1
X_5131_ VGND VPWR _1116_ _1113_ net1654 sg13g2_or2_1
XFILLER_35_2 VPWR VGND sg13g2_fill_1
X_5062_ _1052_ net1736 _1053_ VPWR VGND _0996_ sg13g2_nand3b_1
X_7770__249 VPWR VGND net249 sg13g2_tiehi
X_4013_ _3389_ net1531 VPWR VGND sg13g2_inv_2
X_7703_ net322 VGND VPWR net413 s0.was_valid_out\[21\][0] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_5964_ _1865_ net1386 net513 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_17_clk clknet_3_6__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
X_5895_ _1808_ net582 net1411 VPWR VGND sg13g2_nand2b_1
X_4915_ _0840_ _0920_ net1734 _0921_ VPWR VGND sg13g2_nand3_1
X_7634_ net52 VGND VPWR _0112_ s0.shift_out\[27\][0] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4846_ _0855_ _0854_ net1501 VPWR VGND sg13g2_nand2b_1
X_7565_ VGND VPWR net1209 net404 _3308_ _3252_ sg13g2_a21oi_1
X_6516_ _2362_ net608 net1316 VPWR VGND sg13g2_nand2b_1
X_4777_ VGND VPWR net1182 _0725_ _0797_ net1595 sg13g2_a21oi_1
X_7496_ net1210 net1329 _3246_ VPWR VGND sg13g2_nor2b_1
X_6447_ net1324 VPWR _2299_ VGND _2265_ _2298_ sg13g2_o21ai_1
X_6378_ _2235_ VPWR _2236_ VGND _2226_ _2227_ sg13g2_o21ai_1
X_5329_ _1290_ net1204 _1289_ VPWR VGND sg13g2_nand2_1
XFILLER_44_758 VPWR VGND sg13g2_fill_1
XFILLER_16_438 VPWR VGND sg13g2_decap_8
XFILLER_16_449 VPWR VGND sg13g2_fill_1
XFILLER_19_1000 VPWR VGND sg13g2_decap_8
XFILLER_40_997 VPWR VGND sg13g2_decap_8
XFILLER_7_136 VPWR VGND sg13g2_fill_1
XFILLER_22_72 VPWR VGND sg13g2_fill_1
XFILLER_26_1026 VPWR VGND sg13g2_fill_2
Xfanout1165 _3544_ net1165 VPWR VGND sg13g2_buf_8
Xfanout1176 net1177 net1176 VPWR VGND sg13g2_buf_8
Xfanout1198 net1199 net1198 VPWR VGND sg13g2_buf_8
Xfanout1187 net1189 net1187 VPWR VGND sg13g2_buf_8
XFILLER_47_574 VPWR VGND sg13g2_fill_1
X_4700_ _0719_ net1495 _0720_ _0721_ VPWR VGND sg13g2_a21o_1
X_5680_ net1623 net458 _1611_ VPWR VGND sg13g2_nor2_1
X_4631_ _0662_ net1508 _0663_ _0664_ VPWR VGND sg13g2_a21o_1
X_4562_ VPWR _0143_ net776 VGND sg13g2_inv_1
X_7350_ _3112_ net1224 net769 VPWR VGND sg13g2_nand2_1
X_4493_ s0.data_out\[25\]\[6\] s0.data_out\[24\]\[6\] net1528 _0538_ VPWR VGND sg13g2_mux2_1
X_6301_ _0308_ _2172_ _2173_ _3493_ net1611 VPWR VGND sg13g2_a22oi_1
X_7281_ _3053_ net1232 _3054_ _3055_ VPWR VGND sg13g2_a21o_1
X_6232_ _2094_ VPWR _2109_ VGND net1707 _2101_ sg13g2_o21ai_1
Xclkbuf_leaf_6_clk clknet_3_3__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
X_6163_ net1376 VPWR _2051_ VGND _1990_ _2050_ sg13g2_o21ai_1
X_5114_ _1098_ VPWR _1099_ VGND _1089_ _1090_ sg13g2_o21ai_1
X_6094_ _1983_ net1372 net675 VPWR VGND sg13g2_nand2_1
X_5045_ _1039_ VPWR _1040_ VGND net1734 net511 sg13g2_o21ai_1
XFILLER_25_213 VPWR VGND sg13g2_fill_2
X_6996_ _2793_ VPWR _2794_ VGND net1256 _3528_ sg13g2_o21ai_1
X_5947_ VGND VPWR net1635 net1398 _1851_ net1393 sg13g2_a21oi_1
XFILLER_34_780 VPWR VGND sg13g2_fill_1
XFILLER_22_931 VPWR VGND sg13g2_fill_1
X_7617_ net1720 net430 _3353_ VPWR VGND sg13g2_nor2_1
X_5878_ VGND VPWR net1406 _1788_ _1791_ _1790_ sg13g2_a21oi_1
X_4829_ _0838_ net1500 _0837_ VPWR VGND sg13g2_nand2b_1
X_7548_ _3294_ VPWR _3295_ VGND net1721 net659 sg13g2_o21ai_1
XFILLER_49_1004 VPWR VGND sg13g2_decap_8
X_7479_ s0.data_out\[1\]\[0\] s0.data_out\[0\]\[0\] net1214 _3229_ VPWR VGND sg13g2_mux2_1
XFILLER_4_139 VPWR VGND sg13g2_fill_2
XFILLER_1_824 VPWR VGND sg13g2_decap_8
XFILLER_1_1006 VPWR VGND sg13g2_decap_8
XFILLER_17_714 VPWR VGND sg13g2_fill_1
XFILLER_44_544 VPWR VGND sg13g2_fill_1
XFILLER_17_83 VPWR VGND sg13g2_decap_4
XFILLER_12_474 VPWR VGND sg13g2_fill_1
XFILLER_39_316 VPWR VGND sg13g2_fill_2
Xhold1 s0.genblk1\[26\].modules.bubble VPWR VGND net370 sg13g2_dlygate4sd3_1
XFILLER_48_872 VPWR VGND sg13g2_decap_8
XFILLER_47_360 VPWR VGND sg13g2_fill_2
X_6850_ VGND VPWR net1270 _2657_ _2660_ _2659_ sg13g2_a21oi_1
X_6781_ net1276 net1342 _2603_ VPWR VGND sg13g2_nor2b_1
X_5801_ _0260_ _1720_ _1721_ _3473_ net1630 VPWR VGND sg13g2_a22oi_1
X_3993_ VPWR _3369_ net425 VGND sg13g2_inv_1
X_5732_ VGND VPWR _1542_ _1656_ _1657_ net1414 sg13g2_a21oi_1
X_5663_ net1424 VPWR _1598_ VGND _1528_ _1597_ sg13g2_o21ai_1
X_7402_ s0.data_out\[2\]\[4\] s0.data_out\[1\]\[4\] net1226 _3164_ VPWR VGND sg13g2_mux2_1
X_4614_ _0645_ net1509 _0646_ _0647_ VPWR VGND sg13g2_a21o_1
X_5594_ VGND VPWR _1399_ _1530_ _1531_ net1424 sg13g2_a21oi_1
X_4545_ net1538 VPWR _0586_ VGND _0521_ _0585_ sg13g2_o21ai_1
Xhold401 s0.data_out\[3\]\[1\] VPWR VGND net770 sg13g2_dlygate4sd3_1
X_7333_ _3096_ _3097_ _3098_ VPWR VGND sg13g2_nor2_1
Xhold445 s0.data_out\[19\]\[3\] VPWR VGND net814 sg13g2_dlygate4sd3_1
Xhold423 s0.data_out\[17\]\[5\] VPWR VGND net792 sg13g2_dlygate4sd3_1
Xhold412 s0.data_out\[4\]\[0\] VPWR VGND net781 sg13g2_dlygate4sd3_1
Xhold434 _0017_ VPWR VGND net803 sg13g2_dlygate4sd3_1
Xhold456 s0.valid_out\[13\][0] VPWR VGND net825 sg13g2_dlygate4sd3_1
Xhold467 s0.data_out\[20\]\[6\] VPWR VGND net836 sg13g2_dlygate4sd3_1
X_4476_ net1521 net1167 _0521_ VPWR VGND sg13g2_nor2_1
X_7264_ VGND VPWR net1239 _3035_ _3038_ _3037_ sg13g2_a21oi_1
X_7195_ _2974_ VPWR _2975_ VGND net1172 _2973_ sg13g2_o21ai_1
X_6215_ VGND VPWR _1974_ _2091_ _2092_ net1365 sg13g2_a21oi_1
X_6146_ net1370 net1345 _2035_ VPWR VGND sg13g2_nor2b_1
X_6077_ _1965_ VPWR _1969_ VGND s0.was_valid_out\[11\][0] net1375 sg13g2_o21ai_1
XFILLER_39_872 VPWR VGND sg13g2_fill_1
X_5028_ _0998_ _1000_ _1026_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_577 VPWR VGND sg13g2_decap_4
XFILLER_41_547 VPWR VGND sg13g2_fill_2
XFILLER_41_536 VPWR VGND sg13g2_fill_1
X_6979_ VGND VPWR _2777_ _2776_ net1700 sg13g2_or2_1
XFILLER_22_783 VPWR VGND sg13g2_fill_1
XFILLER_6_927 VPWR VGND sg13g2_fill_1
XFILLER_6_938 VPWR VGND sg13g2_decap_8
XFILLER_1_621 VPWR VGND sg13g2_decap_8
XFILLER_49_647 VPWR VGND sg13g2_decap_8
XFILLER_48_146 VPWR VGND sg13g2_fill_1
XFILLER_17_511 VPWR VGND sg13g2_decap_4
XFILLER_45_886 VPWR VGND sg13g2_decap_8
XFILLER_40_591 VPWR VGND sg13g2_fill_2
X_4330_ net1535 net1348 _0387_ VPWR VGND sg13g2_nor2b_1
XFILLER_5_993 VPWR VGND sg13g2_decap_8
X_4261_ _3625_ net1668 _3624_ VPWR VGND sg13g2_nand2_1
XFILLER_5_75 VPWR VGND sg13g2_fill_1
X_6000_ s0.data_out\[13\]\[5\] s0.data_out\[12\]\[5\] net1389 _1901_ VPWR VGND sg13g2_mux2_1
X_4192_ VGND VPWR _3372_ _3385_ _3559_ net1560 sg13g2_a21oi_1
X_7951_ net360 VGND VPWR _0085_ s0.valid_out\[1\][0] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_36_820 VPWR VGND sg13g2_fill_1
X_6902_ _2601_ VPWR _2712_ VGND net1280 _3526_ sg13g2_o21ai_1
X_7882_ net128 VGND VPWR _0016_ s0.data_out\[7\]\[0\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_35_330 VPWR VGND sg13g2_fill_2
X_6833_ net1274 VPWR _2646_ VGND net1642 net1264 sg13g2_o21ai_1
X_6764_ _2586_ net719 net1291 VPWR VGND sg13g2_nand2b_1
X_6695_ _0008_ _2522_ _2523_ _3510_ net1600 VPWR VGND sg13g2_a22oi_1
X_5715_ _1640_ net1413 _1639_ VPWR VGND sg13g2_nand2b_1
X_5646_ net1692 _1548_ _1583_ VPWR VGND sg13g2_nor2_1
X_5577_ net1744 VPWR _1517_ VGND net636 _1511_ sg13g2_o21ai_1
Xhold220 s0.data_out\[10\]\[1\] VPWR VGND net589 sg13g2_dlygate4sd3_1
X_4528_ VGND VPWR _0567_ _0571_ _0573_ _0572_ sg13g2_a21oi_1
Xhold242 _0702_ VPWR VGND net611 sg13g2_dlygate4sd3_1
Xhold253 _0126_ VPWR VGND net622 sg13g2_dlygate4sd3_1
Xhold231 _0174_ VPWR VGND net600 sg13g2_dlygate4sd3_1
X_7316_ net1585 _3057_ _3085_ VPWR VGND sg13g2_nor2_1
Xhold264 _0115_ VPWR VGND net633 sg13g2_dlygate4sd3_1
X_4459_ _0504_ net1528 s0.data_out\[24\]\[0\] VPWR VGND sg13g2_nand2_1
Xhold286 s0.data_out\[16\]\[2\] VPWR VGND net655 sg13g2_dlygate4sd3_1
Xhold275 s0.data_out\[15\]\[5\] VPWR VGND net644 sg13g2_dlygate4sd3_1
X_7247_ VGND VPWR net1243 _3018_ _3021_ _3020_ sg13g2_a21oi_1
Xhold297 s0.data_out\[5\]\[5\] VPWR VGND net666 sg13g2_dlygate4sd3_1
Xfanout1709 ui_in[1] net1709 VPWR VGND sg13g2_buf_8
X_7178_ VPWR _0053_ net717 VGND sg13g2_inv_1
X_6129_ VGND VPWR _1918_ _2017_ _2018_ net1380 sg13g2_a21oi_1
XFILLER_41_366 VPWR VGND sg13g2_fill_1
X_7759__261 VPWR VGND net261 sg13g2_tiehi
XFILLER_2_952 VPWR VGND sg13g2_decap_8
XFILLER_49_411 VPWR VGND sg13g2_decap_4
XFILLER_18_831 VPWR VGND sg13g2_decap_4
X_5500_ net1664 _1447_ _1449_ VPWR VGND sg13g2_nor2_1
X_6480_ net1699 _2325_ _2326_ VPWR VGND sg13g2_nor2_1
X_5431_ _1384_ VPWR _1385_ VGND net1744 net767 sg13g2_o21ai_1
X_5362_ VGND VPWR _1209_ _1322_ _1323_ net1451 sg13g2_a21oi_1
X_4313_ net1575 _3599_ _0374_ VPWR VGND sg13g2_nor2_1
X_7101_ _2887_ net1248 _2886_ VPWR VGND sg13g2_nand2b_1
X_7032_ _2830_ s0.data_out\[4\]\[5\] net1268 VPWR VGND sg13g2_nand2b_1
X_5293_ net1463 VPWR _1262_ VGND _1202_ _1261_ sg13g2_o21ai_1
X_4244_ _3608_ net1556 s0.data_out\[26\]\[6\] VPWR VGND sg13g2_nand2_1
X_4175_ _3548_ net1687 net1165 VPWR VGND sg13g2_nand2_1
XFILLER_28_606 VPWR VGND sg13g2_fill_2
X_7934_ net72 VGND VPWR net617 s0.data_out\[3\]\[4\] clknet_leaf_9_clk sg13g2_dfrbpq_2
XFILLER_35_39 VPWR VGND sg13g2_fill_2
X_7865_ net147 VGND VPWR net484 s0.data_out\[9\]\[7\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_7796_ net221 VGND VPWR _0274_ s0.data_out\[14\]\[5\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_6816_ _2632_ VPWR _2633_ VGND net1176 _2631_ sg13g2_o21ai_1
X_6747_ _2567_ net1272 _2568_ _2569_ VPWR VGND sg13g2_a21o_1
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
X_6678_ _2510_ VPWR _2511_ VGND net1728 net806 sg13g2_o21ai_1
X_5629_ net1664 _1563_ _1566_ VPWR VGND sg13g2_nor2_1
Xfanout1506 net1507 net1506 VPWR VGND sg13g2_buf_1
Xfanout1517 net1518 net1517 VPWR VGND sg13g2_buf_2
Xfanout1539 net785 net1539 VPWR VGND sg13g2_buf_2
Xfanout1528 net1532 net1528 VPWR VGND sg13g2_buf_8
XFILLER_47_948 VPWR VGND sg13g2_decap_8
XFILLER_42_686 VPWR VGND sg13g2_fill_2
XFILLER_14_399 VPWR VGND sg13g2_fill_2
XFILLER_25_83 VPWR VGND sg13g2_fill_1
XFILLER_6_521 VPWR VGND sg13g2_fill_2
XFILLER_29_1013 VPWR VGND sg13g2_decap_8
XFILLER_37_436 VPWR VGND sg13g2_fill_1
XFILLER_46_981 VPWR VGND sg13g2_decap_8
XFILLER_25_609 VPWR VGND sg13g2_fill_2
X_5980_ VPWR VGND _1879_ _1880_ _1872_ net1574 _1881_ _1864_ sg13g2_a221oi_1
XFILLER_45_480 VPWR VGND sg13g2_fill_1
X_4931_ VPWR _0178_ _0933_ VGND sg13g2_inv_1
X_7650_ net35 VGND VPWR net502 s0.data_out\[26\]\[3\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_4862_ _0871_ net538 net1505 VPWR VGND sg13g2_nand2b_1
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
X_6601_ _2435_ net1289 net554 VPWR VGND sg13g2_nand2_1
XFILLER_32_163 VPWR VGND sg13g2_fill_2
X_7581_ VGND VPWR _3318_ _3319_ _3401_ net1209 sg13g2_a21oi_2
X_4793_ _0164_ _0808_ _0809_ _3434_ net1594 VPWR VGND sg13g2_a22oi_1
X_6532_ net1298 net1344 _2378_ VPWR VGND sg13g2_nor2b_1
X_6463_ _2311_ VPWR _2312_ VGND net1311 _2188_ sg13g2_o21ai_1
X_5414_ _1371_ VPWR _1372_ VGND net1743 net678 sg13g2_o21ai_1
X_6394_ net1663 _2250_ _2252_ VPWR VGND sg13g2_nor2_1
XFILLER_0_719 VPWR VGND sg13g2_decap_8
X_5345_ net1570 _1305_ _1306_ VPWR VGND sg13g2_and2_1
X_5276_ _1175_ VPWR _1249_ VGND _1223_ _1225_ sg13g2_o21ai_1
X_4227_ _3590_ VPWR _3591_ VGND net1555 _3410_ sg13g2_o21ai_1
X_7015_ _2813_ net536 net1267 VPWR VGND sg13g2_nand2b_1
XFILLER_28_414 VPWR VGND sg13g2_fill_2
X_4158_ VPWR _3534_ net794 VGND sg13g2_inv_1
XFILLER_44_918 VPWR VGND sg13g2_decap_8
X_4089_ VPWR _3465_ net813 VGND sg13g2_inv_1
XFILLER_15_119 VPWR VGND sg13g2_fill_1
X_7917_ net90 VGND VPWR _0051_ s0.shift_out\[4\][0] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_7848_ net165 VGND VPWR _0326_ s0.data_out\[10\]\[2\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_7779_ net239 VGND VPWR _0257_ s0.data_out\[15\]\[0\] clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_3_557 VPWR VGND sg13g2_fill_1
XFILLER_11_96 VPWR VGND sg13g2_fill_2
X_7756__264 VPWR VGND net264 sg13g2_tiehi
Xfanout1303 net1304 net1303 VPWR VGND sg13g2_buf_8
Xfanout1314 net1318 net1314 VPWR VGND sg13g2_buf_8
Xfanout1336 net1337 net1336 VPWR VGND sg13g2_buf_8
Xfanout1347 s0.data_new_delayed\[3\] net1347 VPWR VGND sg13g2_buf_8
Xfanout1325 net1327 net1325 VPWR VGND sg13g2_buf_2
Xfanout1369 net1371 net1369 VPWR VGND sg13g2_buf_1
XFILLER_4_1004 VPWR VGND sg13g2_decap_8
Xfanout1358 net1359 net1358 VPWR VGND sg13g2_buf_8
XFILLER_47_745 VPWR VGND sg13g2_decap_8
XFILLER_46_233 VPWR VGND sg13g2_fill_2
X_7973__29 VPWR VGND net29 sg13g2_tiehi
XFILLER_28_992 VPWR VGND sg13g2_decap_8
XFILLER_14_130 VPWR VGND sg13g2_fill_1
XFILLER_43_984 VPWR VGND sg13g2_decap_8
X_7763__257 VPWR VGND net257 sg13g2_tiehi
X_5130_ net1664 _1106_ _1115_ VPWR VGND sg13g2_nor2_1
XFILLER_42_1010 VPWR VGND sg13g2_decap_8
XFILLER_2_590 VPWR VGND sg13g2_decap_8
X_5061_ net1483 VPWR _1052_ VGND _0993_ _1051_ sg13g2_o21ai_1
X_4012_ VPWR _3388_ net1534 VGND sg13g2_inv_1
XFILLER_38_745 VPWR VGND sg13g2_decap_8
X_5963_ _1863_ VPWR _1864_ VGND net1193 _1861_ sg13g2_o21ai_1
X_7702_ net323 VGND VPWR _0180_ s0.data_out\[22\]\[7\] clknet_leaf_41_clk sg13g2_dfrbpq_2
X_4914_ net1501 VPWR _0920_ VGND _0836_ _0919_ sg13g2_o21ai_1
X_5894_ _1805_ net1394 _1806_ _1807_ VPWR VGND sg13g2_a21o_1
XFILLER_34_984 VPWR VGND sg13g2_decap_8
X_7633_ net53 VGND VPWR _0111_ s0.genblk1\[26\].modules.bubble clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
X_4845_ s0.data_out\[21\]\[0\] s0.data_out\[22\]\[0\] net1506 _0854_ VPWR VGND sg13g2_mux2_1
X_7564_ VPWR _0093_ net734 VGND sg13g2_inv_1
X_4776_ VGND VPWR net1496 s0.data_out\[22\]\[0\] _0796_ _0727_ sg13g2_a21oi_1
X_6515_ _2359_ net1298 _2360_ _2361_ VPWR VGND sg13g2_a21o_1
X_7495_ s0.data_out\[1\]\[7\] s0.data_out\[0\]\[7\] net1215 _3245_ VPWR VGND sg13g2_mux2_1
X_6446_ net1312 s0.data_out\[9\]\[5\] _2298_ VPWR VGND sg13g2_and2_1
X_6377_ _2235_ _2234_ net1691 _2211_ net1699 VPWR VGND sg13g2_a22oi_1
XFILLER_0_516 VPWR VGND sg13g2_decap_8
XFILLER_0_527 VPWR VGND sg13g2_decap_8
X_5328_ _1177_ VPWR _1289_ VGND net1454 _3464_ sg13g2_o21ai_1
X_5259_ _1125_ VPWR _1232_ VGND net1466 _3458_ sg13g2_o21ai_1
XFILLER_29_701 VPWR VGND sg13g2_decap_4
XFILLER_17_918 VPWR VGND sg13g2_fill_1
XFILLER_25_995 VPWR VGND sg13g2_decap_8
XFILLER_11_111 VPWR VGND sg13g2_fill_1
XFILLER_40_976 VPWR VGND sg13g2_decap_8
XFILLER_4_800 VPWR VGND sg13g2_decap_8
XFILLER_4_899 VPWR VGND sg13g2_decap_8
XFILLER_26_1005 VPWR VGND sg13g2_decap_8
Xfanout1177 _3395_ net1177 VPWR VGND sg13g2_buf_8
Xfanout1188 net1189 net1188 VPWR VGND sg13g2_buf_8
Xfanout1199 _3379_ net1199 VPWR VGND sg13g2_buf_8
Xfanout1166 _3544_ net1166 VPWR VGND sg13g2_buf_8
XFILLER_14_8 VPWR VGND sg13g2_decap_8
XFILLER_43_770 VPWR VGND sg13g2_fill_1
XFILLER_16_995 VPWR VGND sg13g2_decap_8
XFILLER_15_483 VPWR VGND sg13g2_fill_1
XFILLER_15_494 VPWR VGND sg13g2_decap_4
X_4630_ net1508 net1344 _0663_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_1009 VPWR VGND sg13g2_decap_8
XFILLER_30_486 VPWR VGND sg13g2_fill_2
X_4561_ _0598_ VPWR _0599_ VGND net1716 net775 sg13g2_o21ai_1
X_6300_ net1611 net444 _2173_ VPWR VGND sg13g2_nor2_1
X_7280_ net1232 net1344 _3054_ VPWR VGND sg13g2_nor2b_1
X_4492_ _0537_ net1530 net489 VPWR VGND sg13g2_nand2_1
X_6231_ VPWR VGND _2107_ net1711 _2105_ net1707 _2108_ _2101_ sg13g2_a221oi_1
X_6162_ net1366 s0.data_out\[11\]\[0\] _2050_ VPWR VGND sg13g2_and2_1
X_5113_ _1098_ _1097_ net1692 _1074_ net1697 VPWR VGND sg13g2_a22oi_1
XFILLER_33_0 VPWR VGND sg13g2_fill_2
X_6093_ net1367 net1354 _1982_ VPWR VGND sg13g2_nor2b_1
X_5044_ _1038_ VPWR _1039_ VGND net1178 _1037_ sg13g2_o21ai_1
XFILLER_26_704 VPWR VGND sg13g2_fill_1
XFILLER_27_29 VPWR VGND sg13g2_fill_2
XFILLER_25_225 VPWR VGND sg13g2_fill_2
X_6995_ _2793_ net1256 net505 VPWR VGND sg13g2_nand2_1
X_5946_ _1848_ _1849_ _1850_ VPWR VGND sg13g2_nor2_1
X_5877_ VGND VPWR _1670_ _1789_ _1790_ net1407 sg13g2_a21oi_1
XFILLER_40_239 VPWR VGND sg13g2_fill_2
X_7616_ net570 net1583 _3352_ _0100_ VPWR VGND sg13g2_a21o_1
X_4828_ VGND VPWR net1487 _0835_ _0837_ _0836_ sg13g2_a21oi_1
XFILLER_22_987 VPWR VGND sg13g2_decap_8
X_7547_ _3293_ VPWR _3294_ VGND net1202 _3292_ sg13g2_o21ai_1
X_4759_ s0.data_out\[23\]\[4\] s0.data_out\[22\]\[4\] net1503 _0780_ VPWR VGND sg13g2_mux2_1
X_7478_ _3228_ net1202 _3227_ VPWR VGND sg13g2_nand2_1
X_6429_ net1308 net549 _2285_ VPWR VGND sg13g2_and2_1
XFILLER_1_803 VPWR VGND sg13g2_decap_8
XFILLER_0_346 VPWR VGND sg13g2_fill_2
XFILLER_49_829 VPWR VGND sg13g2_decap_8
X_7753__267 VPWR VGND net267 sg13g2_tiehi
XFILLER_44_567 VPWR VGND sg13g2_fill_1
XFILLER_25_770 VPWR VGND sg13g2_fill_2
XFILLER_13_921 VPWR VGND sg13g2_fill_1
XFILLER_25_792 VPWR VGND sg13g2_fill_1
XFILLER_13_998 VPWR VGND sg13g2_decap_8
XFILLER_4_641 VPWR VGND sg13g2_fill_2
XFILLER_0_880 VPWR VGND sg13g2_decap_8
Xhold2 s0.genblk1\[2\].modules.bubble VPWR VGND net371 sg13g2_dlygate4sd3_1
XFILLER_48_851 VPWR VGND sg13g2_decap_8
X_6780_ s0.data_out\[7\]\[5\] s0.data_out\[6\]\[5\] net1281 _2602_ VPWR VGND sg13g2_mux2_1
X_3992_ VPWR _3368_ net412 VGND sg13g2_inv_1
XFILLER_23_718 VPWR VGND sg13g2_fill_1
X_5800_ net1630 _1657_ _1721_ VPWR VGND sg13g2_nor2_1
X_5731_ _1656_ net612 net1422 VPWR VGND sg13g2_nand2b_1
X_5662_ net1197 _3475_ _1597_ VPWR VGND sg13g2_nor2_1
X_4613_ net1508 net1329 _0646_ VPWR VGND sg13g2_nor2b_1
X_5593_ _1530_ s0.data_out\[15\]\[1\] net1432 VPWR VGND sg13g2_nand2b_1
X_7401_ _3161_ _3162_ _3163_ VPWR VGND sg13g2_nor2_1
X_7332_ net1640 net1225 _3097_ VPWR VGND sg13g2_nor2b_1
X_4544_ net1521 net478 _0585_ VPWR VGND sg13g2_and2_1
Xhold402 s0.valid_out\[25\][0] VPWR VGND net771 sg13g2_dlygate4sd3_1
Xhold435 s0.data_out\[9\]\[5\] VPWR VGND net804 sg13g2_dlygate4sd3_1
X_7263_ VGND VPWR _2930_ _3036_ _3037_ net1239 sg13g2_a21oi_1
Xhold413 _2957_ VPWR VGND net782 sg13g2_dlygate4sd3_1
Xhold424 s0.data_out\[4\]\[5\] VPWR VGND net793 sg13g2_dlygate4sd3_1
Xhold457 s0.shift_out\[26\][0] VPWR VGND net826 sg13g2_dlygate4sd3_1
Xhold468 s0.data_out\[20\]\[6\] VPWR VGND net837 sg13g2_dlygate4sd3_1
X_4475_ _0519_ VPWR _0520_ VGND net1529 _3422_ sg13g2_o21ai_1
Xhold446 _0212_ VPWR VGND net815 sg13g2_dlygate4sd3_1
X_6214_ _2091_ net523 net1372 VPWR VGND sg13g2_nand2b_1
X_7194_ VGND VPWR net1172 _2914_ _2974_ net1585 sg13g2_a21oi_1
X_6145_ s0.data_out\[12\]\[4\] s0.data_out\[11\]\[4\] net1375 _2034_ VPWR VGND sg13g2_mux2_1
X_6076_ net450 _1967_ _1968_ VPWR VGND sg13g2_nor2_1
X_5027_ _1001_ _1024_ _1025_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_512 VPWR VGND sg13g2_decap_4
X_6978_ VGND VPWR net1260 _2773_ _2776_ _2775_ sg13g2_a21oi_1
X_5929_ _1836_ VPWR _1837_ VGND net1748 net588 sg13g2_o21ai_1
XFILLER_21_250 VPWR VGND sg13g2_decap_8
XFILLER_21_261 VPWR VGND sg13g2_fill_2
XFILLER_5_416 VPWR VGND sg13g2_fill_1
XFILLER_0_143 VPWR VGND sg13g2_fill_1
XFILLER_49_626 VPWR VGND sg13g2_decap_8
XFILLER_1_688 VPWR VGND sg13g2_decap_8
XFILLER_23_1019 VPWR VGND sg13g2_decap_8
XFILLER_45_865 VPWR VGND sg13g2_decap_8
XFILLER_28_94 VPWR VGND sg13g2_fill_2
XFILLER_32_537 VPWR VGND sg13g2_fill_1
XFILLER_8_265 VPWR VGND sg13g2_decap_4
XFILLER_8_298 VPWR VGND sg13g2_fill_1
XFILLER_5_972 VPWR VGND sg13g2_decap_8
X_4260_ VGND VPWR net1558 _3623_ _3624_ _3619_ sg13g2_a21oi_1
X_4191_ net1546 _3553_ _3558_ VPWR VGND sg13g2_nor2_1
X_7950_ net42 VGND VPWR _0084_ s0.was_valid_out\[1\][0] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_7881_ net129 VGND VPWR _0015_ s0.shift_out\[7\][0] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_6901_ _2711_ net1275 _2710_ VPWR VGND sg13g2_nand2b_1
X_6832_ _0023_ net631 _2645_ _3517_ net1602 VPWR VGND sg13g2_a22oi_1
X_7808__208 VPWR VGND net208 sg13g2_tiehi
X_6763_ _2583_ net1275 _2584_ _2585_ VPWR VGND sg13g2_a21o_1
X_6694_ net1600 _2489_ _2523_ VPWR VGND sg13g2_nor2_1
X_5714_ VGND VPWR net1401 _1638_ _1639_ _1637_ sg13g2_a21oi_1
X_5645_ _1582_ _1581_ net1674 _1574_ net1683 VPWR VGND sg13g2_a22oi_1
Xhold210 s0.data_out\[23\]\[6\] VPWR VGND net579 sg13g2_dlygate4sd3_1
X_5576_ _1514_ _1515_ _1516_ VPWR VGND sg13g2_nor2_1
X_7315_ net1243 VPWR _3084_ VGND _3054_ _3083_ sg13g2_o21ai_1
X_4527_ _0488_ VPWR _0572_ VGND _0544_ _0547_ sg13g2_o21ai_1
Xhold232 s0.data_out\[24\]\[2\] VPWR VGND net601 sg13g2_dlygate4sd3_1
Xhold221 _0325_ VPWR VGND net590 sg13g2_dlygate4sd3_1
Xhold243 s0.data_out\[14\]\[3\] VPWR VGND net612 sg13g2_dlygate4sd3_1
Xhold276 s0.data_out\[19\]\[6\] VPWR VGND net645 sg13g2_dlygate4sd3_1
Xhold265 s0.data_out\[19\]\[2\] VPWR VGND net634 sg13g2_dlygate4sd3_1
X_4458_ net1521 net1356 _0503_ VPWR VGND sg13g2_nor2b_1
Xhold287 _0247_ VPWR VGND net656 sg13g2_dlygate4sd3_1
Xhold254 s0.data_out\[10\]\[0\] VPWR VGND net623 sg13g2_dlygate4sd3_1
X_7246_ VGND VPWR _2900_ _3019_ _3020_ net1242 sg13g2_a21oi_1
Xhold298 _0045_ VPWR VGND net667 sg13g2_dlygate4sd3_1
X_7177_ _2960_ VPWR _2961_ VGND net1716 net716 sg13g2_o21ai_1
X_6128_ _2017_ s0.data_out\[11\]\[7\] net1387 VPWR VGND sg13g2_nand2b_1
X_4389_ _0444_ net1533 _0445_ _0446_ VPWR VGND sg13g2_a21o_1
X_6059_ net1392 VPWR _1954_ VGND _1902_ _1953_ sg13g2_o21ai_1
XFILLER_27_854 VPWR VGND sg13g2_fill_1
XFILLER_42_846 VPWR VGND sg13g2_fill_1
XFILLER_14_548 VPWR VGND sg13g2_fill_2
X_7898__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_14_74 VPWR VGND sg13g2_fill_1
XFILLER_14_85 VPWR VGND sg13g2_fill_1
XFILLER_5_246 VPWR VGND sg13g2_fill_1
XFILLER_2_931 VPWR VGND sg13g2_decap_8
XFILLER_33_868 VPWR VGND sg13g2_fill_2
X_5430_ _1383_ net1744 _1384_ VPWR VGND _1323_ sg13g2_nand3b_1
XFILLER_9_574 VPWR VGND sg13g2_fill_1
X_5361_ _1322_ net753 net1455 VPWR VGND sg13g2_nand2b_1
X_4312_ net1558 VPWR _0373_ VGND _3602_ _0372_ sg13g2_o21ai_1
X_5292_ net1204 _3460_ _1261_ VPWR VGND sg13g2_nor2_1
X_7100_ VGND VPWR net1240 _2884_ _2886_ _2885_ sg13g2_a21oi_1
X_4243_ net1558 _3605_ _3606_ _3607_ VPWR VGND sg13g2_nor3_1
X_7814__201 VPWR VGND net201 sg13g2_tiehi
X_7031_ _2827_ net1252 _2828_ _2829_ VPWR VGND sg13g2_a21o_1
X_4174_ VGND VPWR net1571 net1166 net5 _3547_ sg13g2_a21oi_1
XFILLER_28_629 VPWR VGND sg13g2_fill_1
XFILLER_49_990 VPWR VGND sg13g2_decap_8
X_7933_ net73 VGND VPWR _0067_ s0.data_out\[3\]\[3\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_7864_ net148 VGND VPWR _0342_ s0.data_out\[9\]\[6\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_6815_ VGND VPWR net1176 _2597_ _2632_ net1601 sg13g2_a21oi_1
X_7795_ net222 VGND VPWR _0273_ s0.data_out\[14\]\[4\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_6746_ net1272 net1347 _2568_ VPWR VGND sg13g2_nor2b_1
X_6677_ _2455_ _2509_ net1731 _2510_ VPWR VGND sg13g2_nand3_1
X_5628_ VGND VPWR _1565_ _1556_ net1655 sg13g2_or2_1
X_5559_ net1429 s0.data_out\[16\]\[6\] _1501_ VPWR VGND sg13g2_and2_1
Xfanout1507 s0.valid_out\[22\][0] net1507 VPWR VGND sg13g2_buf_1
Xfanout1518 s0.valid_out\[23\][0] net1518 VPWR VGND sg13g2_buf_8
Xfanout1529 net1532 net1529 VPWR VGND sg13g2_buf_1
X_7229_ s0.data_out\[2\]\[0\] s0.data_out\[3\]\[0\] net1247 _3003_ VPWR VGND sg13g2_mux2_1
XFILLER_47_927 VPWR VGND sg13g2_decap_8
XFILLER_19_629 VPWR VGND sg13g2_decap_4
XFILLER_42_621 VPWR VGND sg13g2_fill_2
XFILLER_41_120 VPWR VGND sg13g2_fill_2
XFILLER_14_345 VPWR VGND sg13g2_fill_2
XFILLER_26_183 VPWR VGND sg13g2_fill_1
XFILLER_41_153 VPWR VGND sg13g2_fill_1
XFILLER_6_566 VPWR VGND sg13g2_fill_2
XFILLER_46_960 VPWR VGND sg13g2_decap_8
XFILLER_18_640 VPWR VGND sg13g2_fill_1
X_4930_ _0932_ VPWR _0933_ VGND net1734 net755 sg13g2_o21ai_1
XFILLER_17_150 VPWR VGND sg13g2_fill_2
XFILLER_36_1007 VPWR VGND sg13g2_decap_8
X_4861_ _0868_ net1482 _0869_ _0870_ VPWR VGND sg13g2_a21o_1
X_6600_ net1730 net383 _0002_ VPWR VGND sg13g2_and2_1
X_7580_ VGND VPWR net1214 net404 _3318_ net1209 sg13g2_a21oi_1
X_4792_ net1594 _0747_ _0809_ VPWR VGND sg13g2_nor2_1
XFILLER_20_348 VPWR VGND sg13g2_fill_1
X_6531_ _2373_ _2375_ net1676 _2377_ VPWR VGND sg13g2_nand3_1
X_6462_ VPWR _2311_ _2310_ VGND sg13g2_inv_1
X_6393_ _2251_ _2250_ net1663 _2243_ net1653 VPWR VGND sg13g2_a22oi_1
X_5413_ _1290_ _1370_ net1743 _1371_ VPWR VGND sg13g2_nand3_1
X_5344_ _1304_ VPWR _1305_ VGND net1203 _1302_ sg13g2_o21ai_1
X_5275_ _1226_ _1243_ _1248_ VPWR VGND sg13g2_nor2b_1
X_4226_ _3590_ net1557 net452 VPWR VGND sg13g2_nand2_1
X_7014_ _2810_ net1251 _2811_ _2812_ VPWR VGND sg13g2_a21o_1
X_4157_ VPWR _3533_ net505 VGND sg13g2_inv_1
X_4088_ _3464_ s0.data_out\[17\]\[2\] VPWR VGND sg13g2_inv_2
XFILLER_37_982 VPWR VGND sg13g2_decap_8
X_7916_ net91 VGND VPWR _0050_ s0.genblk1\[3\].modules.bubble clknet_leaf_2_clk sg13g2_dfrbpq_1
X_7749__272 VPWR VGND net272 sg13g2_tiehi
X_7847_ net166 VGND VPWR net590 s0.data_out\[10\]\[1\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_11_315 VPWR VGND sg13g2_fill_2
X_7778_ net240 VGND VPWR _0256_ s0.shift_out\[15\][0] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_7895__114 VPWR VGND net114 sg13g2_tiehi
X_6729_ _2551_ net1278 net694 VPWR VGND sg13g2_nand2_1
XFILLER_11_42 VPWR VGND sg13g2_fill_2
Xfanout1304 s0.valid_out\[8\][0] net1304 VPWR VGND sg13g2_buf_8
Xfanout1337 s0.data_new_delayed\[6\] net1337 VPWR VGND sg13g2_buf_8
Xfanout1326 net1327 net1326 VPWR VGND sg13g2_buf_1
Xfanout1348 s0.data_new_delayed\[2\] net1348 VPWR VGND sg13g2_buf_8
Xfanout1315 net1318 net1315 VPWR VGND sg13g2_buf_8
Xfanout1359 s0.data_new_delayed\[0\] net1359 VPWR VGND sg13g2_buf_8
XFILLER_47_724 VPWR VGND sg13g2_decap_8
XFILLER_28_971 VPWR VGND sg13g2_decap_8
XFILLER_15_621 VPWR VGND sg13g2_fill_2
XFILLER_43_963 VPWR VGND sg13g2_decap_8
XFILLER_27_492 VPWR VGND sg13g2_fill_2
XFILLER_30_668 VPWR VGND sg13g2_fill_2
X_5060_ net1469 net837 _1051_ VPWR VGND sg13g2_and2_1
X_4011_ VPWR _3387_ net1230 VGND sg13g2_inv_1
XFILLER_26_919 VPWR VGND sg13g2_fill_2
XFILLER_19_993 VPWR VGND sg13g2_decap_8
X_5962_ _1863_ net1193 _1862_ VPWR VGND sg13g2_nand2_1
X_7701_ net324 VGND VPWR net553 s0.data_out\[22\]\[6\] clknet_leaf_41_clk sg13g2_dfrbpq_2
X_4913_ net1180 _3444_ _0919_ VPWR VGND sg13g2_nor2_1
XFILLER_18_481 VPWR VGND sg13g2_fill_1
XFILLER_18_492 VPWR VGND sg13g2_fill_1
XFILLER_34_963 VPWR VGND sg13g2_decap_8
X_5893_ net1394 net1341 _1806_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_440 VPWR VGND sg13g2_decap_4
X_7632_ net54 VGND VPWR _0110_ s0.valid_out\[27\][0] clknet_leaf_0_clk sg13g2_dfrbpq_2
X_4844_ _0853_ net1501 _0852_ VPWR VGND sg13g2_nand2b_1
X_7563_ _3306_ VPWR _3307_ VGND net1722 net733 sg13g2_o21ai_1
X_4775_ VGND VPWR _0791_ _0794_ _0160_ _0795_ sg13g2_a21oi_1
X_6514_ net1298 net1334 _2360_ VPWR VGND sg13g2_nor2b_1
X_7494_ s0.data_out\[0\]\[7\] s0.data_out\[1\]\[7\] net1225 _3244_ VPWR VGND sg13g2_mux2_1
X_6445_ VPWR _0328_ _2297_ VGND sg13g2_inv_1
X_6376_ VGND VPWR net1320 _2231_ _2234_ _2233_ sg13g2_a21oi_1
X_5327_ VGND VPWR net1437 _1286_ _1288_ _1287_ sg13g2_a21oi_1
X_5258_ _1231_ net1462 _1230_ VPWR VGND sg13g2_nand2b_1
X_5189_ net1199 _3451_ _1166_ VPWR VGND sg13g2_nor2_1
X_4209_ _3572_ VPWR _3573_ VGND net1554 _3417_ sg13g2_o21ai_1
XFILLER_24_440 VPWR VGND sg13g2_fill_2
XFILLER_25_974 VPWR VGND sg13g2_decap_8
XFILLER_40_955 VPWR VGND sg13g2_decap_8
XFILLER_11_123 VPWR VGND sg13g2_fill_2
XFILLER_11_134 VPWR VGND sg13g2_fill_2
XFILLER_4_834 VPWR VGND sg13g2_fill_1
XFILLER_4_878 VPWR VGND sg13g2_decap_8
XFILLER_3_388 VPWR VGND sg13g2_fill_1
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
Xfanout1167 net1169 net1167 VPWR VGND sg13g2_buf_8
Xfanout1178 net1179 net1178 VPWR VGND sg13g2_buf_8
Xfanout1189 _3387_ net1189 VPWR VGND sg13g2_buf_8
XFILLER_34_226 VPWR VGND sg13g2_fill_1
XFILLER_15_440 VPWR VGND sg13g2_fill_1
X_4560_ _0597_ net1716 _0598_ VPWR VGND _0542_ sg13g2_nand3b_1
XFILLER_31_999 VPWR VGND sg13g2_decap_8
X_4491_ VGND VPWR net1537 _0533_ _0536_ _0535_ sg13g2_a21oi_1
X_6230_ _2107_ _3383_ _2106_ VPWR VGND sg13g2_nand2_1
X_6161_ VGND VPWR _2044_ _2048_ _0292_ _2049_ sg13g2_a21oi_1
X_5112_ VGND VPWR net1475 _1094_ _1097_ _1096_ sg13g2_a21oi_1
X_6092_ VGND VPWR _1981_ _1980_ net1698 sg13g2_or2_1
X_5043_ VGND VPWR net1178 _0954_ _1038_ net1607 sg13g2_a21oi_1
Xfanout1690 net1694 net1690 VPWR VGND sg13g2_buf_8
X_6994_ _2777_ VPWR _2792_ VGND net1703 _2784_ sg13g2_o21ai_1
XFILLER_25_237 VPWR VGND sg13g2_decap_4
X_5945_ net1645 net1389 _1849_ VPWR VGND sg13g2_nor2b_1
X_5876_ _1789_ s0.data_out\[13\]\[6\] net1410 VPWR VGND sg13g2_nand2b_1
X_7746__275 VPWR VGND net275 sg13g2_tiehi
X_7615_ VGND VPWR _3330_ _3331_ _3352_ net1583 sg13g2_a21oi_1
X_4827_ net1487 net1351 _0836_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_454 VPWR VGND sg13g2_fill_2
X_7546_ VGND VPWR net1201 _3215_ _3293_ net1583 sg13g2_a21oi_1
X_4758_ net1494 net1344 _0779_ VPWR VGND sg13g2_nor2b_1
X_7477_ s0.data_out\[0\]\[0\] s0.data_out\[1\]\[0\] net1225 _3227_ VPWR VGND sg13g2_mux2_1
X_4689_ _0711_ VPWR _0713_ VGND s0.was_valid_out\[22\][0] net1503 sg13g2_o21ai_1
X_7892__117 VPWR VGND net117 sg13g2_tiehi
X_6428_ VPWR _0324_ _2284_ VGND sg13g2_inv_1
XFILLER_1_859 VPWR VGND sg13g2_decap_8
X_6359_ _2217_ net549 net1360 VPWR VGND sg13g2_nand2b_1
XFILLER_49_808 VPWR VGND sg13g2_decap_8
XFILLER_48_329 VPWR VGND sg13g2_fill_2
XFILLER_17_705 VPWR VGND sg13g2_fill_2
XFILLER_16_226 VPWR VGND sg13g2_decap_4
XFILLER_12_443 VPWR VGND sg13g2_fill_1
XFILLER_13_977 VPWR VGND sg13g2_decap_8
XFILLER_24_292 VPWR VGND sg13g2_decap_8
XFILLER_32_1010 VPWR VGND sg13g2_decap_8
XFILLER_12_498 VPWR VGND sg13g2_decap_4
XFILLER_48_830 VPWR VGND sg13g2_decap_8
XFILLER_39_318 VPWR VGND sg13g2_fill_1
Xhold3 s0.genblk1\[19\].modules.bubble VPWR VGND net372 sg13g2_dlygate4sd3_1
XFILLER_47_362 VPWR VGND sg13g2_fill_1
XFILLER_35_513 VPWR VGND sg13g2_decap_4
XFILLER_47_395 VPWR VGND sg13g2_fill_2
X_3991_ VPWR _3367_ net437 VGND sg13g2_inv_1
X_5730_ _1653_ net1403 _1654_ _1655_ VPWR VGND sg13g2_a21o_1
X_5661_ VPWR _0245_ _1596_ VGND sg13g2_inv_1
X_7400_ _3154_ _3151_ _3162_ VPWR VGND _3152_ sg13g2_nand3b_1
X_4612_ s0.data_out\[24\]\[7\] s0.data_out\[23\]\[7\] net1515 _0645_ VPWR VGND sg13g2_mux2_1
X_5592_ _1527_ net1412 _1528_ _1529_ VPWR VGND sg13g2_a21o_1
X_4543_ VPWR _0139_ net763 VGND sg13g2_inv_1
X_7331_ net1230 VPWR _3096_ VGND net1639 net1218 sg13g2_o21ai_1
Xhold425 s0.data_out\[3\]\[3\] VPWR VGND net794 sg13g2_dlygate4sd3_1
Xhold436 s0.data_out\[18\]\[7\] VPWR VGND net805 sg13g2_dlygate4sd3_1
Xhold414 s0.data_out\[16\]\[0\] VPWR VGND net783 sg13g2_dlygate4sd3_1
X_7262_ _3036_ net568 net1247 VPWR VGND sg13g2_nand2b_1
Xhold403 s0.data_out\[15\]\[6\] VPWR VGND net772 sg13g2_dlygate4sd3_1
X_4474_ _0519_ net1529 net478 VPWR VGND sg13g2_nand2_1
Xhold447 s0.data_out\[23\]\[1\] VPWR VGND net816 sg13g2_dlygate4sd3_1
Xhold458 s0.valid_out\[5\][0] VPWR VGND net827 sg13g2_dlygate4sd3_1
X_6213_ _2088_ net1322 _2089_ _2090_ VPWR VGND sg13g2_a21o_1
X_7193_ VGND VPWR net1242 net503 _2973_ _2911_ sg13g2_a21oi_1
X_6144_ _2033_ net1372 net787 VPWR VGND sg13g2_nand2_1
X_6075_ _1966_ VPWR _1967_ VGND net1380 _1849_ sg13g2_o21ai_1
X_5026_ _1009_ VPWR _1024_ VGND _1017_ _1019_ sg13g2_o21ai_1
X_6977_ VGND VPWR _2668_ _2774_ _2775_ net1260 sg13g2_a21oi_1
X_5928_ _1835_ VPWR _1836_ VGND net1195 _1834_ sg13g2_o21ai_1
XFILLER_16_1016 VPWR VGND sg13g2_decap_8
XFILLER_16_1027 VPWR VGND sg13g2_fill_2
XFILLER_21_240 VPWR VGND sg13g2_decap_4
X_5859_ _1770_ net1391 _1771_ _1772_ VPWR VGND sg13g2_a21o_1
XFILLER_10_969 VPWR VGND sg13g2_decap_8
X_7529_ _3278_ _3243_ _3279_ VPWR VGND _3259_ sg13g2_nand3b_1
XFILLER_0_100 VPWR VGND sg13g2_fill_1
XFILLER_49_605 VPWR VGND sg13g2_decap_8
XFILLER_45_800 VPWR VGND sg13g2_fill_1
XFILLER_45_844 VPWR VGND sg13g2_decap_8
XFILLER_17_524 VPWR VGND sg13g2_fill_1
XFILLER_44_398 VPWR VGND sg13g2_fill_2
XFILLER_5_951 VPWR VGND sg13g2_decap_8
X_4190_ _3554_ VPWR _3557_ VGND net524 net1554 sg13g2_o21ai_1
XFILLER_39_115 VPWR VGND sg13g2_fill_1
XFILLER_39_104 VPWR VGND sg13g2_fill_2
X_7880_ net130 VGND VPWR _0014_ s0.genblk1\[6\].modules.bubble clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_6900_ VGND VPWR net1265 _2708_ _2710_ _2709_ sg13g2_a21oi_1
XFILLER_35_332 VPWR VGND sg13g2_fill_1
X_6831_ net1602 net415 _2645_ VPWR VGND sg13g2_nor2_1
XFILLER_39_1027 VPWR VGND sg13g2_fill_2
XFILLER_36_877 VPWR VGND sg13g2_fill_2
X_6762_ net1275 net1334 _2584_ VPWR VGND sg13g2_nor2b_1
X_6693_ net1296 VPWR _2522_ VGND _2486_ _2521_ sg13g2_o21ai_1
X_5713_ s0.data_out\[15\]\[0\] s0.data_out\[14\]\[0\] net1408 _1638_ VPWR VGND sg13g2_mux2_1
X_5644_ VGND VPWR net1426 _1578_ _1581_ _1580_ sg13g2_a21oi_1
X_7743__278 VPWR VGND net278 sg13g2_tiehi
X_7314_ net1188 _3539_ _3083_ VPWR VGND sg13g2_nor2_1
Xhold211 s0.data_out\[5\]\[2\] VPWR VGND net580 sg13g2_dlygate4sd3_1
X_5575_ VGND VPWR _3365_ _3376_ _1515_ net1428 sg13g2_a21oi_1
Xhold200 _0083_ VPWR VGND net569 sg13g2_dlygate4sd3_1
X_4526_ VGND VPWR _0556_ _0564_ _0571_ _0548_ sg13g2_a21oi_1
Xhold233 _0151_ VPWR VGND net602 sg13g2_dlygate4sd3_1
Xhold222 s0.data_out\[20\]\[2\] VPWR VGND net591 sg13g2_dlygate4sd3_1
Xhold244 _0272_ VPWR VGND net613 sg13g2_dlygate4sd3_1
XFILLER_49_28 VPWR VGND sg13g2_fill_2
XFILLER_46_1009 VPWR VGND sg13g2_decap_8
Xhold277 _0215_ VPWR VGND net646 sg13g2_dlygate4sd3_1
X_4457_ _0502_ net1185 _0501_ VPWR VGND sg13g2_nand2_1
Xhold266 _0211_ VPWR VGND net635 sg13g2_dlygate4sd3_1
Xhold255 s0.data_out\[13\]\[2\] VPWR VGND net624 sg13g2_dlygate4sd3_1
X_7245_ _3019_ net735 net1245 VPWR VGND sg13g2_nand2b_1
Xhold299 s0.data_out\[5\]\[4\] VPWR VGND net668 sg13g2_dlygate4sd3_1
X_7176_ _2959_ VPWR _2960_ VGND net1170 _2958_ sg13g2_o21ai_1
Xhold288 s0.data_out\[14\]\[0\] VPWR VGND net657 sg13g2_dlygate4sd3_1
X_6127_ _2014_ net1370 _2015_ _2016_ VPWR VGND sg13g2_a21o_1
X_4388_ net1533 net1338 _0445_ VPWR VGND sg13g2_nor2b_1
XFILLER_46_608 VPWR VGND sg13g2_fill_2
X_6058_ net1382 s0.data_out\[12\]\[5\] _1953_ VPWR VGND sg13g2_and2_1
X_5009_ VGND VPWR _0886_ _1006_ _1007_ net1484 sg13g2_a21oi_1
XFILLER_14_538 VPWR VGND sg13g2_fill_1
XFILLER_2_910 VPWR VGND sg13g2_decap_8
XFILLER_7_1025 VPWR VGND sg13g2_decap_4
XFILLER_2_987 VPWR VGND sg13g2_decap_8
XFILLER_1_486 VPWR VGND sg13g2_fill_1
XFILLER_36_107 VPWR VGND sg13g2_decap_4
XFILLER_44_195 VPWR VGND sg13g2_decap_4
XFILLER_32_324 VPWR VGND sg13g2_fill_1
XFILLER_13_560 VPWR VGND sg13g2_fill_1
XFILLER_9_542 VPWR VGND sg13g2_fill_2
X_7697__328 VPWR VGND net328 sg13g2_tiehi
X_5360_ _1319_ net1441 _1320_ _1321_ VPWR VGND sg13g2_a21o_1
X_4311_ net1544 s0.data_out\[26\]\[7\] _0372_ VPWR VGND sg13g2_and2_1
X_5291_ _0211_ _1259_ _1260_ _3455_ net1619 VPWR VGND sg13g2_a22oi_1
XFILLER_4_280 VPWR VGND sg13g2_fill_2
X_4242_ net1563 s0.data_out\[26\]\[6\] _3606_ VPWR VGND sg13g2_nor2_1
X_7030_ net1252 net1338 _2828_ VPWR VGND sg13g2_nor2b_1
X_4173_ s0.data_out\[27\]\[2\] net1166 _3547_ VPWR VGND sg13g2_nor2_1
X_7932_ net74 VGND VPWR _0066_ s0.data_out\[3\]\[2\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_7863_ net149 VGND VPWR _0341_ s0.data_out\[9\]\[5\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_6814_ VGND VPWR net1276 net518 _2631_ _2593_ sg13g2_a21oi_1
X_7794_ net223 VGND VPWR net613 s0.data_out\[14\]\[3\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_11_508 VPWR VGND sg13g2_fill_2
X_6745_ s0.data_out\[7\]\[3\] s0.data_out\[6\]\[3\] net1279 _2567_ VPWR VGND sg13g2_mux2_1
XFILLER_32_891 VPWR VGND sg13g2_fill_1
XFILLER_13_1019 VPWR VGND sg13g2_decap_8
X_6676_ net1294 VPWR _2509_ VGND _2451_ _2508_ sg13g2_o21ai_1
X_5627_ _1564_ _1563_ net1665 _1556_ net1654 VPWR VGND sg13g2_a22oi_1
XFILLER_3_707 VPWR VGND sg13g2_fill_2
X_5558_ VPWR _0238_ _1500_ VGND sg13g2_inv_1
X_4509_ _0443_ VPWR _0554_ VGND net1543 _3427_ sg13g2_o21ai_1
X_5489_ _1438_ net527 net1446 VPWR VGND sg13g2_nand2b_1
X_7228_ VGND VPWR net1228 _3000_ _3002_ _3001_ sg13g2_a21oi_1
Xfanout1508 net1511 net1508 VPWR VGND sg13g2_buf_2
Xfanout1519 net1520 net1519 VPWR VGND sg13g2_buf_2
XFILLER_47_906 VPWR VGND sg13g2_decap_8
X_7159_ net1649 _2936_ _2945_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_38_clk clknet_3_4__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_27_663 VPWR VGND sg13g2_decap_8
XFILLER_15_814 VPWR VGND sg13g2_fill_2
XFILLER_25_63 VPWR VGND sg13g2_fill_1
XFILLER_10_585 VPWR VGND sg13g2_fill_2
XFILLER_6_589 VPWR VGND sg13g2_fill_2
XFILLER_2_784 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_3_5__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_33_600 VPWR VGND sg13g2_fill_1
X_4860_ net1482 net1330 _0869_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_165 VPWR VGND sg13g2_fill_1
X_6530_ _2376_ _2373_ _2375_ VPWR VGND sg13g2_nand2_1
X_4791_ net1513 VPWR _0808_ VGND _0744_ _0807_ sg13g2_o21ai_1
XFILLER_20_327 VPWR VGND sg13g2_fill_2
XFILLER_13_390 VPWR VGND sg13g2_fill_1
X_6461_ _2308_ _2309_ _2310_ VPWR VGND sg13g2_nor2_1
X_6392_ VGND VPWR net1323 _2247_ _2250_ _2249_ sg13g2_a21oi_1
X_5412_ net1449 VPWR _1370_ VGND _1287_ _1369_ sg13g2_o21ai_1
X_5343_ _1304_ net1203 _1303_ VPWR VGND sg13g2_nand2_1
X_5274_ _1226_ _1243_ _1244_ _1246_ _1247_ VPWR VGND sg13g2_nor4_1
X_4225_ VGND VPWR net1564 _3410_ _3589_ _3588_ sg13g2_a21oi_1
X_7013_ net1251 net1333 _2811_ VPWR VGND sg13g2_nor2b_1
X_7888__122 VPWR VGND net122 sg13g2_tiehi
X_4156_ VPWR _3532_ net536 VGND sg13g2_inv_1
XFILLER_28_416 VPWR VGND sg13g2_fill_1
XFILLER_37_961 VPWR VGND sg13g2_decap_8
X_4087_ _3463_ net542 VPWR VGND sg13g2_inv_2
X_7915_ net92 VGND VPWR _0049_ s0.valid_out\[4\][0] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_7846_ net167 VGND VPWR _0324_ s0.data_out\[10\]\[0\] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_12_806 VPWR VGND sg13g2_fill_1
X_7777_ net241 VGND VPWR _0255_ s0.genblk1\[14\].modules.bubble clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_4989_ _0985_ net1468 _0986_ _0987_ VPWR VGND sg13g2_a21o_1
X_6728_ VGND VPWR _2550_ _2549_ net1696 sg13g2_or2_1
X_6659_ _2491_ net1286 _2492_ _2493_ VPWR VGND sg13g2_a21o_1
XFILLER_20_894 VPWR VGND sg13g2_fill_2
XFILLER_3_515 VPWR VGND sg13g2_fill_2
XFILLER_3_504 VPWR VGND sg13g2_fill_1
Xfanout1305 net1313 net1305 VPWR VGND sg13g2_buf_8
Xfanout1316 net1318 net1316 VPWR VGND sg13g2_buf_2
Xfanout1327 s0.shift_out\[10\][0] net1327 VPWR VGND sg13g2_buf_2
Xfanout1338 net1339 net1338 VPWR VGND sg13g2_buf_8
XFILLER_47_703 VPWR VGND sg13g2_decap_8
Xfanout1349 net822 net1349 VPWR VGND sg13g2_buf_8
XFILLER_46_235 VPWR VGND sg13g2_fill_1
XFILLER_43_942 VPWR VGND sg13g2_decap_8
XFILLER_42_474 VPWR VGND sg13g2_fill_2
X_7804__212 VPWR VGND net212 sg13g2_tiehi
XFILLER_7_898 VPWR VGND sg13g2_fill_2
X_7811__205 VPWR VGND net205 sg13g2_tiehi
X_4010_ VPWR _3386_ net1561 VGND sg13g2_inv_1
XFILLER_28_4 VPWR VGND sg13g2_fill_2
XFILLER_38_758 VPWR VGND sg13g2_decap_4
XFILLER_25_419 VPWR VGND sg13g2_decap_4
X_5961_ _1746_ VPWR _1862_ VGND net1397 _3490_ sg13g2_o21ai_1
X_7700_ net325 VGND VPWR _0178_ s0.data_out\[22\]\[5\] clknet_leaf_41_clk sg13g2_dfrbpq_2
X_4912_ _0174_ _0917_ _0918_ _3440_ net1605 VPWR VGND sg13g2_a22oi_1
X_5892_ s0.data_out\[14\]\[5\] s0.data_out\[13\]\[5\] net1400 _1805_ VPWR VGND sg13g2_mux2_1
X_7631_ net56 VGND VPWR net677 s0.was_valid_out\[27\][0] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4843_ VGND VPWR net1486 _0850_ _0852_ _0851_ sg13g2_a21oi_1
X_7562_ _3305_ VPWR _3306_ VGND net1201 _3304_ sg13g2_o21ai_1
X_4774_ VGND VPWR _0795_ net1566 net375 sg13g2_or2_1
X_6513_ s0.data_out\[9\]\[6\] s0.data_out\[8\]\[6\] net1304 _2359_ VPWR VGND sg13g2_mux2_1
X_7493_ _3242_ VPWR _3243_ VGND _3234_ _3235_ sg13g2_o21ai_1
Xclkbuf_leaf_9_clk clknet_3_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_6444_ _2296_ VPWR _2297_ VGND net1738 net747 sg13g2_o21ai_1
X_6375_ VGND VPWR _2110_ _2232_ _2233_ net1320 sg13g2_a21oi_1
X_5326_ net1437 net1350 _1287_ VPWR VGND sg13g2_nor2b_1
X_5257_ VGND VPWR net1450 _1228_ _1230_ _1229_ sg13g2_a21oi_1
X_7637__49 VPWR VGND net49 sg13g2_tiehi
X_4208_ _3572_ net1555 net621 VPWR VGND sg13g2_nand2_1
X_5188_ VPWR _0203_ _1165_ VGND sg13g2_inv_1
XFILLER_29_725 VPWR VGND sg13g2_decap_8
X_4139_ VPWR _3515_ net593 VGND sg13g2_inv_1
XFILLER_19_1014 VPWR VGND sg13g2_decap_8
XFILLER_40_934 VPWR VGND sg13g2_decap_8
X_7829_ net185 VGND VPWR _0307_ s0.data_out\[11\]\[2\] clknet_leaf_26_clk sg13g2_dfrbpq_2
XFILLER_22_20 VPWR VGND sg13g2_fill_2
XFILLER_4_824 VPWR VGND sg13g2_fill_2
XFILLER_47_511 VPWR VGND sg13g2_fill_1
Xfanout1179 net1180 net1179 VPWR VGND sg13g2_buf_1
Xfanout1168 net1169 net1168 VPWR VGND sg13g2_buf_8
XFILLER_31_901 VPWR VGND sg13g2_decap_8
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_31_978 VPWR VGND sg13g2_decap_8
X_4490_ VGND VPWR _0424_ _0534_ _0535_ net1537 sg13g2_a21oi_1
X_7739__283 VPWR VGND net283 sg13g2_tiehi
X_6160_ VGND VPWR _2049_ net1568 net377 sg13g2_or2_1
X_5111_ VGND VPWR _0974_ _1095_ _1096_ net1476 sg13g2_a21oi_1
XFILLER_33_2 VPWR VGND sg13g2_fill_1
X_6091_ VGND VPWR net1377 _1977_ _1980_ _1979_ sg13g2_a21oi_1
X_5042_ VGND VPWR net1470 s0.data_out\[20\]\[2\] _1037_ _0952_ sg13g2_a21oi_1
Xfanout1680 net1681 net1680 VPWR VGND sg13g2_buf_2
X_7885__125 VPWR VGND net125 sg13g2_tiehi
Xfanout1691 net1694 net1691 VPWR VGND sg13g2_buf_8
XFILLER_38_588 VPWR VGND sg13g2_fill_1
X_6993_ VPWR VGND _2790_ net1710 _2788_ net1703 _2791_ _2784_ sg13g2_a221oi_1
XFILLER_25_227 VPWR VGND sg13g2_fill_1
X_5944_ net1393 VPWR _1848_ VGND net1644 net1384 sg13g2_o21ai_1
XFILLER_34_750 VPWR VGND sg13g2_fill_2
X_5875_ _1786_ net1395 _1787_ _1788_ VPWR VGND sg13g2_a21o_1
X_7614_ VGND VPWR _3349_ _3350_ _0099_ _3351_ sg13g2_a21oi_1
X_4826_ s0.data_out\[22\]\[2\] s0.data_out\[21\]\[2\] net1491 _0835_ VPWR VGND sg13g2_mux2_1
X_7545_ VGND VPWR net1212 net459 _3292_ _3217_ sg13g2_a21oi_1
X_4757_ _0775_ _0777_ net1671 _0778_ VPWR VGND sg13g2_nand3_1
X_7476_ VGND VPWR net1218 _3225_ _3226_ _3222_ sg13g2_a21oi_1
X_4688_ VGND VPWR net1181 _0604_ _0712_ _0711_ sg13g2_a21oi_1
XFILLER_49_1018 VPWR VGND sg13g2_decap_8
X_6427_ _2283_ VPWR _2284_ VGND net1738 net623 sg13g2_o21ai_1
X_6358_ _2215_ net1308 _2213_ _2216_ VPWR VGND sg13g2_a21o_1
XFILLER_1_838 VPWR VGND sg13g2_decap_8
X_5309_ net1205 _3457_ _1274_ VPWR VGND sg13g2_nor2_1
X_6289_ VPWR _0305_ _2164_ VGND sg13g2_inv_1
XFILLER_16_205 VPWR VGND sg13g2_fill_2
X_7801__215 VPWR VGND net215 sg13g2_tiehi
Xhold4 s0.genblk1\[13\].modules.bubble VPWR VGND net373 sg13g2_dlygate4sd3_1
XFILLER_48_886 VPWR VGND sg13g2_decap_8
X_3990_ VPWR _3366_ net428 VGND sg13g2_inv_1
X_5660_ _1595_ VPWR _1596_ VGND net1743 net783 sg13g2_o21ai_1
X_4611_ _0644_ net1516 net662 VPWR VGND sg13g2_nand2_1
X_5591_ net1412 net1354 _1528_ VPWR VGND sg13g2_nor2b_1
XFILLER_30_274 VPWR VGND sg13g2_fill_2
XFILLER_8_982 VPWR VGND sg13g2_decap_8
X_4542_ _0583_ VPWR _0584_ VGND net1725 net762 sg13g2_o21ai_1
X_7330_ _0071_ _3094_ _3095_ _3535_ net1582 VPWR VGND sg13g2_a22oi_1
Xhold415 s0.data_out\[20\]\[6\] VPWR VGND net784 sg13g2_dlygate4sd3_1
X_4473_ net1701 _0500_ _0518_ VPWR VGND sg13g2_nor2_1
Xhold426 s0.data_out\[3\]\[0\] VPWR VGND net795 sg13g2_dlygate4sd3_1
X_7261_ _3033_ net1231 _3034_ _3035_ VPWR VGND sg13g2_a21o_1
Xhold404 _1733_ VPWR VGND net773 sg13g2_dlygate4sd3_1
Xhold448 _0162_ VPWR VGND net817 sg13g2_dlygate4sd3_1
Xhold437 s0.data_out\[8\]\[0\] VPWR VGND net806 sg13g2_dlygate4sd3_1
Xhold459 s0.valid_out\[2\][0] VPWR VGND net828 sg13g2_dlygate4sd3_1
X_6212_ net1321 net1351 _2089_ VPWR VGND sg13g2_nor2b_1
X_7192_ VPWR _0056_ net671 VGND sg13g2_inv_1
X_6143_ _2031_ VPWR _2032_ VGND net1694 _2003_ sg13g2_o21ai_1
X_6074_ VPWR _1966_ _1965_ VGND sg13g2_inv_1
XFILLER_39_853 VPWR VGND sg13g2_fill_2
X_5025_ _0983_ _1001_ _1022_ _1023_ VPWR VGND sg13g2_or3_1
XFILLER_0_1020 VPWR VGND sg13g2_decap_8
X_6976_ _2774_ s0.data_out\[4\]\[2\] net1266 VPWR VGND sg13g2_nand2b_1
X_5927_ VGND VPWR _3381_ _1801_ _1835_ net1629 sg13g2_a21oi_1
X_5858_ net1391 net1169 _1771_ VPWR VGND sg13g2_nor2_1
X_4809_ net1512 VPWR _0822_ VGND _0755_ _0821_ sg13g2_o21ai_1
XFILLER_22_797 VPWR VGND sg13g2_fill_2
X_5789_ net1195 _3481_ _1712_ VPWR VGND sg13g2_nor2_1
X_7528_ _3267_ _3274_ _3276_ _3277_ _3278_ VPWR VGND sg13g2_nor4_1
X_7459_ _3211_ VPWR _3212_ VGND net1209 _3206_ sg13g2_o21ai_1
XFILLER_45_823 VPWR VGND sg13g2_decap_8
XFILLER_17_547 VPWR VGND sg13g2_fill_2
XFILLER_28_96 VPWR VGND sg13g2_fill_1
XFILLER_44_84 VPWR VGND sg13g2_fill_2
X_7729__293 VPWR VGND net293 sg13g2_tiehi
XFILLER_9_735 VPWR VGND sg13g2_fill_1
XFILLER_8_278 VPWR VGND sg13g2_fill_1
XFILLER_5_930 VPWR VGND sg13g2_decap_8
X_7736__286 VPWR VGND net286 sg13g2_tiehi
XFILLER_48_683 VPWR VGND sg13g2_decap_8
X_6830_ net1285 VPWR _2644_ VGND _2577_ _2643_ sg13g2_o21ai_1
XFILLER_39_1006 VPWR VGND sg13g2_decap_8
X_7882__128 VPWR VGND net128 sg13g2_tiehi
X_6761_ s0.data_out\[7\]\[6\] s0.data_out\[6\]\[6\] net1281 _2583_ VPWR VGND sg13g2_mux2_1
X_5712_ net1401 net1358 _1637_ VPWR VGND sg13g2_nor2b_1
X_6692_ net1176 _3518_ _2521_ VPWR VGND sg13g2_nor2_1
X_5643_ VGND VPWR _1453_ _1579_ _1580_ net1427 sg13g2_a21oi_1
X_5574_ net1415 _1508_ _1514_ VPWR VGND sg13g2_nor2_1
Xhold201 s0.data_out\[0\]\[0\] VPWR VGND net570 sg13g2_dlygate4sd3_1
X_4525_ _0569_ VPWR _0570_ VGND _0527_ _0529_ sg13g2_o21ai_1
X_7313_ _0067_ _3081_ _3082_ _3534_ net1585 VPWR VGND sg13g2_a22oi_1
Xhold223 _0199_ VPWR VGND net592 sg13g2_dlygate4sd3_1
Xhold212 _0042_ VPWR VGND net581 sg13g2_dlygate4sd3_1
Xhold234 s0.data_out\[14\]\[1\] VPWR VGND net603 sg13g2_dlygate4sd3_1
Xhold245 s0.data_out\[1\]\[3\] VPWR VGND net614 sg13g2_dlygate4sd3_1
X_4456_ net626 net637 net1543 _0501_ VPWR VGND sg13g2_mux2_1
Xhold278 s0.data_out\[19\]\[0\] VPWR VGND net647 sg13g2_dlygate4sd3_1
Xhold267 s0.was_valid_out\[16\][0] VPWR VGND net636 sg13g2_dlygate4sd3_1
Xhold256 _1946_ VPWR VGND net625 sg13g2_dlygate4sd3_1
X_7244_ _3016_ net1232 _3017_ _3018_ VPWR VGND sg13g2_a21o_1
X_4387_ s0.data_out\[26\]\[5\] s0.data_out\[25\]\[5\] net1540 _0444_ VPWR VGND sg13g2_mux2_1
X_7175_ VGND VPWR net1170 _2888_ _2959_ net1581 sg13g2_a21oi_1
Xhold289 _1824_ VPWR VGND net658 sg13g2_dlygate4sd3_1
X_6126_ net1371 net1330 _2015_ VPWR VGND sg13g2_nor2b_1
X_6057_ _0285_ _1951_ _1952_ _3484_ net1628 VPWR VGND sg13g2_a22oi_1
XFILLER_39_694 VPWR VGND sg13g2_fill_1
X_5008_ _1006_ net509 net1490 VPWR VGND sg13g2_nand2b_1
XFILLER_26_300 VPWR VGND sg13g2_decap_4
XFILLER_41_347 VPWR VGND sg13g2_fill_1
X_6959_ _0035_ _2759_ _2760_ _3519_ net1597 VPWR VGND sg13g2_a22oi_1
XFILLER_14_98 VPWR VGND sg13g2_fill_2
XFILLER_2_966 VPWR VGND sg13g2_decap_8
XFILLER_7_1004 VPWR VGND sg13g2_decap_8
XFILLER_17_311 VPWR VGND sg13g2_fill_2
XFILLER_18_867 VPWR VGND sg13g2_fill_2
XFILLER_13_572 VPWR VGND sg13g2_fill_2
X_4310_ _0119_ _0370_ _0371_ _3400_ net1575 VPWR VGND sg13g2_a22oi_1
X_5290_ net1619 _1182_ _1260_ VPWR VGND sg13g2_nor2_1
X_4241_ net472 net1563 _3605_ VPWR VGND sg13g2_nor2b_1
X_4172_ VGND VPWR _3415_ net1165 net4 _3546_ sg13g2_a21oi_1
X_7931_ net75 VGND VPWR _0065_ s0.data_out\[3\]\[1\] clknet_leaf_2_clk sg13g2_dfrbpq_2
XFILLER_35_130 VPWR VGND sg13g2_fill_1
XFILLER_24_826 VPWR VGND sg13g2_decap_8
X_7862_ net150 VGND VPWR _0340_ s0.data_out\[9\]\[4\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_23_347 VPWR VGND sg13g2_fill_1
X_7793_ net224 VGND VPWR _0271_ s0.data_out\[14\]\[2\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_6813_ _0019_ _2629_ _2630_ _3515_ net1598 VPWR VGND sg13g2_a22oi_1
X_6744_ _2566_ net1279 net796 VPWR VGND sg13g2_nand2_1
X_6675_ net1283 s0.data_out\[7\]\[0\] _2508_ VPWR VGND sg13g2_and2_1
XFILLER_31_380 VPWR VGND sg13g2_fill_1
X_5626_ VGND VPWR net1428 _1560_ _1563_ _1562_ sg13g2_a21oi_1
X_5557_ _1499_ VPWR _1500_ VGND net1745 net792 sg13g2_o21ai_1
X_4508_ _0553_ net1537 _0552_ VPWR VGND sg13g2_nand2b_1
X_5488_ _1435_ net1429 _1436_ _1437_ VPWR VGND sg13g2_a21o_1
X_4439_ _0485_ _0486_ _0487_ VPWR VGND sg13g2_nor2_1
X_7227_ net1228 net1356 _3001_ VPWR VGND sg13g2_nor2b_1
Xfanout1509 net1511 net1509 VPWR VGND sg13g2_buf_1
X_7158_ VGND VPWR _2944_ _2942_ net1658 sg13g2_or2_1
X_7089_ VGND VPWR _3361_ _2872_ _0048_ _2877_ sg13g2_a21oi_1
X_6109_ _1997_ VPWR _1998_ VGND net1373 _3489_ sg13g2_o21ai_1
XFILLER_18_119 VPWR VGND sg13g2_fill_1
XFILLER_42_645 VPWR VGND sg13g2_fill_2
XFILLER_41_122 VPWR VGND sg13g2_fill_1
XFILLER_15_859 VPWR VGND sg13g2_fill_1
XFILLER_41_144 VPWR VGND sg13g2_decap_4
XFILLER_6_568 VPWR VGND sg13g2_fill_1
XFILLER_29_1027 VPWR VGND sg13g2_fill_2
XFILLER_2_763 VPWR VGND sg13g2_decap_8
XFILLER_49_211 VPWR VGND sg13g2_fill_2
X_7733__289 VPWR VGND net289 sg13g2_tiehi
XFILLER_46_995 VPWR VGND sg13g2_decap_8
XFILLER_33_623 VPWR VGND sg13g2_decap_4
X_4790_ net1496 net530 _0807_ VPWR VGND sg13g2_and2_1
XFILLER_20_306 VPWR VGND sg13g2_fill_2
XFILLER_21_829 VPWR VGND sg13g2_fill_2
XFILLER_32_188 VPWR VGND sg13g2_fill_1
X_6460_ net1641 net1304 _2309_ VPWR VGND sg13g2_nor2b_1
X_6391_ VGND VPWR _2119_ _2248_ _2249_ net1323 sg13g2_a21oi_1
X_5411_ net1206 _3464_ _1369_ VPWR VGND sg13g2_nor2_1
X_7649__36 VPWR VGND net36 sg13g2_tiehi
X_5342_ s0.data_out\[17\]\[0\] s0.data_out\[18\]\[0\] net1454 _1303_ VPWR VGND sg13g2_mux2_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
X_5273_ _1245_ VPWR _1246_ VGND net1692 _1206_ sg13g2_o21ai_1
X_7012_ s0.data_out\[5\]\[6\] s0.data_out\[4\]\[6\] net1255 _2810_ VPWR VGND sg13g2_mux2_1
X_4224_ _3409_ _3385_ net1561 _3588_ VPWR VGND sg13g2_a21o_1
X_4155_ VPWR _3531_ net780 VGND sg13g2_inv_1
X_4086_ VPWR _3462_ net585 VGND sg13g2_inv_1
X_7914_ net94 VGND VPWR net401 s0.was_valid_out\[4\][0] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_7845_ net168 VGND VPWR _0323_ s0.shift_out\[10\][0] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_36_494 VPWR VGND sg13g2_decap_8
X_4988_ net1468 net1330 _0986_ VPWR VGND sg13g2_nor2b_1
X_7776_ net242 VGND VPWR _0254_ s0.valid_out\[15\][0] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_6727_ VGND VPWR net1282 _2546_ _2549_ _2548_ sg13g2_a21oi_1
X_6658_ net1286 net1339 _2492_ VPWR VGND sg13g2_nor2b_1
X_5609_ _1546_ s0.data_out\[15\]\[3\] net1432 VPWR VGND sg13g2_nand2b_1
X_6589_ net1641 net1291 _2426_ VPWR VGND sg13g2_nor2b_1
Xfanout1328 net1329 net1328 VPWR VGND sg13g2_buf_8
Xfanout1317 net1318 net1317 VPWR VGND sg13g2_buf_1
Xfanout1306 net1313 net1306 VPWR VGND sg13g2_buf_1
Xfanout1339 net1342 net1339 VPWR VGND sg13g2_buf_8
XFILLER_4_1018 VPWR VGND sg13g2_decap_8
XFILLER_47_759 VPWR VGND sg13g2_decap_8
XFILLER_43_921 VPWR VGND sg13g2_decap_8
X_7687__339 VPWR VGND net339 sg13g2_tiehi
XFILLER_27_461 VPWR VGND sg13g2_fill_1
XFILLER_15_623 VPWR VGND sg13g2_fill_1
XFILLER_43_998 VPWR VGND sg13g2_decap_8
X_7646__39 VPWR VGND net39 sg13g2_tiehi
XFILLER_42_1024 VPWR VGND sg13g2_decap_4
X_5960_ VGND VPWR net1378 _1859_ _1861_ _1860_ sg13g2_a21oi_1
X_5891_ _1804_ net1399 net582 VPWR VGND sg13g2_nand2_1
X_4911_ net1605 _0848_ _0918_ VPWR VGND sg13g2_nor2_1
X_7630_ net204 VGND VPWR _0108_ s0.module0.bubble clknet_leaf_11_clk sg13g2_dfrbpq_1
X_4842_ net1486 net1359 _0851_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_475 VPWR VGND sg13g2_fill_1
XFILLER_34_998 VPWR VGND sg13g2_decap_8
X_7561_ VGND VPWR net1200 _3260_ _3305_ net1587 sg13g2_a21oi_1
X_4773_ VGND VPWR _0789_ _0792_ _0794_ _0793_ sg13g2_a21oi_1
X_6512_ _2358_ net1303 net608 VPWR VGND sg13g2_nand2_1
X_7492_ _3242_ _3241_ net1686 _3220_ net1695 VPWR VGND sg13g2_a22oi_1
X_6443_ _2261_ _2295_ net1738 _2296_ VPWR VGND sg13g2_nand3_1
X_6374_ _2232_ net544 net1360 VPWR VGND sg13g2_nand2b_1
X_5325_ _1285_ VPWR _1286_ VGND net1443 _3461_ sg13g2_o21ai_1
X_5256_ net1450 net1341 _1229_ VPWR VGND sg13g2_nor2b_1
X_4207_ VGND VPWR net1564 _3417_ _3571_ _3570_ sg13g2_a21oi_1
X_5187_ _1164_ VPWR _1165_ VGND net1742 net784 sg13g2_o21ai_1
X_4138_ VPWR _3514_ net802 VGND sg13g2_inv_1
XFILLER_29_759 VPWR VGND sg13g2_fill_1
X_4069_ VPWR _3445_ net627 VGND sg13g2_inv_1
XFILLER_12_604 VPWR VGND sg13g2_fill_2
XFILLER_24_442 VPWR VGND sg13g2_fill_1
X_7828_ net186 VGND VPWR _0306_ s0.data_out\[11\]\[1\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_7759_ net261 VGND VPWR _0237_ s0.data_out\[17\]\[4\] clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_20_681 VPWR VGND sg13g2_fill_1
XFILLER_4_814 VPWR VGND sg13g2_fill_2
X_7693__332 VPWR VGND net332 sg13g2_tiehi
XFILLER_26_1019 VPWR VGND sg13g2_decap_8
X_7636__50 VPWR VGND net50 sg13g2_tiehi
Xfanout1169 _3411_ net1169 VPWR VGND sg13g2_buf_8
XFILLER_15_431 VPWR VGND sg13g2_fill_2
X_7878__133 VPWR VGND net133 sg13g2_tiehi
X_5110_ _1095_ _3392_ s0.data_out\[19\]\[3\] VPWR VGND sg13g2_nand2_1
X_6090_ VGND VPWR _1858_ _1978_ _1979_ net1376 sg13g2_a21oi_1
X_5041_ VPWR _0185_ _1036_ VGND sg13g2_inv_1
XFILLER_38_556 VPWR VGND sg13g2_fill_1
Xfanout1692 net1693 net1692 VPWR VGND sg13g2_buf_8
Xfanout1670 net1671 net1670 VPWR VGND sg13g2_buf_8
Xfanout1681 ui_in[4] net1681 VPWR VGND sg13g2_buf_8
X_6992_ _2790_ _2789_ net1260 VPWR VGND sg13g2_nand2b_1
X_5943_ _0276_ _1846_ _1847_ _3476_ net1629 VPWR VGND sg13g2_a22oi_1
X_5874_ net1395 net1336 _1787_ VPWR VGND sg13g2_nor2b_1
X_7613_ VGND VPWR _3351_ net1565 net382 sg13g2_or2_1
X_4825_ _0834_ net1491 s0.data_out\[21\]\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_21_456 VPWR VGND sg13g2_fill_1
XFILLER_21_489 VPWR VGND sg13g2_decap_4
X_7544_ _0089_ _3290_ _3291_ _3542_ net1583 VPWR VGND sg13g2_a22oi_1
X_4756_ _0777_ net1181 _0776_ VPWR VGND sg13g2_nand2_1
X_7475_ _3223_ net1208 _3224_ _3225_ VPWR VGND sg13g2_a21o_1
X_4687_ VGND VPWR net1634 net1503 _0711_ _0710_ sg13g2_a21oi_1
X_6426_ _2225_ _2282_ net1738 _2283_ VPWR VGND sg13g2_nand3_1
XFILLER_1_817 VPWR VGND sg13g2_decap_8
X_6357_ _2214_ VPWR _2215_ VGND net1315 _3498_ sg13g2_o21ai_1
X_5308_ _0215_ _1272_ _1273_ _3452_ net1617 VPWR VGND sg13g2_a22oi_1
X_6288_ _2163_ VPWR _2164_ VGND net1740 net786 sg13g2_o21ai_1
X_5239_ _1210_ net1448 _1211_ _1212_ VPWR VGND sg13g2_a21o_1
X_7633__53 VPWR VGND net53 sg13g2_tiehi
XFILLER_17_76 VPWR VGND sg13g2_fill_2
XFILLER_0_894 VPWR VGND sg13g2_decap_8
Xhold5 s0.genblk1\[24\].modules.bubble VPWR VGND net374 sg13g2_dlygate4sd3_1
XFILLER_48_865 VPWR VGND sg13g2_decap_8
XFILLER_47_397 VPWR VGND sg13g2_fill_1
XFILLER_43_581 VPWR VGND sg13g2_fill_2
X_4610_ VPWR VGND net1688 _0635_ _0642_ net1696 _0643_ _0618_ sg13g2_a221oi_1
X_5590_ s0.data_out\[16\]\[1\] s0.data_out\[15\]\[1\] net1419 _1527_ VPWR VGND sg13g2_mux2_1
XFILLER_8_961 VPWR VGND sg13g2_decap_8
X_4541_ _0514_ _0582_ net1725 _0583_ VPWR VGND sg13g2_nand3_1
Xhold405 s0.data_out\[25\]\[5\] VPWR VGND net774 sg13g2_dlygate4sd3_1
Xhold416 s0.shift_out\[25\][0] VPWR VGND net785 sg13g2_dlygate4sd3_1
X_4472_ _0517_ net1571 _0515_ VPWR VGND sg13g2_xnor2_1
X_7260_ net1231 net1329 _3034_ VPWR VGND sg13g2_nor2b_1
Xhold427 s0.data_out\[6\]\[3\] VPWR VGND net796 sg13g2_dlygate4sd3_1
Xhold438 s0.data_out\[6\]\[5\] VPWR VGND net807 sg13g2_dlygate4sd3_1
X_6211_ s0.data_out\[11\]\[2\] s0.data_out\[10\]\[2\] net1360 _2088_ VPWR VGND sg13g2_mux2_1
X_7191_ _2971_ VPWR _2972_ VGND net1723 net670 sg13g2_o21ai_1
Xhold449 s0.data_out\[8\]\[4\] VPWR VGND net818 sg13g2_dlygate4sd3_1
X_6142_ _2031_ net1675 _2030_ VPWR VGND sg13g2_nand2_1
XFILLER_31_0 VPWR VGND sg13g2_fill_1
X_6073_ _1963_ _1964_ _1965_ VPWR VGND sg13g2_nor2_1
X_5024_ _1017_ _1021_ _1009_ _1022_ VPWR VGND sg13g2_nand3_1
XFILLER_39_898 VPWR VGND sg13g2_fill_2
X_6975_ _2771_ net1250 _2772_ _2773_ VPWR VGND sg13g2_a21o_1
X_5926_ VGND VPWR net1394 net574 _1834_ _1799_ sg13g2_a21oi_1
XFILLER_34_581 VPWR VGND sg13g2_fill_2
X_5857_ _1769_ VPWR _1770_ VGND net1400 _3479_ sg13g2_o21ai_1
X_4808_ net1493 net558 _0821_ VPWR VGND sg13g2_and2_1
X_5788_ VPWR _0257_ _1711_ VGND sg13g2_inv_1
X_7527_ VGND VPWR _3261_ _3265_ _3277_ net1669 sg13g2_a21oi_1
X_4739_ _0760_ net1505 net552 VPWR VGND sg13g2_nand2_1
X_7458_ net1202 VPWR _3211_ VGND net507 net1224 sg13g2_o21ai_1
X_6409_ _2267_ s0.data_out\[9\]\[5\] net1362 VPWR VGND sg13g2_nand2b_1
XFILLER_1_614 VPWR VGND sg13g2_decap_8
X_7389_ _3151_ _3150_ net1648 _3144_ net1659 VPWR VGND sg13g2_a22oi_1
XFILLER_48_106 VPWR VGND sg13g2_fill_2
X_7868__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_28_64 VPWR VGND sg13g2_fill_2
XFILLER_17_515 VPWR VGND sg13g2_fill_1
XFILLER_45_879 VPWR VGND sg13g2_decap_8
XFILLER_8_224 VPWR VGND sg13g2_fill_1
X_7875__136 VPWR VGND net136 sg13g2_tiehi
XFILLER_4_441 VPWR VGND sg13g2_fill_2
XFILLER_5_986 VPWR VGND sg13g2_decap_8
XFILLER_4_496 VPWR VGND sg13g2_fill_2
XFILLER_0_691 VPWR VGND sg13g2_decap_8
XFILLER_48_662 VPWR VGND sg13g2_decap_8
XFILLER_36_868 VPWR VGND sg13g2_fill_2
X_6760_ _2582_ net1280 net719 VPWR VGND sg13g2_nand2_1
XFILLER_44_890 VPWR VGND sg13g2_decap_8
X_5711_ _1636_ net1197 _1635_ VPWR VGND sg13g2_nand2_1
X_6691_ _0007_ _2519_ _2520_ _3511_ net1599 VPWR VGND sg13g2_a22oi_1
X_5642_ _1579_ s0.data_out\[15\]\[5\] net1433 VPWR VGND sg13g2_nand2b_1
XFILLER_31_584 VPWR VGND sg13g2_fill_1
X_5573_ VGND VPWR _1513_ _1512_ _1510_ sg13g2_or2_1
Xhold202 s0.valid_out\[0\][0] VPWR VGND net571 sg13g2_dlygate4sd3_1
X_7312_ net1585 _3020_ _3082_ VPWR VGND sg13g2_nor2_1
X_4524_ _0548_ _0565_ _0566_ _0568_ _0569_ VPWR VGND sg13g2_nor4_1
Xhold213 s0.data_out\[13\]\[5\] VPWR VGND net582 sg13g2_dlygate4sd3_1
Xhold235 s0.data_out\[3\]\[7\] VPWR VGND net604 sg13g2_dlygate4sd3_1
Xhold224 s0.data_out\[7\]\[3\] VPWR VGND net593 sg13g2_dlygate4sd3_1
Xhold246 _3299_ VPWR VGND net615 sg13g2_dlygate4sd3_1
X_7243_ net1232 net1167 _3017_ VPWR VGND sg13g2_nor2_1
X_4455_ VGND VPWR net1538 _0497_ _0500_ _0499_ sg13g2_a21oi_1
Xhold257 s0.data_out\[24\]\[0\] VPWR VGND net626 sg13g2_dlygate4sd3_1
Xhold268 s0.data_out\[25\]\[0\] VPWR VGND net637 sg13g2_dlygate4sd3_1
X_4386_ _0443_ net1542 s0.data_out\[25\]\[5\] VPWR VGND sg13g2_nand2_1
X_7174_ VGND VPWR net1240 s0.data_out\[3\]\[1\] _2958_ _2885_ sg13g2_a21oi_1
Xhold279 _1254_ VPWR VGND net648 sg13g2_dlygate4sd3_1
X_6125_ s0.data_out\[12\]\[7\] s0.data_out\[11\]\[7\] net1375 _2014_ VPWR VGND sg13g2_mux2_1
X_6056_ net1628 _1897_ _1952_ VPWR VGND sg13g2_nor2_1
XFILLER_22_1022 VPWR VGND sg13g2_decap_8
X_5007_ _1003_ net1468 _1004_ _1005_ VPWR VGND sg13g2_a21o_1
XFILLER_26_356 VPWR VGND sg13g2_fill_1
XFILLER_27_868 VPWR VGND sg13g2_fill_2
XFILLER_42_827 VPWR VGND sg13g2_fill_1
X_6958_ net1597 _2701_ _2760_ VPWR VGND sg13g2_nor2_1
X_6889_ _2697_ net1264 _2698_ _2699_ VPWR VGND sg13g2_a21o_1
X_5909_ VGND VPWR net1390 s0.data_out\[13\]\[0\] _1821_ _1762_ sg13g2_a21oi_1
XFILLER_6_717 VPWR VGND sg13g2_fill_2
XFILLER_5_238 VPWR VGND sg13g2_fill_2
XFILLER_2_945 VPWR VGND sg13g2_decap_8
XFILLER_1_433 VPWR VGND sg13g2_fill_2
XFILLER_39_74 VPWR VGND sg13g2_fill_2
XFILLER_39_63 VPWR VGND sg13g2_fill_2
XFILLER_18_835 VPWR VGND sg13g2_fill_2
XFILLER_29_150 VPWR VGND sg13g2_fill_2
XFILLER_9_566 VPWR VGND sg13g2_fill_2
X_4240_ VGND VPWR net1558 _3603_ _3604_ _3599_ sg13g2_a21oi_1
X_4171_ s0.data_out\[27\]\[1\] net1165 _3546_ VPWR VGND sg13g2_nor2_1
X_7930_ net76 VGND VPWR _0064_ s0.data_out\[3\]\[0\] clknet_leaf_2_clk sg13g2_dfrbpq_2
X_7861_ net151 VGND VPWR _0339_ s0.data_out\[9\]\[3\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_6812_ net1598 _2571_ _2630_ VPWR VGND sg13g2_nor2_1
X_7792_ net225 VGND VPWR _0270_ s0.data_out\[14\]\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_6743_ _2550_ VPWR _2565_ VGND net1703 _2557_ sg13g2_o21ai_1
X_6674_ VGND VPWR _2503_ _2506_ _0003_ _2507_ sg13g2_a21oi_1
X_5625_ VGND VPWR _1441_ _1561_ _1562_ net1428 sg13g2_a21oi_1
X_5556_ _1498_ VPWR _1499_ VGND net1207 _1497_ sg13g2_o21ai_1
X_4507_ VGND VPWR net1519 _0550_ _0552_ _0551_ sg13g2_a21oi_1
X_5487_ net1429 net1330 _1436_ VPWR VGND sg13g2_nor2b_1
X_4438_ net1641 _3389_ _0486_ VPWR VGND sg13g2_nor2_1
X_7226_ s0.data_out\[3\]\[0\] s0.data_out\[2\]\[0\] net1235 _3000_ VPWR VGND sg13g2_mux2_1
X_4369_ net1534 net1328 _0426_ VPWR VGND sg13g2_nor2b_1
X_7157_ _2943_ _2942_ net1659 _2936_ net1647 VPWR VGND sg13g2_a22oi_1
X_7088_ net1716 VPWR _2877_ VGND _2874_ _2876_ sg13g2_o21ai_1
X_6108_ _1997_ net1372 s0.data_out\[11\]\[3\] VPWR VGND sg13g2_nand2_1
X_6039_ VPWR _0281_ _1938_ VGND sg13g2_inv_1
XFILLER_42_602 VPWR VGND sg13g2_fill_2
XFILLER_26_142 VPWR VGND sg13g2_fill_1
XFILLER_27_687 VPWR VGND sg13g2_fill_1
XFILLER_25_76 VPWR VGND sg13g2_decap_8
XFILLER_30_819 VPWR VGND sg13g2_decap_8
X_7726__297 VPWR VGND net297 sg13g2_tiehi
XFILLER_22_392 VPWR VGND sg13g2_fill_1
X_7658__26 VPWR VGND net26 sg13g2_tiehi
XFILLER_29_1006 VPWR VGND sg13g2_decap_8
XFILLER_2_742 VPWR VGND sg13g2_decap_8
X_7872__139 VPWR VGND net139 sg13g2_tiehi
XFILLER_46_974 VPWR VGND sg13g2_decap_8
XFILLER_45_451 VPWR VGND sg13g2_fill_1
XFILLER_18_698 VPWR VGND sg13g2_fill_2
XFILLER_21_819 VPWR VGND sg13g2_fill_1
XFILLER_9_330 VPWR VGND sg13g2_decap_4
XFILLER_9_352 VPWR VGND sg13g2_fill_2
XFILLER_12_1010 VPWR VGND sg13g2_decap_8
X_6390_ _2248_ net832 net1362 VPWR VGND sg13g2_nand2b_1
X_5410_ VPWR _0222_ net809 VGND sg13g2_inv_1
X_5341_ VGND VPWR net1436 _1300_ _1302_ _1301_ sg13g2_a21oi_1
X_5272_ _1233_ _1231_ net1674 _1245_ VPWR VGND sg13g2_a21o_1
X_7011_ _2809_ net1253 net536 VPWR VGND sg13g2_nand2_1
X_4223_ VGND VPWR _3577_ _3586_ _3587_ _3569_ sg13g2_a21oi_1
X_4154_ VPWR _3530_ net752 VGND sg13g2_inv_1
X_4085_ VPWR _3461_ s0.data_out\[18\]\[2\] VGND sg13g2_inv_1
X_7913_ net95 VGND VPWR net567 s0.data_out\[5\]\[7\] clknet_leaf_6_clk sg13g2_dfrbpq_2
XFILLER_37_996 VPWR VGND sg13g2_decap_8
X_7844_ net169 VGND VPWR _0322_ s0.data_new_delayed\[7\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_36_484 VPWR VGND sg13g2_fill_2
X_7775_ net244 VGND VPWR net406 s0.was_valid_out\[15\][0] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_4987_ s0.data_out\[21\]\[7\] s0.data_out\[20\]\[7\] net1478 _0985_ VPWR VGND sg13g2_mux2_1
X_6726_ VGND VPWR _2435_ _2547_ _2548_ net1282 sg13g2_a21oi_1
X_6657_ s0.data_out\[8\]\[5\] s0.data_out\[7\]\[5\] net1292 _2491_ VPWR VGND sg13g2_mux2_1
X_6588_ net1297 VPWR _2425_ VGND net1641 net1287 sg13g2_o21ai_1
X_5608_ _1543_ net1413 _1544_ _1545_ VPWR VGND sg13g2_a21o_1
XFILLER_3_517 VPWR VGND sg13g2_fill_1
X_5539_ _0234_ _1484_ _1485_ _3465_ net1619 VPWR VGND sg13g2_a22oi_1
XFILLER_11_89 VPWR VGND sg13g2_fill_2
Xfanout1318 s0.valid_out\[9\][0] net1318 VPWR VGND sg13g2_buf_2
Xfanout1329 net1332 net1329 VPWR VGND sg13g2_buf_8
X_7209_ VGND VPWR net1191 _2869_ _2986_ _2985_ sg13g2_a21oi_1
Xfanout1307 net1308 net1307 VPWR VGND sg13g2_buf_2
XFILLER_47_738 VPWR VGND sg13g2_decap_8
X_7732__290 VPWR VGND net290 sg13g2_tiehi
XFILLER_27_451 VPWR VGND sg13g2_fill_2
XFILLER_28_985 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_fill_2
XFILLER_36_75 VPWR VGND sg13g2_fill_2
XFILLER_15_613 VPWR VGND sg13g2_fill_1
XFILLER_43_977 VPWR VGND sg13g2_decap_8
XFILLER_42_498 VPWR VGND sg13g2_fill_1
XFILLER_42_476 VPWR VGND sg13g2_fill_1
XFILLER_14_156 VPWR VGND sg13g2_fill_1
XFILLER_11_863 VPWR VGND sg13g2_fill_1
XFILLER_42_1003 VPWR VGND sg13g2_decap_8
XFILLER_38_738 VPWR VGND sg13g2_decap_8
XFILLER_46_793 VPWR VGND sg13g2_decap_8
X_5890_ _1802_ VPWR _1803_ VGND _3381_ _1800_ sg13g2_o21ai_1
X_4910_ net1501 VPWR _0917_ VGND _0845_ _0916_ sg13g2_o21ai_1
XFILLER_33_410 VPWR VGND sg13g2_fill_2
XFILLER_34_933 VPWR VGND sg13g2_fill_2
X_4841_ s0.data_out\[22\]\[0\] s0.data_out\[21\]\[0\] net1491 _0850_ VPWR VGND sg13g2_mux2_1
XFILLER_34_977 VPWR VGND sg13g2_decap_8
XFILLER_33_487 VPWR VGND sg13g2_fill_1
X_7560_ VGND VPWR net1213 net439 _3304_ _3263_ sg13g2_a21oi_1
X_4772_ _0712_ VPWR _0793_ VGND _0767_ _0769_ sg13g2_o21ai_1
X_6511_ VGND VPWR net1309 _2354_ _2357_ _2356_ sg13g2_a21oi_1
X_7491_ VGND VPWR net1200 _3236_ _3241_ _3240_ sg13g2_a21oi_1
X_6442_ net1320 VPWR _2295_ VGND _2257_ _2294_ sg13g2_o21ai_1
X_6373_ _2229_ net1308 _2230_ _2231_ VPWR VGND sg13g2_a21o_1
X_5324_ _1285_ net1443 s0.data_out\[17\]\[2\] VPWR VGND sg13g2_nand2_1
X_5255_ s0.data_out\[19\]\[5\] s0.data_out\[18\]\[5\] net1455 _1228_ VPWR VGND sg13g2_mux2_1
X_7645__40 VPWR VGND net40 sg13g2_tiehi
X_4206_ _3386_ VPWR _3570_ VGND net1564 s0.data_out\[26\]\[1\] sg13g2_o21ai_1
X_5186_ _1163_ net1742 _1164_ VPWR VGND _1105_ sg13g2_nand3b_1
X_4137_ VPWR _3513_ net649 VGND sg13g2_inv_1
X_4068_ _3444_ s0.data_out\[21\]\[2\] VPWR VGND sg13g2_inv_2
X_7686__340 VPWR VGND net340 sg13g2_tiehi
XFILLER_25_922 VPWR VGND sg13g2_fill_2
XFILLER_36_281 VPWR VGND sg13g2_fill_1
X_7827_ net187 VGND VPWR _0305_ s0.data_out\[11\]\[0\] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_25_988 VPWR VGND sg13g2_decap_8
XFILLER_40_969 VPWR VGND sg13g2_decap_8
X_7758_ net262 VGND VPWR net543 s0.data_out\[17\]\[3\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_6709_ _2534_ net1634 net1281 VPWR VGND sg13g2_nand2_1
X_7689_ net337 VGND VPWR _0167_ s0.data_out\[23\]\[6\] clknet_leaf_42_clk sg13g2_dfrbpq_2
XFILLER_47_579 VPWR VGND sg13g2_fill_2
XFILLER_47_557 VPWR VGND sg13g2_fill_2
XFILLER_16_922 VPWR VGND sg13g2_fill_2
XFILLER_16_988 VPWR VGND sg13g2_decap_8
XFILLER_15_498 VPWR VGND sg13g2_fill_2
XFILLER_30_446 VPWR VGND sg13g2_decap_4
XFILLER_11_660 VPWR VGND sg13g2_fill_1
X_5040_ _1035_ VPWR _1036_ VGND net1734 net629 sg13g2_o21ai_1
XFILLER_38_502 VPWR VGND sg13g2_decap_8
Xfanout1660 net1662 net1660 VPWR VGND sg13g2_buf_8
Xfanout1671 net1672 net1671 VPWR VGND sg13g2_buf_8
Xfanout1682 net1685 net1682 VPWR VGND sg13g2_buf_8
Xfanout1693 net1694 net1693 VPWR VGND sg13g2_buf_8
XFILLER_19_760 VPWR VGND sg13g2_fill_2
X_6991_ s0.data_out\[4\]\[0\] s0.data_out\[5\]\[0\] net1266 _2789_ VPWR VGND sg13g2_mux2_1
XFILLER_26_719 VPWR VGND sg13g2_fill_1
X_5942_ net1631 _1783_ _1847_ VPWR VGND sg13g2_nor2_1
XFILLER_18_281 VPWR VGND sg13g2_fill_2
XFILLER_22_903 VPWR VGND sg13g2_fill_1
X_5873_ s0.data_out\[14\]\[6\] s0.data_out\[13\]\[6\] net1400 _1786_ VPWR VGND sg13g2_mux2_1
X_7612_ VGND VPWR net1648 _3321_ _3350_ net1640 sg13g2_a21oi_1
X_4824_ net1736 net389 _0171_ VPWR VGND sg13g2_and2_1
X_4755_ s0.data_out\[22\]\[5\] s0.data_out\[23\]\[5\] net1516 _0776_ VPWR VGND sg13g2_mux2_1
X_7543_ net1583 _3222_ _3291_ VPWR VGND sg13g2_nor2_1
X_4686_ net1513 VPWR _0710_ VGND net1641 net1493 sg13g2_o21ai_1
X_7474_ net1208 net1352 _3224_ VPWR VGND sg13g2_nor2b_1
X_6425_ net1319 VPWR _2282_ VGND _2221_ _2281_ sg13g2_o21ai_1
X_6356_ _2214_ net1314 net549 VPWR VGND sg13g2_nand2_1
X_5307_ net1617 _1214_ _1273_ VPWR VGND sg13g2_nor2_1
X_6287_ _2107_ _2162_ net1740 _2163_ VPWR VGND sg13g2_nand3_1
X_5238_ net1448 net1336 _1211_ VPWR VGND sg13g2_nor2b_1
X_5169_ net1475 VPWR _1151_ VGND _1070_ _1150_ sg13g2_o21ai_1
XFILLER_33_32 VPWR VGND sg13g2_fill_2
XFILLER_21_991 VPWR VGND sg13g2_decap_8
XFILLER_32_1024 VPWR VGND sg13g2_decap_4
XFILLER_3_177 VPWR VGND sg13g2_fill_2
XFILLER_3_188 VPWR VGND sg13g2_fill_2
XFILLER_0_873 VPWR VGND sg13g2_decap_8
XFILLER_48_844 VPWR VGND sg13g2_decap_8
Xhold6 s0.genblk1\[23\].modules.bubble VPWR VGND net375 sg13g2_dlygate4sd3_1
XFILLER_43_571 VPWR VGND sg13g2_fill_1
XFILLER_30_276 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_10_clk clknet_3_2__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_4540_ net1538 VPWR _0582_ VGND _0509_ _0581_ sg13g2_o21ai_1
Xhold406 s0.data_out\[25\]\[6\] VPWR VGND net775 sg13g2_dlygate4sd3_1
X_4471_ VGND VPWR _0516_ _0515_ net1571 sg13g2_or2_1
Xhold417 s0.data_out\[11\]\[0\] VPWR VGND net786 sg13g2_dlygate4sd3_1
Xhold428 s0.data_out\[21\]\[5\] VPWR VGND net797 sg13g2_dlygate4sd3_1
Xhold439 s0.data_out\[18\]\[1\] VPWR VGND net808 sg13g2_dlygate4sd3_1
X_6210_ _2087_ net1360 net523 VPWR VGND sg13g2_nand2_1
X_7190_ _2970_ VPWR _2971_ VGND net1173 _2969_ sg13g2_o21ai_1
X_6141_ VGND VPWR net1379 _2027_ _2030_ _2029_ sg13g2_a21oi_1
X_6072_ net1643 net1375 _1964_ VPWR VGND sg13g2_nor2b_1
X_5023_ _1018_ _1019_ _1020_ _1021_ VPWR VGND sg13g2_nor3_1
XFILLER_39_855 VPWR VGND sg13g2_fill_1
XFILLER_38_343 VPWR VGND sg13g2_fill_2
Xfanout1490 s0.valid_out\[21\][0] net1490 VPWR VGND sg13g2_buf_8
XFILLER_26_516 VPWR VGND sg13g2_fill_2
X_6974_ net1250 net1349 _2772_ VPWR VGND sg13g2_nor2b_1
X_5925_ _0272_ _1832_ _1833_ _3479_ net1626 VPWR VGND sg13g2_a22oi_1
X_5856_ _1769_ net1398 net757 VPWR VGND sg13g2_nand2_1
X_7683__343 VPWR VGND net343 sg13g2_tiehi
X_4807_ _0167_ _0819_ _0820_ _3433_ net1593 VPWR VGND sg13g2_a22oi_1
XFILLER_21_276 VPWR VGND sg13g2_fill_1
XFILLER_21_287 VPWR VGND sg13g2_fill_2
X_5787_ _1710_ VPWR _1711_ VGND net1747 net679 sg13g2_o21ai_1
X_7526_ _3275_ VPWR _3276_ VGND net1686 _3241_ sg13g2_o21ai_1
X_4738_ VGND VPWR net1512 _0756_ _0759_ _0758_ sg13g2_a21oi_1
X_7457_ VGND VPWR _3210_ net1214 net507 sg13g2_or2_1
X_4669_ _0152_ _0696_ _0697_ _3429_ net1589 VPWR VGND sg13g2_a22oi_1
X_6408_ _2264_ net1312 _2265_ _2266_ VPWR VGND sg13g2_a21o_1
X_7388_ VGND VPWR net1230 _3147_ _3150_ _3149_ sg13g2_a21oi_1
XFILLER_1_648 VPWR VGND sg13g2_decap_4
X_6339_ _2201_ VPWR _0318_ VGND net1637 net1167 sg13g2_o21ai_1
XFILLER_49_619 VPWR VGND sg13g2_decap_8
X_7690__336 VPWR VGND net336 sg13g2_tiehi
XFILLER_28_54 VPWR VGND sg13g2_fill_2
XFILLER_45_858 VPWR VGND sg13g2_decap_8
XFILLER_17_549 VPWR VGND sg13g2_fill_1
XFILLER_44_31 VPWR VGND sg13g2_fill_2
X_7909__99 VPWR VGND net99 sg13g2_tiehi
XFILLER_8_236 VPWR VGND sg13g2_fill_1
XFILLER_12_276 VPWR VGND sg13g2_fill_2
XFILLER_12_287 VPWR VGND sg13g2_fill_2
XFILLER_8_269 VPWR VGND sg13g2_fill_1
XFILLER_8_258 VPWR VGND sg13g2_decap_8
XFILLER_5_965 VPWR VGND sg13g2_decap_8
XFILLER_0_670 VPWR VGND sg13g2_decap_8
XFILLER_48_641 VPWR VGND sg13g2_decap_8
X_5710_ s0.data_out\[14\]\[0\] s0.data_out\[15\]\[0\] net1419 _1635_ VPWR VGND sg13g2_mux2_1
X_6690_ net1599 _2464_ _2520_ VPWR VGND sg13g2_nor2_1
XFILLER_31_530 VPWR VGND sg13g2_fill_2
X_5641_ _1576_ net1415 _1577_ _1578_ VPWR VGND sg13g2_a21o_1
X_5572_ net405 net1421 _1512_ VPWR VGND sg13g2_nor2_1
X_7311_ net1243 VPWR _3081_ VGND _3017_ _3080_ sg13g2_o21ai_1
X_4523_ VGND VPWR _0561_ _0563_ _0568_ net1679 sg13g2_a21oi_1
Xhold214 _0286_ VPWR VGND net583 sg13g2_dlygate4sd3_1
Xhold203 s0.data_out\[27\]\[0\] VPWR VGND net572 sg13g2_dlygate4sd3_1
Xhold225 _0019_ VPWR VGND net594 sg13g2_dlygate4sd3_1
X_7242_ _3015_ VPWR _3016_ VGND net1237 _3534_ sg13g2_o21ai_1
Xhold258 s0.data_out\[20\]\[7\] VPWR VGND net627 sg13g2_dlygate4sd3_1
X_4454_ VGND VPWR _0393_ _0498_ _0499_ net1538 sg13g2_a21oi_1
Xhold269 _0137_ VPWR VGND net638 sg13g2_dlygate4sd3_1
Xhold236 _0071_ VPWR VGND net605 sg13g2_dlygate4sd3_1
Xhold247 s0.data_out\[3\]\[4\] VPWR VGND net616 sg13g2_dlygate4sd3_1
X_4385_ VGND VPWR net1550 _0439_ _0442_ _0441_ sg13g2_a21oi_1
X_7173_ VPWR _0052_ net782 VGND sg13g2_inv_1
X_6124_ _2013_ net1374 net586 VPWR VGND sg13g2_nand2_1
X_6055_ net1392 VPWR _1951_ VGND _1894_ _1950_ sg13g2_o21ai_1
X_5006_ net1468 net1340 _1004_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_1001 VPWR VGND sg13g2_decap_8
X_6957_ net1274 VPWR _2759_ VGND _2698_ _2758_ sg13g2_o21ai_1
X_6888_ net1264 net1328 _2698_ VPWR VGND sg13g2_nor2b_1
X_5908_ VGND VPWR _1818_ _1819_ _0268_ _1820_ sg13g2_a21oi_1
XFILLER_22_563 VPWR VGND sg13g2_fill_1
X_5839_ VGND VPWR net1402 _1749_ _1752_ _1751_ sg13g2_a21oi_1
X_7509_ _3257_ _3258_ _3256_ _3259_ VPWR VGND sg13g2_nand3_1
XFILLER_2_924 VPWR VGND sg13g2_decap_8
XFILLER_49_438 VPWR VGND sg13g2_fill_1
XFILLER_17_313 VPWR VGND sg13g2_fill_1
XFILLER_29_195 VPWR VGND sg13g2_decap_4
XFILLER_40_360 VPWR VGND sg13g2_fill_2
XFILLER_45_1012 VPWR VGND sg13g2_decap_8
X_4170_ VGND VPWR net1570 net1165 net3 _3545_ sg13g2_a21oi_1
XFILLER_49_983 VPWR VGND sg13g2_decap_8
X_7860_ net152 VGND VPWR net486 s0.data_out\[9\]\[2\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_6811_ net1284 VPWR _2629_ VGND _2568_ _2628_ sg13g2_o21ai_1
X_7791_ net226 VGND VPWR _0269_ s0.data_out\[14\]\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_6742_ VPWR VGND _2563_ net1710 _2561_ net1703 _2564_ _2557_ sg13g2_a221oi_1
X_6673_ VGND VPWR _2507_ net1566 net376 sg13g2_or2_1
X_7680__346 VPWR VGND net346 sg13g2_tiehi
XFILLER_32_883 VPWR VGND sg13g2_fill_1
X_5624_ _1561_ s0.data_out\[15\]\[6\] net1434 VPWR VGND sg13g2_nand2b_1
X_5555_ VGND VPWR net1207 _1458_ _1498_ net1623 sg13g2_a21oi_1
X_7858__154 VPWR VGND net154 sg13g2_tiehi
X_4506_ net1519 net1338 _0551_ VPWR VGND sg13g2_nor2b_1
X_5486_ s0.data_out\[17\]\[7\] s0.data_out\[16\]\[7\] net1433 _1435_ VPWR VGND sg13g2_mux2_1
X_4437_ net1537 VPWR _0485_ VGND net1641 net1519 sg13g2_o21ai_1
X_7225_ _3415_ _2998_ _2999_ VPWR VGND sg13g2_nor2_1
X_7156_ VGND VPWR net1248 _2939_ _2942_ _2941_ sg13g2_a21oi_1
X_4368_ s0.data_out\[26\]\[7\] s0.data_out\[25\]\[7\] net1540 _0425_ VPWR VGND sg13g2_mux2_1
X_6107_ VPWR VGND _1994_ net1712 _1992_ net1707 _1996_ _1988_ sg13g2_a221oi_1
X_4299_ net1545 s0.data_out\[26\]\[4\] _0363_ VPWR VGND sg13g2_and2_1
X_7087_ _2876_ _2873_ _2875_ VPWR VGND sg13g2_nand2_1
XFILLER_46_408 VPWR VGND sg13g2_fill_2
X_6038_ _1937_ VPWR _1938_ VGND net1740 net732 sg13g2_o21ai_1
X_7865__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_42_647 VPWR VGND sg13g2_fill_1
XFILLER_26_198 VPWR VGND sg13g2_fill_2
XFILLER_25_55 VPWR VGND sg13g2_decap_4
XFILLER_2_798 VPWR VGND sg13g2_decap_8
XFILLER_46_953 VPWR VGND sg13g2_decap_8
X_5340_ net1436 net1358 _1301_ VPWR VGND sg13g2_nor2b_1
X_5271_ net1683 _1241_ _1244_ VPWR VGND sg13g2_nor2_1
X_4222_ _3585_ VPWR _3586_ VGND net1701 _3576_ sg13g2_o21ai_1
X_7010_ VGND VPWR net1259 _2805_ _2808_ _2807_ sg13g2_a21oi_1
X_4153_ VPWR _3529_ net580 VGND sg13g2_inv_1
X_4084_ VPWR _3460_ net487 VGND sg13g2_inv_1
XFILLER_49_780 VPWR VGND sg13g2_decap_8
X_7912_ net96 VGND VPWR _0046_ s0.data_out\[5\]\[6\] clknet_leaf_3_clk sg13g2_dfrbpq_2
XFILLER_37_975 VPWR VGND sg13g2_decap_8
X_7843_ net170 VGND VPWR _0321_ s0.data_new_delayed\[6\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_4986_ _0984_ net1480 net627 VPWR VGND sg13g2_nand2_1
XFILLER_23_146 VPWR VGND sg13g2_fill_1
X_7774_ net245 VGND VPWR net528 s0.data_out\[16\]\[7\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_11_308 VPWR VGND sg13g2_fill_2
X_6725_ _2547_ net532 net1289 VPWR VGND sg13g2_nand2b_1
X_6656_ VGND VPWR net1296 _2487_ _2490_ _2489_ sg13g2_a21oi_1
X_6587_ _0343_ _2423_ _2424_ _3503_ net1615 VPWR VGND sg13g2_a22oi_1
X_5607_ net1413 s0.data_new_delayed\[3\] _1544_ VPWR VGND sg13g2_nor2b_1
X_5538_ net1620 _1404_ _1485_ VPWR VGND sg13g2_nor2_1
X_5469_ _1418_ net1206 _1417_ VPWR VGND sg13g2_nand2_1
X_7871__140 VPWR VGND net140 sg13g2_tiehi
X_7208_ _2983_ _2984_ _2985_ VPWR VGND sg13g2_nor2_1
Xfanout1319 net1320 net1319 VPWR VGND sg13g2_buf_8
Xfanout1308 net1313 net1308 VPWR VGND sg13g2_buf_8
X_7139_ _2925_ net1173 _2924_ VPWR VGND sg13g2_nand2_1
XFILLER_47_717 VPWR VGND sg13g2_decap_8
XFILLER_28_920 VPWR VGND sg13g2_fill_1
XFILLER_15_603 VPWR VGND sg13g2_fill_1
XFILLER_43_956 VPWR VGND sg13g2_decap_8
XFILLER_35_1011 VPWR VGND sg13g2_decap_8
XFILLER_10_352 VPWR VGND sg13g2_decap_4
XFILLER_10_363 VPWR VGND sg13g2_decap_8
XFILLER_19_931 VPWR VGND sg13g2_fill_1
XFILLER_18_452 VPWR VGND sg13g2_decap_4
XFILLER_19_986 VPWR VGND sg13g2_decap_8
XFILLER_46_772 VPWR VGND sg13g2_decap_8
X_4840_ VGND VPWR net1500 _0846_ _0849_ _0848_ sg13g2_a21oi_1
X_7972__67 VPWR VGND net67 sg13g2_tiehi
X_6510_ VGND VPWR _2237_ _2355_ _2356_ net1309 sg13g2_a21oi_1
X_4771_ VGND VPWR _0778_ _0785_ _0792_ _0770_ sg13g2_a21oi_1
X_7490_ net1200 _3239_ _3240_ VPWR VGND sg13g2_nor2_1
X_6441_ net1308 s0.data_out\[9\]\[4\] _2294_ VPWR VGND sg13g2_and2_1
X_6372_ net1308 net1168 _2230_ VPWR VGND sg13g2_nor2_1
X_5323_ net1744 net393 _0219_ VPWR VGND sg13g2_and2_1
X_7855__157 VPWR VGND net157 sg13g2_tiehi
X_5254_ _1227_ net1455 net700 VPWR VGND sg13g2_nand2_1
X_5185_ net1474 VPWR _1163_ VGND _1102_ _1162_ sg13g2_o21ai_1
X_4205_ net1695 _3568_ _3569_ VPWR VGND sg13g2_nor2_1
X_4136_ VPWR _3512_ net674 VGND sg13g2_inv_1
X_4067_ VPWR _3443_ net534 VGND sg13g2_inv_1
XFILLER_37_794 VPWR VGND sg13g2_fill_2
X_7826_ net188 VGND VPWR _0304_ s0.shift_out\[11\][0] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_948 VPWR VGND sg13g2_decap_8
X_7757_ net263 VGND VPWR _0235_ s0.data_out\[17\]\[2\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_4969_ net1470 net1358 _0967_ VPWR VGND sg13g2_nor2b_1
X_6708_ net1288 VPWR _2533_ VGND net1642 net1277 sg13g2_o21ai_1
X_7688_ net338 VGND VPWR _0166_ s0.data_out\[23\]\[5\] clknet_leaf_41_clk sg13g2_dfrbpq_2
X_6639_ VGND VPWR net1297 _2470_ _2473_ _2472_ sg13g2_a21oi_1
XFILLER_43_720 VPWR VGND sg13g2_fill_1
XFILLER_16_934 VPWR VGND sg13g2_fill_1
XFILLER_28_783 VPWR VGND sg13g2_fill_2
XFILLER_15_433 VPWR VGND sg13g2_fill_1
XFILLER_30_425 VPWR VGND sg13g2_fill_2
XFILLER_7_665 VPWR VGND sg13g2_fill_2
XFILLER_7_698 VPWR VGND sg13g2_fill_2
XFILLER_3_893 VPWR VGND sg13g2_decap_8
Xfanout1650 net1652 net1650 VPWR VGND sg13g2_buf_8
XFILLER_26_4 VPWR VGND sg13g2_fill_2
Xfanout1661 net1662 net1661 VPWR VGND sg13g2_buf_1
X_7642__44 VPWR VGND net44 sg13g2_tiehi
Xfanout1683 net1684 net1683 VPWR VGND sg13g2_buf_8
Xfanout1694 ui_in[3] net1694 VPWR VGND sg13g2_buf_8
Xfanout1672 ui_in[5] net1672 VPWR VGND sg13g2_buf_8
X_6990_ _2788_ net1260 _2787_ VPWR VGND sg13g2_nand2b_1
X_5941_ net1406 VPWR _1846_ VGND _1780_ _1845_ sg13g2_o21ai_1
XFILLER_18_293 VPWR VGND sg13g2_fill_2
X_5872_ _1785_ net1399 net738 VPWR VGND sg13g2_nand2_1
X_7611_ _3323_ VPWR _3349_ VGND _3324_ _3348_ sg13g2_o21ai_1
X_4823_ net1604 _0826_ _0827_ _0170_ VPWR VGND sg13g2_nor3_1
XFILLER_22_937 VPWR VGND sg13g2_fill_1
X_7542_ net1218 VPWR _3290_ VGND _3224_ _3289_ sg13g2_o21ai_1
X_4754_ _0775_ net1512 _0774_ VPWR VGND sg13g2_nand2b_1
X_7473_ s0.data_out\[1\]\[1\] s0.data_out\[0\]\[1\] net1214 _3223_ VPWR VGND sg13g2_mux2_1
X_4685_ _0156_ _0708_ _0709_ _3425_ net1593 VPWR VGND sg13g2_a22oi_1
X_6424_ net1307 s0.data_out\[9\]\[0\] _2281_ VPWR VGND sg13g2_and2_1
X_6355_ net1307 net1355 _2213_ VPWR VGND sg13g2_nor2b_1
X_5306_ net1461 VPWR _1272_ VGND _1211_ _1271_ sg13g2_o21ai_1
X_6286_ net1365 VPWR _2162_ VGND _2103_ _2161_ sg13g2_o21ai_1
X_5237_ s0.data_out\[19\]\[6\] s0.data_out\[18\]\[6\] net1453 _1210_ VPWR VGND sg13g2_mux2_1
X_5168_ net1198 _3455_ _1150_ VPWR VGND sg13g2_nor2_1
X_4119_ VPWR _3495_ net586 VGND sg13g2_inv_1
X_5099_ net1458 net1358 _1084_ VPWR VGND sg13g2_nor2b_1
XFILLER_17_78 VPWR VGND sg13g2_fill_1
X_7809_ net207 VGND VPWR _0287_ s0.data_out\[13\]\[6\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_12_436 VPWR VGND sg13g2_decap_8
XFILLER_13_948 VPWR VGND sg13g2_fill_1
XFILLER_24_285 VPWR VGND sg13g2_decap_8
XFILLER_9_919 VPWR VGND sg13g2_fill_2
XFILLER_32_1003 VPWR VGND sg13g2_decap_8
XFILLER_20_491 VPWR VGND sg13g2_fill_2
XFILLER_0_852 VPWR VGND sg13g2_decap_8
Xhold7 s0.genblk1\[8\].modules.bubble VPWR VGND net376 sg13g2_dlygate4sd3_1
XFILLER_48_823 VPWR VGND sg13g2_decap_8
XFILLER_15_263 VPWR VGND sg13g2_fill_2
XFILLER_31_767 VPWR VGND sg13g2_fill_2
XFILLER_8_996 VPWR VGND sg13g2_decap_8
Xhold407 _0599_ VPWR VGND net776 sg13g2_dlygate4sd3_1
X_4470_ _0514_ VPWR _0515_ VGND net1185 _0512_ sg13g2_o21ai_1
Xhold418 s0.data_out\[11\]\[4\] VPWR VGND net787 sg13g2_dlygate4sd3_1
Xhold429 s0.data_out\[26\]\[0\] VPWR VGND net798 sg13g2_dlygate4sd3_1
X_6140_ VGND VPWR _1900_ _2028_ _2029_ net1379 sg13g2_a21oi_1
X_7676__351 VPWR VGND net351 sg13g2_tiehi
X_6071_ net1379 VPWR _1963_ VGND net1643 net1370 sg13g2_o21ai_1
XFILLER_39_801 VPWR VGND sg13g2_fill_1
XFILLER_38_311 VPWR VGND sg13g2_fill_2
X_5022_ net1690 _0980_ _1020_ VPWR VGND sg13g2_nor2_1
XFILLER_39_878 VPWR VGND sg13g2_fill_2
Xfanout1491 s0.valid_out\[21\][0] net1491 VPWR VGND sg13g2_buf_8
Xfanout1480 net1481 net1480 VPWR VGND sg13g2_buf_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
X_6973_ s0.data_out\[5\]\[2\] s0.data_out\[4\]\[2\] net1255 _2771_ VPWR VGND sg13g2_mux2_1
X_5924_ net1626 _1774_ _1833_ VPWR VGND sg13g2_nor2_1
XFILLER_34_550 VPWR VGND sg13g2_fill_2
X_7918__89 VPWR VGND net89 sg13g2_tiehi
X_5855_ _1753_ VPWR _1768_ VGND net1707 _1760_ sg13g2_o21ai_1
X_4806_ net1593 _0765_ _0820_ VPWR VGND sg13g2_nor2_1
XFILLER_10_907 VPWR VGND sg13g2_fill_1
XFILLER_10_918 VPWR VGND sg13g2_fill_2
XFILLER_16_1009 VPWR VGND sg13g2_decap_8
XFILLER_21_244 VPWR VGND sg13g2_fill_1
X_5786_ _1636_ _1709_ net1747 _1710_ VPWR VGND sg13g2_nand3_1
X_7525_ _3269_ _3273_ net1677 _3275_ VPWR VGND sg13g2_nand3_1
X_4737_ VGND VPWR _0644_ _0757_ _0758_ net1512 sg13g2_a21oi_1
X_7456_ _3208_ VPWR _3209_ VGND net1220 _3097_ sg13g2_o21ai_1
X_4668_ net1592 _0641_ _0697_ VPWR VGND sg13g2_nor2_1
X_6407_ net1312 net1340 _2265_ VPWR VGND sg13g2_nor2b_1
X_4599_ _0631_ _0504_ net1525 _0632_ VPWR VGND sg13g2_a21o_1
X_7387_ VGND VPWR _3032_ _3148_ _3149_ net1230 sg13g2_a21oi_1
X_6338_ _2201_ net1637 net1688 VPWR VGND sg13g2_nand2_1
XFILLER_48_108 VPWR VGND sg13g2_fill_1
X_6269_ s0.data_out\[11\]\[5\] s0.data_out\[10\]\[5\] net1362 _2146_ VPWR VGND sg13g2_mux2_1
XFILLER_28_66 VPWR VGND sg13g2_fill_1
XFILLER_45_837 VPWR VGND sg13g2_decap_8
XFILLER_12_211 VPWR VGND sg13g2_fill_2
XFILLER_13_778 VPWR VGND sg13g2_fill_2
XFILLER_13_789 VPWR VGND sg13g2_fill_1
XFILLER_5_944 VPWR VGND sg13g2_decap_8
XFILLER_4_443 VPWR VGND sg13g2_fill_1
XFILLER_48_620 VPWR VGND sg13g2_decap_4
XFILLER_48_697 VPWR VGND sg13g2_decap_8
X_5640_ net1415 net1340 _1577_ VPWR VGND sg13g2_nor2b_1
X_5571_ _1510_ VPWR _1511_ VGND net1428 _1390_ sg13g2_o21ai_1
X_7310_ net1188 _3540_ _3080_ VPWR VGND sg13g2_nor2_1
X_4522_ VPWR _0567_ _0566_ VGND sg13g2_inv_1
X_7241_ _3015_ net1237 net735 VPWR VGND sg13g2_nand2_1
Xhold226 s0.data_out\[2\]\[5\] VPWR VGND net595 sg13g2_dlygate4sd3_1
X_4453_ _0498_ net481 net1543 VPWR VGND sg13g2_nand2b_1
Xhold204 _0113_ VPWR VGND net573 sg13g2_dlygate4sd3_1
Xhold215 s0.data_out\[5\]\[6\] VPWR VGND net584 sg13g2_dlygate4sd3_1
Xhold259 _0204_ VPWR VGND net628 sg13g2_dlygate4sd3_1
Xhold237 s0.data_out\[15\]\[2\] VPWR VGND net606 sg13g2_dlygate4sd3_1
Xhold248 _0068_ VPWR VGND net617 sg13g2_dlygate4sd3_1
X_4384_ VGND VPWR _3629_ _0440_ _0441_ net1550 sg13g2_a21oi_1
X_7172_ _2956_ VPWR _2957_ VGND net1723 net781 sg13g2_o21ai_1
X_6123_ VGND VPWR net1380 _2009_ _2012_ _2011_ sg13g2_a21oi_1
X_6054_ net1384 net418 _1950_ VPWR VGND sg13g2_and2_1
X_5005_ s0.data_out\[21\]\[5\] s0.data_out\[20\]\[5\] net1478 _1003_ VPWR VGND sg13g2_mux2_1
XFILLER_26_325 VPWR VGND sg13g2_fill_2
X_6956_ net1263 net566 _2758_ VPWR VGND sg13g2_and2_1
X_5907_ VGND VPWR _1820_ net1568 net395 sg13g2_or2_1
X_6887_ s0.data_out\[6\]\[7\] s0.data_out\[5\]\[7\] net1268 _2697_ VPWR VGND sg13g2_mux2_1
XFILLER_10_704 VPWR VGND sg13g2_fill_2
XFILLER_14_68 VPWR VGND sg13g2_fill_1
X_5838_ VGND VPWR _1642_ _1750_ _1751_ net1402 sg13g2_a21oi_1
X_5769_ _1694_ net1417 _1693_ VPWR VGND sg13g2_nand2b_1
X_7508_ VGND VPWR _3258_ _3255_ net1659 sg13g2_or2_1
XFILLER_5_207 VPWR VGND sg13g2_fill_2
X_7439_ VGND VPWR net1222 s0.data_out\[1\]\[5\] _3195_ _3156_ sg13g2_a21oi_1
XFILLER_2_903 VPWR VGND sg13g2_decap_8
XFILLER_7_1018 VPWR VGND sg13g2_decap_8
XFILLER_39_76 VPWR VGND sg13g2_fill_1
XFILLER_29_152 VPWR VGND sg13g2_fill_1
XFILLER_9_568 VPWR VGND sg13g2_fill_1
XFILLER_4_273 VPWR VGND sg13g2_fill_1
X_7673__354 VPWR VGND net354 sg13g2_tiehi
XFILLER_49_962 VPWR VGND sg13g2_decap_8
XFILLER_36_623 VPWR VGND sg13g2_fill_1
X_6810_ net1175 _3521_ _2628_ VPWR VGND sg13g2_nor2_1
X_7790_ net227 VGND VPWR _0268_ s0.shift_out\[14\][0] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_35_177 VPWR VGND sg13g2_fill_1
X_6741_ _2563_ net1177 _2562_ VPWR VGND sg13g2_nand2_1
X_6672_ _2428_ _2504_ _2505_ _2506_ VPWR VGND sg13g2_nor3_1
XFILLER_31_350 VPWR VGND sg13g2_fill_1
XFILLER_32_862 VPWR VGND sg13g2_fill_2
X_5623_ _1558_ net1416 _1559_ _1560_ VPWR VGND sg13g2_a21o_1
X_5554_ VGND VPWR net1426 net457 _1497_ _1455_ sg13g2_a21oi_1
X_4505_ s0.data_out\[25\]\[5\] s0.data_out\[24\]\[5\] net1528 _0550_ VPWR VGND sg13g2_mux2_1
X_5485_ _1434_ net1434 net527 VPWR VGND sg13g2_nand2_1
X_4436_ _0132_ _0483_ _0484_ _3398_ net1579 VPWR VGND sg13g2_a22oi_1
X_7224_ _2997_ VPWR _2998_ VGND net1190 _2995_ sg13g2_o21ai_1
X_4367_ _0424_ net1542 net556 VPWR VGND sg13g2_nand2_1
X_7155_ VGND VPWR _2809_ _2940_ _2941_ net1248 sg13g2_a21oi_1
X_7969__106 VPWR VGND net106 sg13g2_tiehi
X_6106_ _1981_ VPWR _1995_ VGND net1707 _1988_ sg13g2_o21ai_1
X_4298_ _0116_ net453 _0362_ _3410_ net1576 VPWR VGND sg13g2_a22oi_1
X_7086_ net1170 VPWR _2875_ VGND s0.was_valid_out\[3\][0] net1253 sg13g2_o21ai_1
X_6037_ _1936_ VPWR _1937_ VGND net1192 _1935_ sg13g2_o21ai_1
XFILLER_27_623 VPWR VGND sg13g2_fill_2
XFILLER_42_604 VPWR VGND sg13g2_fill_1
XFILLER_26_155 VPWR VGND sg13g2_fill_1
XFILLER_41_114 VPWR VGND sg13g2_fill_1
X_6939_ net1273 VPWR _2745_ VGND _2679_ _2744_ sg13g2_o21ai_1
XFILLER_10_512 VPWR VGND sg13g2_fill_2
XFILLER_41_88 VPWR VGND sg13g2_fill_1
XFILLER_2_777 VPWR VGND sg13g2_decap_8
XFILLER_46_932 VPWR VGND sg13g2_decap_8
XFILLER_17_100 VPWR VGND sg13g2_fill_1
XFILLER_18_645 VPWR VGND sg13g2_decap_8
XFILLER_18_667 VPWR VGND sg13g2_decap_4
XFILLER_33_615 VPWR VGND sg13g2_fill_2
X_5270_ _1243_ _1234_ _1242_ VPWR VGND sg13g2_nand2_1
X_4221_ net1570 VPWR _3585_ VGND _3579_ _3584_ sg13g2_o21ai_1
X_4152_ VPWR _3528_ net693 VGND sg13g2_inv_1
X_4083_ VPWR _3459_ net499 VGND sg13g2_inv_1
XFILLER_37_932 VPWR VGND sg13g2_fill_2
X_7911_ net97 VGND VPWR net667 s0.data_out\[5\]\[5\] clknet_leaf_13_clk sg13g2_dfrbpq_2
XFILLER_36_475 VPWR VGND sg13g2_fill_1
X_7842_ net171 VGND VPWR _0320_ s0.data_new_delayed\[5\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_4985_ _0973_ _0982_ _0983_ VPWR VGND sg13g2_nor2_1
X_7773_ net246 VGND VPWR _0251_ s0.data_out\[16\]\[6\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_23_136 VPWR VGND sg13g2_fill_1
X_6724_ _2544_ net1270 _2545_ _2546_ VPWR VGND sg13g2_a21o_1
X_6655_ VGND VPWR _2379_ _2488_ _2489_ net1296 sg13g2_a21oi_1
X_6586_ net1615 _2356_ _2424_ VPWR VGND sg13g2_nor2_1
X_5606_ s0.data_out\[16\]\[3\] s0.data_out\[15\]\[3\] net1419 _1543_ VPWR VGND sg13g2_mux2_1
X_5537_ net1436 VPWR _1484_ VGND _1401_ _1483_ sg13g2_o21ai_1
X_5468_ _1285_ VPWR _1417_ VGND net1443 _3470_ sg13g2_o21ai_1
X_7207_ net1639 net1235 _2984_ VPWR VGND sg13g2_nor2b_1
Xfanout1309 net1313 net1309 VPWR VGND sg13g2_buf_8
X_5399_ VGND VPWR _1360_ net1568 net392 sg13g2_or2_1
X_4419_ _0128_ _0470_ _0471_ _3409_ net1577 VPWR VGND sg13g2_a22oi_1
X_7138_ s0.data_out\[3\]\[4\] s0.data_out\[4\]\[4\] net1254 _2924_ VPWR VGND sg13g2_mux2_1
X_7069_ net1596 _2831_ _2861_ VPWR VGND sg13g2_nor2_1
XFILLER_28_943 VPWR VGND sg13g2_fill_1
XFILLER_43_902 VPWR VGND sg13g2_fill_1
XFILLER_36_44 VPWR VGND sg13g2_fill_1
XFILLER_43_935 VPWR VGND sg13g2_decap_8
XFILLER_14_136 VPWR VGND sg13g2_fill_2
XFILLER_30_629 VPWR VGND sg13g2_fill_2
XFILLER_23_670 VPWR VGND sg13g2_fill_2
XFILLER_7_858 VPWR VGND sg13g2_fill_1
XFILLER_6_357 VPWR VGND sg13g2_fill_1
X_7654__31 VPWR VGND net31 sg13g2_tiehi
X_7670__357 VPWR VGND net357 sg13g2_tiehi
XFILLER_46_751 VPWR VGND sg13g2_decap_8
X_7848__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_33_412 VPWR VGND sg13g2_fill_1
X_4770_ _0790_ VPWR _0791_ VGND _0750_ _0752_ sg13g2_o21ai_1
XFILLER_20_117 VPWR VGND sg13g2_fill_2
XFILLER_9_151 VPWR VGND sg13g2_decap_4
X_6440_ _0327_ net545 _2293_ _3499_ net1609 VPWR VGND sg13g2_a22oi_1
X_6371_ _2228_ VPWR _2229_ VGND net1315 _3499_ sg13g2_o21ai_1
X_5322_ net1624 _1278_ net476 _0218_ VPWR VGND sg13g2_nor3_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_5253_ _1223_ _1224_ _1226_ VPWR VGND _1225_ sg13g2_nand3b_1
X_4204_ VGND VPWR net1560 _3567_ _3568_ _3563_ sg13g2_a21oi_1
X_5184_ net1198 _3452_ _1162_ VPWR VGND sg13g2_nor2_1
XFILLER_29_718 VPWR VGND sg13g2_decap_8
X_4135_ VPWR _3511_ net547 VGND sg13g2_inv_1
X_4066_ VPWR _3442_ net797 VGND sg13g2_inv_1
XFILLER_25_924 VPWR VGND sg13g2_fill_1
X_7825_ net189 VGND VPWR _0303_ s0.genblk1\[10\].modules.bubble clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
XFILLER_19_1007 VPWR VGND sg13g2_decap_8
XFILLER_24_423 VPWR VGND sg13g2_fill_1
XFILLER_25_946 VPWR VGND sg13g2_fill_1
X_4968_ s0.data_out\[21\]\[0\] s0.data_out\[20\]\[0\] net1478 _0966_ VPWR VGND sg13g2_mux2_1
X_7756_ net264 VGND VPWR _0234_ s0.data_out\[17\]\[1\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_6707_ _0011_ _2531_ _2532_ _3507_ net1600 VPWR VGND sg13g2_a22oi_1
X_4899_ _0893_ VPWR _0908_ VGND _0901_ _0904_ sg13g2_o21ai_1
X_7687_ net339 VGND VPWR _0165_ s0.data_out\[23\]\[4\] clknet_leaf_41_clk sg13g2_dfrbpq_2
XFILLER_22_13 VPWR VGND sg13g2_decap_8
X_6638_ VGND VPWR _2358_ _2471_ _2472_ net1297 sg13g2_a21oi_1
XFILLER_3_305 VPWR VGND sg13g2_fill_2
X_6569_ _3394_ _3510_ _2410_ VPWR VGND sg13g2_nor2_1
X_7651__34 VPWR VGND net34 sg13g2_tiehi
XFILLER_47_559 VPWR VGND sg13g2_fill_1
XFILLER_43_710 VPWR VGND sg13g2_fill_1
XFILLER_27_250 VPWR VGND sg13g2_fill_1
XFILLER_43_754 VPWR VGND sg13g2_fill_2
XFILLER_10_150 VPWR VGND sg13g2_fill_2
XFILLER_3_872 VPWR VGND sg13g2_decap_8
Xfanout1651 net1652 net1651 VPWR VGND sg13g2_buf_1
Xfanout1640 net1642 net1640 VPWR VGND sg13g2_buf_1
Xfanout1662 ui_in[6] net1662 VPWR VGND sg13g2_buf_8
Xfanout1673 net1676 net1673 VPWR VGND sg13g2_buf_8
Xfanout1684 net1685 net1684 VPWR VGND sg13g2_buf_8
Xfanout1695 net1696 net1695 VPWR VGND sg13g2_buf_8
X_5940_ net1194 _3482_ _1845_ VPWR VGND sg13g2_nor2_1
XFILLER_19_762 VPWR VGND sg13g2_fill_1
XFILLER_18_283 VPWR VGND sg13g2_fill_1
X_7610_ VGND VPWR _3346_ _3347_ _3348_ _3327_ sg13g2_a21oi_1
X_5871_ VGND VPWR net1406 _1781_ _1784_ _1783_ sg13g2_a21oi_1
X_4822_ VGND VPWR _3369_ _0828_ _0169_ _0833_ sg13g2_a21oi_1
X_7861__151 VPWR VGND net151 sg13g2_tiehi
X_7541_ net1208 net430 _3289_ VPWR VGND sg13g2_and2_1
X_4753_ VGND VPWR net1494 _0772_ _0774_ _0773_ sg13g2_a21oi_1
X_7472_ VGND VPWR _3112_ _3221_ _3222_ net1218 sg13g2_a21oi_1
XFILLER_30_993 VPWR VGND sg13g2_decap_8
X_6423_ VGND VPWR _2275_ _2279_ _0323_ _2280_ sg13g2_a21oi_1
X_4684_ net1593 _0649_ _0709_ VPWR VGND sg13g2_nor2_1
X_7718__305 VPWR VGND net305 sg13g2_tiehi
X_6354_ VGND VPWR _2212_ _2211_ net1699 sg13g2_or2_1
X_5305_ net1448 s0.data_out\[18\]\[6\] _1271_ VPWR VGND sg13g2_and2_1
X_6285_ net1321 s0.data_out\[10\]\[0\] _2161_ VPWR VGND sg13g2_and2_1
X_5236_ _1209_ net1455 net767 VPWR VGND sg13g2_nand2_1
X_5167_ _0198_ _1148_ _1149_ _3450_ net1607 VPWR VGND sg13g2_a22oi_1
X_5098_ s0.data_out\[20\]\[0\] s0.data_out\[19\]\[0\] net1465 _1083_ VPWR VGND sg13g2_mux2_1
X_4118_ VPWR _3494_ net551 VGND sg13g2_inv_1
XFILLER_44_518 VPWR VGND sg13g2_fill_1
X_4049_ VPWR _3425_ net525 VGND sg13g2_inv_1
X_7808_ net208 VGND VPWR net583 s0.data_out\[13\]\[5\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_33_34 VPWR VGND sg13g2_fill_1
XFILLER_40_757 VPWR VGND sg13g2_fill_2
X_7739_ net283 VGND VPWR _0217_ s0.was_valid_out\[18\][0] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_33_56 VPWR VGND sg13g2_fill_2
X_7838__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_0_831 VPWR VGND sg13g2_decap_8
XFILLER_48_802 VPWR VGND sg13g2_decap_8
Xhold8 s0.genblk1\[12\].modules.bubble VPWR VGND net377 sg13g2_dlygate4sd3_1
XFILLER_48_879 VPWR VGND sg13g2_decap_8
X_7845__168 VPWR VGND net168 sg13g2_tiehi
XFILLER_15_275 VPWR VGND sg13g2_fill_2
X_7927__79 VPWR VGND net79 sg13g2_tiehi
XFILLER_31_746 VPWR VGND sg13g2_fill_2
XFILLER_12_982 VPWR VGND sg13g2_decap_8
XFILLER_8_975 VPWR VGND sg13g2_decap_8
XFILLER_11_470 VPWR VGND sg13g2_fill_1
Xhold408 s0.data_out\[15\]\[4\] VPWR VGND net777 sg13g2_dlygate4sd3_1
Xhold419 _0309_ VPWR VGND net788 sg13g2_dlygate4sd3_1
X_6070_ _0288_ _1961_ _1962_ _3482_ net1629 VPWR VGND sg13g2_a22oi_1
X_5021_ net1673 _1008_ _1019_ VPWR VGND sg13g2_nor2_1
Xfanout1481 s0.valid_out\[20\][0] net1481 VPWR VGND sg13g2_buf_8
Xfanout1492 s0.valid_out\[21\][0] net1492 VPWR VGND sg13g2_buf_1
Xfanout1470 net1471 net1470 VPWR VGND sg13g2_buf_2
XFILLER_0_1013 VPWR VGND sg13g2_decap_8
X_6972_ net1716 net384 _0038_ VPWR VGND sg13g2_and2_1
X_5923_ net1402 VPWR _1832_ VGND _1771_ _1831_ sg13g2_o21ai_1
X_5854_ VPWR VGND _1766_ net1712 _1764_ net1707 _1767_ _1760_ sg13g2_a221oi_1
X_4805_ net1512 VPWR _0819_ VGND _0762_ _0818_ sg13g2_o21ai_1
XFILLER_22_746 VPWR VGND sg13g2_decap_4
X_7524_ VGND VPWR _3269_ _3273_ _3274_ net1677 sg13g2_a21oi_1
X_5785_ net1412 VPWR _1709_ VGND _1637_ _1708_ sg13g2_o21ai_1
X_4736_ _0757_ net558 net1516 VPWR VGND sg13g2_nand2b_1
X_7455_ VPWR _3208_ _3207_ VGND sg13g2_inv_1
X_4667_ net1526 VPWR _0696_ VGND _0638_ _0695_ sg13g2_o21ai_1
X_6406_ s0.data_out\[10\]\[5\] s0.data_out\[9\]\[5\] net1317 _2264_ VPWR VGND sg13g2_mux2_1
X_7386_ _3148_ s0.data_out\[1\]\[7\] net1236 VPWR VGND sg13g2_nand2b_1
X_4598_ _0631_ _3389_ s0.data_out\[23\]\[0\] VPWR VGND sg13g2_nand2_1
X_6337_ VGND VPWR net1637 net1572 _0317_ _2200_ sg13g2_a21oi_1
XFILLER_1_628 VPWR VGND sg13g2_decap_4
X_6268_ _2145_ net1362 net493 VPWR VGND sg13g2_nand2_1
X_6199_ VGND VPWR _2079_ _2078_ _2077_ sg13g2_or2_1
X_5219_ s0.data_out\[19\]\[0\] s0.data_out\[18\]\[0\] net1454 _1192_ VPWR VGND sg13g2_mux2_1
XFILLER_44_33 VPWR VGND sg13g2_fill_1
X_7799__218 VPWR VGND net218 sg13g2_tiehi
XFILLER_40_587 VPWR VGND sg13g2_decap_4
X_7917__90 VPWR VGND net90 sg13g2_tiehi
XFILLER_21_790 VPWR VGND sg13g2_fill_1
XFILLER_5_923 VPWR VGND sg13g2_decap_8
XFILLER_48_676 VPWR VGND sg13g2_decap_8
XFILLER_43_392 VPWR VGND sg13g2_fill_2
XFILLER_15_1010 VPWR VGND sg13g2_decap_8
X_5570_ _1510_ _1509_ _1508_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_772 VPWR VGND sg13g2_fill_1
X_4521_ VGND VPWR _0553_ _0555_ _0566_ net1668 sg13g2_a21oi_1
Xhold205 s0.data_out\[13\]\[4\] VPWR VGND net574 sg13g2_dlygate4sd3_1
Xhold216 s0.data_out\[17\]\[7\] VPWR VGND net585 sg13g2_dlygate4sd3_1
X_4452_ _0495_ net1521 _0496_ _0497_ VPWR VGND sg13g2_a21o_1
X_7240_ _2999_ _3013_ _3014_ VPWR VGND sg13g2_nor2_1
Xhold227 _3198_ VPWR VGND net596 sg13g2_dlygate4sd3_1
Xhold249 s0.data_out\[5\]\[0\] VPWR VGND net618 sg13g2_dlygate4sd3_1
Xhold238 _1718_ VPWR VGND net607 sg13g2_dlygate4sd3_1
X_4383_ _0440_ net431 net1556 VPWR VGND sg13g2_nand2b_1
X_7171_ _2955_ VPWR _2956_ VGND net1170 _2954_ sg13g2_o21ai_1
X_6122_ VGND VPWR _1911_ _2010_ _2011_ net1380 sg13g2_a21oi_1
X_6053_ _0284_ _1948_ _1949_ _3485_ net1628 VPWR VGND sg13g2_a22oi_1
X_5004_ _1002_ net1480 net509 VPWR VGND sg13g2_nand2_1
X_6955_ _0034_ _2756_ _2757_ _3520_ net1597 VPWR VGND sg13g2_a22oi_1
X_5906_ VPWR VGND _1795_ _1740_ _1817_ _1777_ _1819_ _1815_ sg13g2_a221oi_1
XFILLER_22_543 VPWR VGND sg13g2_fill_2
X_6886_ _2696_ net1267 net566 VPWR VGND sg13g2_nand2_1
X_5837_ _1750_ net624 net1408 VPWR VGND sg13g2_nand2b_1
X_5768_ VGND VPWR net1404 _1692_ _1693_ _1690_ sg13g2_a21oi_1
X_7507_ VGND VPWR _3257_ _3249_ net1648 sg13g2_or2_1
X_4719_ _0740_ net1572 _0738_ VPWR VGND sg13g2_xnor2_1
X_7438_ _0080_ _3193_ _3194_ _3539_ net1587 VPWR VGND sg13g2_a22oi_1
X_5699_ net1749 VPWR _1627_ VGND _1624_ _1626_ sg13g2_o21ai_1
X_7369_ _3130_ VPWR _3131_ VGND net1226 _3540_ sg13g2_o21ai_1
X_7952__347 VPWR VGND net347 sg13g2_tiehi
XFILLER_2_959 VPWR VGND sg13g2_decap_8
XFILLER_17_304 VPWR VGND sg13g2_decap_8
XFILLER_45_657 VPWR VGND sg13g2_fill_2
XFILLER_38_1021 VPWR VGND sg13g2_decap_8
X_7666__362 VPWR VGND net362 sg13g2_tiehi
XFILLER_13_565 VPWR VGND sg13g2_decap_8
XFILLER_5_742 VPWR VGND sg13g2_fill_2
XFILLER_49_941 VPWR VGND sg13g2_decap_8
XFILLER_1_992 VPWR VGND sg13g2_decap_8
XFILLER_35_101 VPWR VGND sg13g2_fill_1
XFILLER_24_819 VPWR VGND sg13g2_decap_8
X_6740_ s0.data_out\[6\]\[0\] s0.data_out\[7\]\[0\] net1289 _2562_ VPWR VGND sg13g2_mux2_1
X_6671_ _2481_ _2483_ _2505_ VPWR VGND sg13g2_nor2b_1
X_5622_ net1416 net1335 _1559_ VPWR VGND sg13g2_nor2b_1
X_5553_ VPWR _0237_ net682 VGND sg13g2_inv_1
X_4504_ _0549_ net1530 net407 VPWR VGND sg13g2_nand2_1
X_5484_ _1432_ VPWR _1433_ VGND _1420_ _1430_ sg13g2_o21ai_1
X_4435_ net1579 _0429_ _0484_ VPWR VGND sg13g2_nor2_1
X_7223_ _2997_ net1190 _2996_ VPWR VGND sg13g2_nand2_1
X_4366_ VGND VPWR net1549 _0420_ _0423_ _0422_ sg13g2_a21oi_1
X_7154_ _2940_ s0.data_out\[3\]\[6\] net1253 VPWR VGND sg13g2_nand2b_1
X_6105_ _1994_ _1993_ net1376 VPWR VGND sg13g2_nand2b_1
X_7789__228 VPWR VGND net228 sg13g2_tiehi
X_4297_ net1576 net449 _0362_ VPWR VGND sg13g2_nor2_1
X_7085_ net1241 _2868_ _2874_ VPWR VGND sg13g2_nor2_1
X_6036_ VGND VPWR net1192 _1876_ _1936_ net1627 sg13g2_a21oi_1
X_7906__102 VPWR VGND net102 sg13g2_tiehi
XFILLER_41_148 VPWR VGND sg13g2_fill_1
X_6938_ net1262 net693 _2744_ VPWR VGND sg13g2_and2_1
X_6869_ net1262 net1169 _2679_ VPWR VGND sg13g2_nor2_1
XFILLER_41_67 VPWR VGND sg13g2_fill_2
XFILLER_2_756 VPWR VGND sg13g2_decap_8
XFILLER_46_911 VPWR VGND sg13g2_decap_8
XFILLER_18_613 VPWR VGND sg13g2_fill_2
XFILLER_46_988 VPWR VGND sg13g2_decap_8
XFILLER_33_627 VPWR VGND sg13g2_fill_1
XFILLER_14_830 VPWR VGND sg13g2_fill_2
XFILLER_12_1024 VPWR VGND sg13g2_decap_4
X_4220_ _3583_ net1560 _3584_ VPWR VGND sg13g2_nor2b_1
X_4151_ VPWR _3527_ net668 VGND sg13g2_inv_1
X_4082_ VPWR _3458_ net700 VGND sg13g2_inv_1
X_7910_ net98 VGND VPWR net669 s0.data_out\[5\]\[4\] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_7841_ net172 VGND VPWR _0319_ s0.data_new_delayed\[4\] clknet_leaf_13_clk sg13g2_dfrbpq_2
XFILLER_36_432 VPWR VGND sg13g2_fill_1
X_4984_ _0981_ VPWR _0982_ VGND net1573 _0956_ sg13g2_o21ai_1
X_7772_ net247 VGND VPWR _0250_ s0.data_out\[16\]\[5\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_6723_ net1270 net1349 _2545_ VPWR VGND sg13g2_nor2b_1
X_6654_ _2488_ net653 net1303 VPWR VGND sg13g2_nand2b_1
XFILLER_31_170 VPWR VGND sg13g2_fill_1
X_5605_ _1542_ net1422 net765 VPWR VGND sg13g2_nand2_1
X_6585_ net1309 VPWR _2423_ VGND _2353_ _2422_ sg13g2_o21ai_1
X_5536_ net1423 net495 _1483_ VPWR VGND sg13g2_and2_1
X_5467_ VGND VPWR net1423 _1414_ _1416_ _1415_ sg13g2_a21oi_1
X_4418_ net1577 _0413_ _0471_ VPWR VGND sg13g2_nor2_1
X_7206_ net1239 VPWR _2983_ VGND net1639 net1229 sg13g2_o21ai_1
X_5398_ _1278_ _1279_ _1357_ _1358_ _1359_ VPWR VGND sg13g2_nor4_1
XFILLER_28_1020 VPWR VGND sg13g2_decap_8
X_4349_ VPWR VGND _0405_ net1710 _0403_ net1701 _0406_ _0399_ sg13g2_a221oi_1
X_7137_ VGND VPWR net1242 _2922_ _2923_ _2920_ sg13g2_a21oi_1
X_7068_ net1263 VPWR _2860_ VGND _2828_ _2859_ sg13g2_o21ai_1
X_6019_ net1382 net1331 _1920_ VPWR VGND sg13g2_nor2b_1
XFILLER_43_914 VPWR VGND sg13g2_decap_8
XFILLER_36_67 VPWR VGND sg13g2_fill_2
XFILLER_28_999 VPWR VGND sg13g2_decap_8
XFILLER_42_468 VPWR VGND sg13g2_fill_1
X_7663__365 VPWR VGND net365 sg13g2_tiehi
XFILLER_7_826 VPWR VGND sg13g2_fill_2
XFILLER_42_1017 VPWR VGND sg13g2_decap_8
XFILLER_2_597 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_730 VPWR VGND sg13g2_decap_8
XFILLER_33_468 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_40_clk clknet_3_1__leaf_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_6370_ _2228_ net1315 net544 VPWR VGND sg13g2_nand2_1
X_5321_ net1624 _1280_ _1284_ _0217_ VPWR VGND sg13g2_nor3_1
X_5252_ net1654 _1222_ _1225_ VPWR VGND sg13g2_nor2_1
X_5183_ _0202_ _1160_ _1161_ _3446_ net1607 VPWR VGND sg13g2_a22oi_1
X_4203_ _3565_ net1547 _3566_ _3567_ VPWR VGND sg13g2_a21o_1
X_4134_ VPWR _3510_ net818 VGND sg13g2_inv_1
X_7660__24 VPWR VGND net24 sg13g2_tiehi
X_4065_ VPWR _3441_ net538 VGND sg13g2_inv_1
XFILLER_37_785 VPWR VGND sg13g2_fill_1
X_7824_ net190 VGND VPWR _0302_ s0.valid_out\[11\][0] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_7903__105 VPWR VGND net105 sg13g2_tiehi
X_4967_ VGND VPWR _0961_ _0963_ _0965_ net1705 sg13g2_a21oi_1
X_7755_ net265 VGND VPWR _0233_ s0.data_out\[17\]\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_7971__80 VPWR VGND net80 sg13g2_tiehi
X_6706_ net1600 _2479_ _2532_ VPWR VGND sg13g2_nor2_1
X_4898_ _0885_ _0906_ _0866_ _0907_ VPWR VGND sg13g2_nand3_1
X_7686_ net340 VGND VPWR net811 s0.data_out\[23\]\[3\] clknet_leaf_40_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_31_clk clknet_3_5__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
X_6637_ _2471_ s0.data_out\[7\]\[6\] net1304 VPWR VGND sg13g2_nand2b_1
XFILLER_4_807 VPWR VGND sg13g2_decap_8
X_6568_ _0339_ _2408_ _2409_ _3504_ net1608 VPWR VGND sg13g2_a22oi_1
X_5519_ _1465_ _1467_ net1683 _1468_ VPWR VGND sg13g2_nand3_1
X_6499_ net1295 net1168 _2345_ VPWR VGND sg13g2_nor2_1
XFILLER_15_402 VPWR VGND sg13g2_fill_1
XFILLER_27_273 VPWR VGND sg13g2_decap_4
X_7939__66 VPWR VGND net66 sg13g2_tiehi
X_7960__243 VPWR VGND net243 sg13g2_tiehi
XFILLER_30_427 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_22_clk clknet_3_7__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_8_49 VPWR VGND sg13g2_fill_1
XFILLER_7_667 VPWR VGND sg13g2_fill_1
XFILLER_3_851 VPWR VGND sg13g2_decap_8
Xfanout1641 net1642 net1641 VPWR VGND sg13g2_buf_8
XFILLER_26_6 VPWR VGND sg13g2_fill_1
Xfanout1630 net1631 net1630 VPWR VGND sg13g2_buf_8
Xfanout1663 net1667 net1663 VPWR VGND sg13g2_buf_8
Xfanout1652 ui_in[7] net1652 VPWR VGND sg13g2_buf_8
Xfanout1674 net1676 net1674 VPWR VGND sg13g2_buf_8
Xfanout1685 ui_in[4] net1685 VPWR VGND sg13g2_buf_8
Xfanout1696 net1700 net1696 VPWR VGND sg13g2_buf_8
XFILLER_18_251 VPWR VGND sg13g2_decap_8
X_5870_ VGND VPWR _1663_ _1782_ _1783_ net1406 sg13g2_a21oi_1
X_4821_ net1734 VPWR _0833_ VGND _0830_ _0832_ sg13g2_o21ai_1
Xclkbuf_leaf_13_clk clknet_3_3__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_7540_ VPWR _0088_ net800 VGND sg13g2_inv_1
X_4752_ net1494 net1339 _0773_ VPWR VGND sg13g2_nor2b_1
X_7471_ _3221_ net430 net1224 VPWR VGND sg13g2_nand2b_1
X_4683_ net1523 VPWR _0708_ VGND _0646_ _0707_ sg13g2_o21ai_1
XFILLER_30_972 VPWR VGND sg13g2_decap_8
X_6422_ VGND VPWR _2280_ net1567 net388 sg13g2_or2_1
X_6353_ VGND VPWR net1319 _2208_ _2211_ _2210_ sg13g2_a21oi_1
X_6284_ VGND VPWR _2157_ _2159_ _0304_ _2160_ sg13g2_a21oi_1
X_5304_ VPWR _0214_ _1270_ VGND sg13g2_inv_1
X_5235_ _1207_ VPWR _1208_ VGND _1198_ _1199_ sg13g2_o21ai_1
XFILLER_25_1023 VPWR VGND sg13g2_decap_4
X_5166_ net1607 _1081_ _1149_ VPWR VGND sg13g2_nor2_1
X_5097_ VGND VPWR net1475 _1079_ _1082_ _1081_ sg13g2_a21oi_1
XFILLER_17_14 VPWR VGND sg13g2_decap_4
X_4117_ VPWR _3493_ net760 VGND sg13g2_inv_1
X_4048_ VPWR _3424_ net556 VGND sg13g2_inv_1
X_5999_ _1900_ net1387 net746 VPWR VGND sg13g2_nand2_1
X_7807_ net209 VGND VPWR _0285_ s0.data_out\[13\]\[4\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_7738_ net284 VGND VPWR net673 s0.data_out\[19\]\[7\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_7669_ net358 VGND VPWR _0147_ s0.genblk1\[23\].modules.bubble clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_20_493 VPWR VGND sg13g2_fill_1
XFILLER_4_604 VPWR VGND sg13g2_fill_1
XFILLER_0_810 VPWR VGND sg13g2_decap_8
XFILLER_0_887 VPWR VGND sg13g2_decap_8
Xhold9 s0.genblk1\[5\].modules.bubble VPWR VGND net378 sg13g2_dlygate4sd3_1
XFILLER_48_858 VPWR VGND sg13g2_decap_8
XFILLER_16_711 VPWR VGND sg13g2_fill_1
XFILLER_16_722 VPWR VGND sg13g2_fill_2
XFILLER_16_744 VPWR VGND sg13g2_fill_2
XFILLER_31_769 VPWR VGND sg13g2_fill_1
XFILLER_12_972 VPWR VGND sg13g2_fill_1
XFILLER_8_954 VPWR VGND sg13g2_decap_8
Xhold409 s0.data_out\[19\]\[5\] VPWR VGND net778 sg13g2_dlygate4sd3_1
XFILLER_48_1012 VPWR VGND sg13g2_decap_8
X_5020_ VGND VPWR _1014_ _1016_ _1018_ net1682 sg13g2_a21oi_1
Xclkbuf_leaf_2_clk clknet_3_0__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
Xfanout1493 net1497 net1493 VPWR VGND sg13g2_buf_8
Xfanout1482 net1485 net1482 VPWR VGND sg13g2_buf_8
Xfanout1460 s0.shift_out\[19\][0] net1460 VPWR VGND sg13g2_buf_8
Xfanout1471 net1472 net1471 VPWR VGND sg13g2_buf_1
X_6971_ net1591 _2763_ _2764_ _0037_ VPWR VGND sg13g2_nor3_1
X_5922_ net1194 _3485_ _1831_ VPWR VGND sg13g2_nor2_1
XFILLER_34_552 VPWR VGND sg13g2_fill_1
X_5853_ _1766_ net1195 _1765_ VPWR VGND sg13g2_nand2_1
X_4804_ net1493 net552 _0818_ VPWR VGND sg13g2_and2_1
X_5784_ net1401 s0.data_out\[14\]\[0\] _1708_ VPWR VGND sg13g2_and2_1
XFILLER_34_596 VPWR VGND sg13g2_fill_1
X_7523_ _3273_ net1223 _3272_ VPWR VGND sg13g2_nand2b_1
X_4735_ _0754_ net1493 _0755_ _0756_ VPWR VGND sg13g2_a21o_1
XFILLER_21_257 VPWR VGND sg13g2_decap_4
X_7454_ VGND VPWR net1633 net1216 _3207_ _3206_ sg13g2_a21oi_1
X_4666_ net1182 _3434_ _0695_ VPWR VGND sg13g2_nor2_1
X_6405_ _2263_ net1316 s0.data_out\[9\]\[5\] VPWR VGND sg13g2_nand2_1
X_4597_ _0630_ net1525 _0629_ VPWR VGND sg13g2_nand2b_1
X_7385_ _3145_ net1219 _3146_ _3147_ VPWR VGND sg13g2_a21o_1
XFILLER_1_607 VPWR VGND sg13g2_decap_8
X_6336_ net1637 net1349 _2200_ VPWR VGND sg13g2_nor2_1
X_6267_ net1682 _2143_ _2144_ VPWR VGND sg13g2_and2_1
XFILLER_0_139 VPWR VGND sg13g2_decap_4
X_6198_ net1643 net1363 _2078_ VPWR VGND sg13g2_nor2b_1
X_5218_ VGND VPWR net1459 _1188_ _1191_ _1190_ sg13g2_a21oi_1
X_5149_ _1133_ VPWR _1134_ VGND net1692 _1097_ sg13g2_o21ai_1
XFILLER_29_379 VPWR VGND sg13g2_fill_1
XFILLER_40_577 VPWR VGND sg13g2_fill_1
XFILLER_8_217 VPWR VGND sg13g2_fill_2
XFILLER_5_902 VPWR VGND sg13g2_decap_8
XFILLER_5_979 VPWR VGND sg13g2_decap_8
X_7851__162 VPWR VGND net162 sg13g2_tiehi
XFILLER_0_684 VPWR VGND sg13g2_decap_8
XFILLER_48_655 VPWR VGND sg13g2_decap_8
XFILLER_29_891 VPWR VGND sg13g2_fill_1
XFILLER_35_316 VPWR VGND sg13g2_fill_1
XFILLER_16_541 VPWR VGND sg13g2_fill_1
XFILLER_44_883 VPWR VGND sg13g2_decap_8
XFILLER_16_585 VPWR VGND sg13g2_fill_1
X_7708__316 VPWR VGND net316 sg13g2_tiehi
XFILLER_16_596 VPWR VGND sg13g2_fill_2
X_4520_ _0565_ _0556_ _0564_ VPWR VGND sg13g2_nand2_1
Xhold217 s0.data_out\[11\]\[7\] VPWR VGND net586 sg13g2_dlygate4sd3_1
Xhold206 s0.data_out\[13\]\[7\] VPWR VGND net575 sg13g2_dlygate4sd3_1
XFILLER_7_261 VPWR VGND sg13g2_decap_4
X_4451_ net1521 net1352 _0496_ VPWR VGND sg13g2_nor2b_1
Xhold239 s0.data_out\[8\]\[6\] VPWR VGND net608 sg13g2_dlygate4sd3_1
Xhold228 s0.data_out\[12\]\[3\] VPWR VGND net597 sg13g2_dlygate4sd3_1
X_7170_ VGND VPWR net1170 _2894_ _2955_ net1585 sg13g2_a21oi_1
X_6121_ _2010_ s0.data_out\[11\]\[6\] net1387 VPWR VGND sg13g2_nand2b_1
XFILLER_4_990 VPWR VGND sg13g2_decap_8
X_4382_ _0437_ net1534 _0438_ _0439_ VPWR VGND sg13g2_a21o_1
X_7715__309 VPWR VGND net309 sg13g2_tiehi
XFILLER_39_611 VPWR VGND sg13g2_fill_2
X_6052_ net1628 _1887_ _1949_ VPWR VGND sg13g2_nor2_1
X_5003_ _1000_ _0998_ _1001_ VPWR VGND _0999_ sg13g2_nand3b_1
XFILLER_22_1015 VPWR VGND sg13g2_decap_8
Xfanout1290 s0.valid_out\[7\][0] net1290 VPWR VGND sg13g2_buf_1
XFILLER_26_327 VPWR VGND sg13g2_fill_1
X_6954_ net1597 _2694_ _2757_ VPWR VGND sg13g2_nor2_1
XFILLER_26_349 VPWR VGND sg13g2_fill_2
X_5905_ _1818_ _1793_ _1792_ VPWR VGND sg13g2_nand2b_1
X_6885_ VGND VPWR net1274 _2692_ _2695_ _2694_ sg13g2_a21oi_1
XFILLER_14_15 VPWR VGND sg13g2_decap_4
XFILLER_22_533 VPWR VGND sg13g2_fill_2
X_7828__186 VPWR VGND net186 sg13g2_tiehi
XFILLER_10_706 VPWR VGND sg13g2_fill_1
X_5836_ _1747_ net1391 _1748_ _1749_ VPWR VGND sg13g2_a21o_1
X_5767_ s0.data_out\[15\]\[4\] s0.data_out\[14\]\[4\] net1410 _1692_ VPWR VGND sg13g2_mux2_1
X_7506_ _3256_ _3255_ net1659 _3249_ net1648 VPWR VGND sg13g2_a22oi_1
X_4718_ VGND VPWR _0739_ _0738_ net1572 sg13g2_or2_1
X_7914__94 VPWR VGND net94 sg13g2_tiehi
X_5698_ _1626_ _1623_ _1625_ VPWR VGND sg13g2_nand2_1
X_7437_ net1587 _3168_ _3194_ VPWR VGND sg13g2_nor2_1
X_4649_ _0658_ _0660_ _0682_ VPWR VGND sg13g2_nor2b_1
X_7368_ _3130_ net1226 s0.data_out\[1\]\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_2_938 VPWR VGND sg13g2_decap_8
XFILLER_1_426 VPWR VGND sg13g2_decap_8
X_7835__179 VPWR VGND net179 sg13g2_tiehi
X_6319_ net1323 VPWR _2187_ VGND net1646 net1311 sg13g2_o21ai_1
X_7299_ VPWR _0064_ _3071_ VGND sg13g2_inv_1
XFILLER_38_1000 VPWR VGND sg13g2_decap_8
XFILLER_41_897 VPWR VGND sg13g2_fill_1
XFILLER_5_710 VPWR VGND sg13g2_fill_2
XFILLER_4_253 VPWR VGND sg13g2_fill_1
XFILLER_45_1026 VPWR VGND sg13g2_fill_2
XFILLER_1_971 VPWR VGND sg13g2_decap_8
XFILLER_49_920 VPWR VGND sg13g2_decap_8
XFILLER_49_997 VPWR VGND sg13g2_decap_8
X_6670_ _2484_ _2497_ _2499_ _2504_ VPWR VGND sg13g2_nor3_1
X_7721__302 VPWR VGND net302 sg13g2_tiehi
X_5621_ s0.data_out\[16\]\[6\] s0.data_out\[15\]\[6\] net1421 _1558_ VPWR VGND sg13g2_mux2_1
X_5552_ _1495_ VPWR _1496_ VGND net1745 net681 sg13g2_o21ai_1
X_4503_ _0546_ _0544_ _0548_ VPWR VGND _0545_ sg13g2_nand3b_1
X_5483_ _1432_ net1692 _1429_ VPWR VGND sg13g2_nand2_1
X_7911__97 VPWR VGND net97 sg13g2_tiehi
X_4434_ net1550 VPWR _0483_ VGND _0426_ _0482_ sg13g2_o21ai_1
X_7222_ s0.data_out\[2\]\[1\] s0.data_out\[3\]\[1\] net1247 _2996_ VPWR VGND sg13g2_mux2_1
X_4365_ VGND VPWR _3608_ _0421_ _0422_ net1549 sg13g2_a21oi_1
X_7153_ _2937_ net1241 _2938_ _2939_ VPWR VGND sg13g2_a21o_1
X_7084_ _2870_ VPWR _2873_ VGND s0.was_valid_out\[3\][0] net1246 sg13g2_o21ai_1
X_6104_ s0.data_out\[11\]\[0\] s0.data_out\[12\]\[0\] net1386 _1993_ VPWR VGND sg13g2_mux2_1
X_4296_ net1561 VPWR _0361_ VGND _3592_ _0360_ sg13g2_o21ai_1
X_6035_ VGND VPWR net1378 net692 _1935_ _1874_ sg13g2_a21oi_1
XFILLER_27_625 VPWR VGND sg13g2_fill_1
X_6937_ VPWR _0030_ net533 VGND sg13g2_inv_1
X_6868_ _2677_ VPWR _2678_ VGND net1266 _3521_ sg13g2_o21ai_1
XFILLER_10_514 VPWR VGND sg13g2_fill_1
X_5819_ net1630 _1668_ _1736_ VPWR VGND sg13g2_nor2_1
X_7841__172 VPWR VGND net172 sg13g2_tiehi
X_6799_ _2619_ VPWR _2620_ VGND net1177 _2618_ sg13g2_o21ai_1
XFILLER_2_735 VPWR VGND sg13g2_decap_8
XFILLER_46_967 VPWR VGND sg13g2_decap_8
XFILLER_33_617 VPWR VGND sg13g2_fill_1
XFILLER_9_334 VPWR VGND sg13g2_fill_1
X_7705__319 VPWR VGND net319 sg13g2_tiehi
XFILLER_12_1003 VPWR VGND sg13g2_decap_8
XFILLER_13_396 VPWR VGND sg13g2_fill_1
X_4150_ VPWR _3526_ net666 VGND sg13g2_inv_1
X_4081_ VPWR _3457_ net805 VGND sg13g2_inv_1
XFILLER_49_794 VPWR VGND sg13g2_decap_8
X_7840_ net173 VGND VPWR _0318_ s0.data_new_delayed\[3\] clknet_leaf_38_clk sg13g2_dfrbpq_2
XFILLER_37_989 VPWR VGND sg13g2_decap_8
X_4983_ _0981_ net1690 _0980_ VPWR VGND sg13g2_nand2_1
X_7771_ net248 VGND VPWR _0249_ s0.data_out\[16\]\[4\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_6722_ s0.data_out\[7\]\[2\] s0.data_out\[6\]\[2\] net1278 _2544_ VPWR VGND sg13g2_mux2_1
X_7825__189 VPWR VGND net189 sg13g2_tiehi
X_6653_ _2485_ net1286 _2486_ _2487_ VPWR VGND sg13g2_a21o_1
X_5604_ _1525_ _1533_ _1540_ _1541_ VPWR VGND sg13g2_nor3_1
XFILLER_31_193 VPWR VGND sg13g2_fill_2
X_6584_ _3394_ _3507_ _2422_ VPWR VGND sg13g2_nor2_1
X_5535_ VPWR _0233_ net690 VGND sg13g2_inv_1
X_7795__222 VPWR VGND net222 sg13g2_tiehi
X_5466_ net1424 net1350 _1415_ VPWR VGND sg13g2_nor2b_1
X_4417_ net1551 VPWR _0470_ VGND _0410_ _0469_ sg13g2_o21ai_1
X_7205_ _0059_ _2981_ _2982_ _3531_ net1586 VPWR VGND sg13g2_a22oi_1
X_5397_ _1332_ _1334_ _1358_ VPWR VGND sg13g2_nor2b_1
X_4348_ _0405_ _0404_ net1552 VPWR VGND sg13g2_nand2b_1
X_7136_ s0.data_out\[4\]\[4\] s0.data_out\[3\]\[4\] net1245 _2922_ VPWR VGND sg13g2_mux2_1
X_4279_ _3556_ _0346_ _0347_ _0348_ VPWR VGND sg13g2_nor3_1
X_7067_ net1252 s0.data_out\[4\]\[5\] _2859_ VPWR VGND sg13g2_and2_1
X_6018_ s0.data_out\[13\]\[7\] s0.data_out\[12\]\[7\] net1389 _1919_ VPWR VGND sg13g2_mux2_1
XFILLER_27_400 VPWR VGND sg13g2_fill_2
XFILLER_28_912 VPWR VGND sg13g2_fill_1
XFILLER_27_444 VPWR VGND sg13g2_decap_8
XFILLER_28_978 VPWR VGND sg13g2_decap_8
X_7969_ net106 VGND VPWR _0103_ s0.data_out\[0\]\[3\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_27_499 VPWR VGND sg13g2_decap_8
XFILLER_35_1025 VPWR VGND sg13g2_decap_4
XFILLER_38_709 VPWR VGND sg13g2_fill_1
XFILLER_46_786 VPWR VGND sg13g2_decap_8
XFILLER_33_458 VPWR VGND sg13g2_fill_1
X_7779__239 VPWR VGND net239 sg13g2_tiehi
X_5320_ VPWR VGND net1205 _1282_ _1283_ _1278_ _1284_ _1281_ sg13g2_a221oi_1
X_5251_ VGND VPWR _1224_ _1215_ net1664 sg13g2_or2_1
X_4202_ net1547 net1348 _3566_ VPWR VGND sg13g2_nor2b_1
X_5182_ net1606 _1130_ _1161_ VPWR VGND sg13g2_nor2_1
X_4133_ VPWR _3509_ net426 VGND sg13g2_inv_1
XFILLER_3_1012 VPWR VGND sg13g2_decap_8
X_4064_ VPWR _3440_ net599 VGND sg13g2_inv_1
XFILLER_49_591 VPWR VGND sg13g2_decap_8
X_7823_ net192 VGND VPWR _0301_ s0.was_valid_out\[11\][0] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_7754_ net266 VGND VPWR _0232_ s0.shift_out\[17\][0] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_6705_ net1297 VPWR _2531_ VGND _2476_ _2530_ sg13g2_o21ai_1
X_4966_ _0961_ _0963_ net1706 _0964_ VPWR VGND sg13g2_nand3_1
XFILLER_33_981 VPWR VGND sg13g2_decap_8
X_4897_ _0902_ _0903_ _0904_ _0905_ _0906_ VPWR VGND sg13g2_nor4_1
X_7685_ net341 VGND VPWR _0163_ s0.data_out\[23\]\[2\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_6636_ _2468_ net1286 _2469_ _2470_ VPWR VGND sg13g2_a21o_1
X_6567_ net1608 _2348_ _2409_ VPWR VGND sg13g2_nor2_1
XFILLER_3_307 VPWR VGND sg13g2_fill_1
X_5518_ _1467_ _3375_ _1466_ VPWR VGND sg13g2_nand2_1
X_6498_ _2343_ VPWR _2344_ VGND net1302 _3504_ sg13g2_o21ai_1
X_5449_ net1748 net391 _0231_ VPWR VGND sg13g2_and2_1
X_7119_ VGND VPWR _2793_ _2904_ _2905_ net1249 sg13g2_a21oi_1
XFILLER_47_56 VPWR VGND sg13g2_fill_2
XFILLER_43_756 VPWR VGND sg13g2_fill_1
XFILLER_31_929 VPWR VGND sg13g2_fill_1
XFILLER_6_156 VPWR VGND sg13g2_fill_1
Xfanout1642 uio_in[0] net1642 VPWR VGND sg13g2_buf_8
Xfanout1620 net1621 net1620 VPWR VGND sg13g2_buf_8
Xfanout1631 net1632 net1631 VPWR VGND sg13g2_buf_8
Xfanout1653 net1657 net1653 VPWR VGND sg13g2_buf_8
Xfanout1664 net1666 net1664 VPWR VGND sg13g2_buf_8
Xfanout1675 net1676 net1675 VPWR VGND sg13g2_buf_8
Xfanout1697 net1700 net1697 VPWR VGND sg13g2_buf_8
Xfanout1686 net1687 net1686 VPWR VGND sg13g2_buf_8
XFILLER_18_274 VPWR VGND sg13g2_fill_1
X_4820_ _0829_ VPWR _0832_ VGND net1498 _0831_ sg13g2_o21ai_1
X_4751_ s0.data_out\[23\]\[5\] s0.data_out\[22\]\[5\] net1503 _0772_ VPWR VGND sg13g2_mux2_1
X_7470_ VGND VPWR net1201 _3215_ _3220_ _3219_ sg13g2_a21oi_1
X_4682_ net1181 _3432_ _0707_ VPWR VGND sg13g2_nor2_1
X_6421_ _2195_ _2277_ _2278_ _2279_ VPWR VGND sg13g2_nor3_1
X_7792__225 VPWR VGND net225 sg13g2_tiehi
X_6352_ VGND VPWR _2087_ _2209_ _2210_ net1319 sg13g2_a21oi_1
X_6283_ VGND VPWR _2160_ net1567 net390 sg13g2_or2_1
X_5303_ _1269_ VPWR _1270_ VGND net1742 net778 sg13g2_o21ai_1
X_5234_ _1207_ _1206_ net1692 _1183_ net1697 VPWR VGND sg13g2_a22oi_1
X_5165_ net1475 VPWR _1148_ VGND _1078_ _1147_ sg13g2_o21ai_1
XFILLER_25_1002 VPWR VGND sg13g2_decap_8
X_4116_ VPWR _3492_ net675 VGND sg13g2_inv_1
X_5096_ VGND VPWR _0958_ _1080_ _1081_ net1475 sg13g2_a21oi_1
X_4047_ VPWR _3423_ s0.data_out\[25\]\[2\] VGND sg13g2_inv_1
XFILLER_25_723 VPWR VGND sg13g2_fill_1
XFILLER_13_907 VPWR VGND sg13g2_fill_2
X_7806_ net210 VGND VPWR net758 s0.data_out\[13\]\[3\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_5998_ _1899_ net1684 _1898_ VPWR VGND sg13g2_nand2_1
X_4949_ net1736 VPWR _0949_ VGND _0946_ _0948_ sg13g2_o21ai_1
X_7737_ net285 VGND VPWR net646 s0.data_out\[19\]\[6\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_24_299 VPWR VGND sg13g2_decap_8
XFILLER_33_58 VPWR VGND sg13g2_fill_1
X_7668_ net359 VGND VPWR _0146_ s0.valid_out\[24\][0] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_21_984 VPWR VGND sg13g2_decap_8
XFILLER_32_1017 VPWR VGND sg13g2_decap_8
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
X_6619_ _2453_ net1293 _2452_ VPWR VGND sg13g2_nand2b_1
X_7599_ _3332_ _3333_ _3336_ _3337_ VPWR VGND sg13g2_or3_1
XFILLER_0_866 VPWR VGND sg13g2_decap_8
XFILLER_48_837 VPWR VGND sg13g2_decap_8
XFILLER_31_748 VPWR VGND sg13g2_fill_1
XFILLER_7_432 VPWR VGND sg13g2_fill_2
Xfanout1450 net1451 net1450 VPWR VGND sg13g2_buf_8
Xfanout1483 net1485 net1483 VPWR VGND sg13g2_buf_8
Xfanout1472 net1477 net1472 VPWR VGND sg13g2_buf_1
Xfanout1461 net1463 net1461 VPWR VGND sg13g2_buf_8
XFILLER_38_358 VPWR VGND sg13g2_fill_1
Xfanout1494 net1497 net1494 VPWR VGND sg13g2_buf_1
X_6970_ VGND VPWR _3362_ _2765_ _0036_ _2770_ sg13g2_a21oi_1
XFILLER_47_892 VPWR VGND sg13g2_decap_8
X_5921_ _0271_ _1829_ _1830_ _3480_ net1626 VPWR VGND sg13g2_a22oi_1
X_5852_ s0.data_out\[13\]\[0\] s0.data_out\[14\]\[0\] net1408 _1765_ VPWR VGND sg13g2_mux2_1
X_4803_ VPWR _0166_ _0817_ VGND sg13g2_inv_1
X_5783_ VGND VPWR _1703_ _1706_ _0256_ _1707_ sg13g2_a21oi_1
X_7900__109 VPWR VGND net109 sg13g2_tiehi
X_7522_ VGND VPWR net1211 _3270_ _3272_ _3271_ sg13g2_a21oi_1
XFILLER_9_60 VPWR VGND sg13g2_fill_1
X_4734_ net1493 net1329 _0755_ VPWR VGND sg13g2_nor2b_1
X_7926__81 VPWR VGND net81 sg13g2_tiehi
X_7453_ net1220 VPWR _3206_ VGND net1640 net1209 sg13g2_o21ai_1
X_4665_ _0151_ _0693_ _0694_ _3430_ net1589 VPWR VGND sg13g2_a22oi_1
X_6404_ _2259_ _2261_ net1682 _2262_ VPWR VGND sg13g2_nand3_1
X_4596_ VGND VPWR net1510 _0627_ _0629_ _0628_ sg13g2_a21oi_1
X_7384_ net1219 net1328 _3146_ VPWR VGND sg13g2_nor2b_1
X_6335_ VGND VPWR net1638 _3415_ _0316_ _2199_ sg13g2_a21oi_1
X_6266_ VGND VPWR net1368 _2140_ _2143_ _2142_ sg13g2_a21oi_1
X_6197_ net1369 VPWR _2077_ VGND net1326 net1643 sg13g2_o21ai_1
X_5217_ VGND VPWR _1076_ _1189_ _1190_ net1458 sg13g2_a21oi_1
X_5148_ _1133_ net1673 _1131_ VPWR VGND sg13g2_nand2_1
X_5079_ net1736 VPWR _1067_ VGND net651 _1061_ sg13g2_o21ai_1
XFILLER_37_380 VPWR VGND sg13g2_fill_1
XFILLER_25_575 VPWR VGND sg13g2_fill_1
XFILLER_25_586 VPWR VGND sg13g2_fill_2
XFILLER_13_748 VPWR VGND sg13g2_fill_1
XFILLER_21_781 VPWR VGND sg13g2_fill_2
XFILLER_5_958 VPWR VGND sg13g2_decap_8
XFILLER_0_652 VPWR VGND sg13g2_decap_8
XFILLER_0_663 VPWR VGND sg13g2_decap_8
XFILLER_48_634 VPWR VGND sg13g2_decap_8
XFILLER_18_80 VPWR VGND sg13g2_decap_8
XFILLER_47_199 VPWR VGND sg13g2_fill_2
XFILLER_44_840 VPWR VGND sg13g2_decap_4
XFILLER_16_520 VPWR VGND sg13g2_fill_2
XFILLER_44_862 VPWR VGND sg13g2_decap_8
XFILLER_43_394 VPWR VGND sg13g2_fill_1
X_7923__84 VPWR VGND net84 sg13g2_tiehi
Xhold207 _0288_ VPWR VGND net576 sg13g2_dlygate4sd3_1
X_4450_ _0494_ VPWR _0495_ VGND net1529 _3421_ sg13g2_o21ai_1
Xhold218 _0312_ VPWR VGND net587 sg13g2_dlygate4sd3_1
X_4381_ net1534 net1343 _0438_ VPWR VGND sg13g2_nor2b_1
Xhold229 _0296_ VPWR VGND net598 sg13g2_dlygate4sd3_1
X_6120_ _2007_ net1370 _2008_ _2009_ VPWR VGND sg13g2_a21o_1
X_6051_ net1390 VPWR _1948_ VGND _1884_ _1947_ sg13g2_o21ai_1
X_5002_ VGND VPWR _1000_ _0990_ net1653 sg13g2_or2_1
Xfanout1291 s0.valid_out\[7\][0] net1291 VPWR VGND sg13g2_buf_8
Xfanout1280 net1281 net1280 VPWR VGND sg13g2_buf_8
XFILLER_38_155 VPWR VGND sg13g2_fill_1
X_6953_ net1274 VPWR _2756_ VGND _2691_ _2755_ sg13g2_o21ai_1
X_6884_ VGND VPWR _2582_ _2693_ _2694_ net1274 sg13g2_a21oi_1
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
X_5904_ _1817_ _1811_ _1816_ VPWR VGND sg13g2_nand2_1
XFILLER_34_350 VPWR VGND sg13g2_fill_2
X_5835_ net1391 net1350 _1748_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_545 VPWR VGND sg13g2_fill_1
X_5766_ _1691_ net1411 s0.data_out\[14\]\[4\] VPWR VGND sg13g2_nand2_1
X_7505_ _3253_ net1220 _3254_ _3255_ VPWR VGND sg13g2_a21o_1
X_4717_ _0737_ VPWR _0738_ VGND net1182 _0735_ sg13g2_o21ai_1
X_5697_ net1196 VPWR _1625_ VGND s0.was_valid_out\[14\][0] net1421 sg13g2_o21ai_1
X_7436_ net1233 VPWR _3193_ VGND _3165_ _3192_ sg13g2_o21ai_1
X_4648_ _0661_ _0674_ _0676_ _0681_ VPWR VGND sg13g2_nor3_1
XFILLER_2_917 VPWR VGND sg13g2_decap_8
X_4579_ net1727 net375 _0147_ VPWR VGND sg13g2_and2_1
X_7367_ VGND VPWR _3129_ _3111_ net1571 sg13g2_or2_1
X_6318_ _0312_ _2185_ _2186_ _3495_ net1612 VPWR VGND sg13g2_a22oi_1
X_7298_ _3070_ VPWR _3071_ VGND net1718 net795 sg13g2_o21ai_1
X_6249_ _2126_ net1362 net522 VPWR VGND sg13g2_nand2_1
XFILLER_44_103 VPWR VGND sg13g2_fill_2
XFILLER_29_166 VPWR VGND sg13g2_fill_2
XFILLER_29_199 VPWR VGND sg13g2_fill_2
XFILLER_25_350 VPWR VGND sg13g2_decap_8
XFILLER_5_744 VPWR VGND sg13g2_fill_1
X_7920__87 VPWR VGND net87 sg13g2_tiehi
XFILLER_20_70 VPWR VGND sg13g2_fill_1
XFILLER_45_1005 VPWR VGND sg13g2_decap_8
XFILLER_1_950 VPWR VGND sg13g2_decap_8
X_7714__310 VPWR VGND net310 sg13g2_tiehi
XFILLER_49_976 VPWR VGND sg13g2_decap_8
Xhold90 s0.data_out\[0\]\[2\] VPWR VGND net459 sg13g2_dlygate4sd3_1
XFILLER_32_810 VPWR VGND sg13g2_fill_1
X_5620_ _1557_ net1420 s0.data_out\[15\]\[6\] VPWR VGND sg13g2_nand2_1
X_5551_ _1494_ VPWR _1495_ VGND net1207 _1493_ sg13g2_o21ai_1
X_4502_ VPWR _0547_ _0546_ VGND sg13g2_inv_1
X_5482_ _1412_ _1421_ _1422_ _1430_ _1431_ VPWR VGND sg13g2_nor4_1
X_7221_ VGND VPWR net1229 _2993_ _2995_ _2994_ sg13g2_a21oi_1
X_4433_ net1186 _3424_ _0482_ VPWR VGND sg13g2_nor2_1
X_4364_ _0421_ net834 net1557 VPWR VGND sg13g2_nand2b_1
X_7152_ net1241 net1333 _2938_ VPWR VGND sg13g2_nor2b_1
X_7951__360 VPWR VGND net360 sg13g2_tiehi
X_4295_ net1547 net452 _0360_ VPWR VGND sg13g2_and2_1
X_7083_ _2870_ _2871_ _2872_ VPWR VGND sg13g2_nor2_1
X_6103_ _1992_ net1376 _1991_ VPWR VGND sg13g2_nand2b_1
X_7834__180 VPWR VGND net180 sg13g2_tiehi
X_6034_ net373 net1568 _1934_ _0280_ VPWR VGND sg13g2_nor3_1
XFILLER_39_420 VPWR VGND sg13g2_fill_2
X_6936_ _2742_ VPWR _2743_ VGND net1725 net532 sg13g2_o21ai_1
XFILLER_23_876 VPWR VGND sg13g2_fill_1
X_6867_ _2677_ net1269 net693 VPWR VGND sg13g2_nand2_1
XFILLER_34_191 VPWR VGND sg13g2_fill_2
XFILLER_10_526 VPWR VGND sg13g2_fill_2
X_6798_ VGND VPWR net1177 _2562_ _2619_ net1598 sg13g2_a21oi_1
X_5818_ net1418 VPWR _1735_ VGND _1665_ _1734_ sg13g2_o21ai_1
X_5749_ _1674_ s0.data_out\[14\]\[6\] net1420 VPWR VGND sg13g2_nand2b_1
XFILLER_41_69 VPWR VGND sg13g2_fill_1
X_7419_ _3179_ VPWR _3180_ VGND net1719 net721 sg13g2_o21ai_1
XFILLER_49_239 VPWR VGND sg13g2_decap_4
XFILLER_18_604 VPWR VGND sg13g2_decap_4
XFILLER_46_946 VPWR VGND sg13g2_decap_8
XFILLER_45_445 VPWR VGND sg13g2_fill_2
XFILLER_14_832 VPWR VGND sg13g2_fill_1
XFILLER_25_191 VPWR VGND sg13g2_decap_4
XFILLER_41_684 VPWR VGND sg13g2_fill_1
XFILLER_5_563 VPWR VGND sg13g2_fill_1
X_7818__197 VPWR VGND net197 sg13g2_tiehi
X_4080_ VPWR _3456_ net709 VGND sg13g2_inv_1
XFILLER_49_773 VPWR VGND sg13g2_decap_8
XFILLER_37_968 VPWR VGND sg13g2_decap_8
X_4982_ VGND VPWR net1488 _0977_ _0980_ _0979_ sg13g2_a21oi_1
X_7770_ net249 VGND VPWR net467 s0.data_out\[16\]\[3\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_6721_ _2543_ net1278 net532 VPWR VGND sg13g2_nand2_1
X_6652_ net1286 net1344 _2486_ VPWR VGND sg13g2_nor2b_1
X_5603_ VPWR VGND _1539_ net1711 _1537_ net1706 _1540_ _1532_ sg13g2_a221oi_1
X_6583_ VPWR _0342_ _2421_ VGND sg13g2_inv_1
XFILLER_11_17 VPWR VGND sg13g2_fill_2
X_5534_ _1481_ VPWR _1482_ VGND net1743 net689 sg13g2_o21ai_1
X_5465_ _1413_ VPWR _1414_ VGND net1435 _3464_ sg13g2_o21ai_1
X_4416_ net1186 _3422_ _0469_ VPWR VGND sg13g2_nor2_1
X_7204_ net1585 _2935_ _2982_ VPWR VGND sg13g2_nor2_1
X_5396_ _1335_ _1350_ _1351_ _1357_ VPWR VGND sg13g2_nor3_1
X_7135_ _2921_ net1245 net616 VPWR VGND sg13g2_nand2_1
X_4347_ _3581_ VPWR _0404_ VGND net1557 _3420_ sg13g2_o21ai_1
X_4278_ _3613_ _3614_ _0347_ VPWR VGND sg13g2_nor2_1
X_7066_ _0044_ _2857_ _2858_ _3527_ net1597 VPWR VGND sg13g2_a22oi_1
X_6017_ _1918_ net1387 net540 VPWR VGND sg13g2_nand2_1
XFILLER_36_36 VPWR VGND sg13g2_fill_1
XFILLER_36_69 VPWR VGND sg13g2_fill_1
X_7968_ net119 VGND VPWR _0102_ s0.data_out\[0\]\[2\] clknet_leaf_11_clk sg13g2_dfrbpq_2
XFILLER_43_949 VPWR VGND sg13g2_decap_8
XFILLER_14_128 VPWR VGND sg13g2_fill_2
X_7899_ net110 VGND VPWR _0033_ s0.data_out\[6\]\[5\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_6919_ VGND VPWR _2714_ _2722_ _2729_ _2706_ sg13g2_a21oi_1
XFILLER_35_1004 VPWR VGND sg13g2_decap_8
XFILLER_10_301 VPWR VGND sg13g2_fill_1
X_7704__320 VPWR VGND net320 sg13g2_tiehi
XFILLER_22_183 VPWR VGND sg13g2_fill_2
XFILLER_7_828 VPWR VGND sg13g2_fill_1
XFILLER_10_345 VPWR VGND sg13g2_decap_8
Xhold390 s0.data_out\[22\]\[0\] VPWR VGND net759 sg13g2_dlygate4sd3_1
X_7711__313 VPWR VGND net313 sg13g2_tiehi
XFILLER_46_765 VPWR VGND sg13g2_decap_8
XFILLER_45_253 VPWR VGND sg13g2_fill_1
XFILLER_19_979 VPWR VGND sg13g2_decap_8
XFILLER_34_927 VPWR VGND sg13g2_fill_1
XFILLER_42_982 VPWR VGND sg13g2_decap_8
XFILLER_14_673 VPWR VGND sg13g2_fill_1
X_7824__190 VPWR VGND net190 sg13g2_tiehi
XFILLER_9_165 VPWR VGND sg13g2_fill_1
X_5250_ _1223_ _1222_ net1654 _1215_ net1664 VPWR VGND sg13g2_a22oi_1
X_4201_ _3564_ VPWR _3565_ VGND net1555 _3413_ sg13g2_o21ai_1
X_5181_ net1473 VPWR _1160_ VGND _1127_ _1159_ sg13g2_o21ai_1
X_4132_ VPWR _3508_ net608 VGND sg13g2_inv_1
XFILLER_49_570 VPWR VGND sg13g2_decap_8
X_4063_ VPWR _3439_ net530 VGND sg13g2_inv_1
X_7831__183 VPWR VGND net183 sg13g2_tiehi
X_7822_ net193 VGND VPWR net541 s0.data_out\[12\]\[7\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_7948__57 VPWR VGND net57 sg13g2_tiehi
X_4965_ _0963_ net1178 _0962_ VPWR VGND sg13g2_nand2_1
X_7753_ net267 VGND VPWR _0231_ s0.genblk1\[16\].modules.bubble clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_6704_ net1176 _3517_ _2530_ VPWR VGND sg13g2_nor2_1
X_7684_ net342 VGND VPWR net817 s0.data_out\[23\]\[1\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_4896_ net1690 _0864_ _0905_ VPWR VGND sg13g2_nor2_1
X_6635_ net1286 net1337 _2469_ VPWR VGND sg13g2_nor2b_1
X_6566_ net1306 VPWR _2408_ VGND _2345_ _2407_ sg13g2_o21ai_1
X_5517_ _1336_ VPWR _1466_ VGND net1445 _3468_ sg13g2_o21ai_1
X_6497_ _2343_ net1302 net547 VPWR VGND sg13g2_nand2_1
X_5448_ net1623 _1391_ _1392_ _0230_ VPWR VGND sg13g2_nor3_1
X_5379_ _1340_ net681 net1455 VPWR VGND sg13g2_nand2b_1
X_7118_ _2904_ s0.data_out\[3\]\[3\] net1254 VPWR VGND sg13g2_nand2b_1
X_7049_ _2845_ VPWR _2846_ VGND net1726 net618 sg13g2_o21ai_1
XFILLER_31_908 VPWR VGND sg13g2_fill_1
XFILLER_8_29 VPWR VGND sg13g2_fill_1
XFILLER_24_993 VPWR VGND sg13g2_decap_8
XFILLER_12_71 VPWR VGND sg13g2_fill_2
X_7778__240 VPWR VGND net240 sg13g2_tiehi
XFILLER_3_886 VPWR VGND sg13g2_decap_8
Xfanout1621 net1625 net1621 VPWR VGND sg13g2_buf_8
Xfanout1632 _3374_ net1632 VPWR VGND sg13g2_buf_8
Xfanout1610 net1615 net1610 VPWR VGND sg13g2_buf_8
Xfanout1643 net1646 net1643 VPWR VGND sg13g2_buf_8
Xfanout1654 net1656 net1654 VPWR VGND sg13g2_buf_8
Xfanout1665 net1666 net1665 VPWR VGND sg13g2_buf_8
Xfanout1676 ui_in[5] net1676 VPWR VGND sg13g2_buf_8
Xfanout1698 net1700 net1698 VPWR VGND sg13g2_buf_1
Xfanout1687 net1689 net1687 VPWR VGND sg13g2_buf_8
XFILLER_19_743 VPWR VGND sg13g2_fill_1
X_7785__233 VPWR VGND net233 sg13g2_tiehi
XFILLER_15_982 VPWR VGND sg13g2_decap_8
X_4750_ _0771_ net1505 s0.data_out\[22\]\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_33_289 VPWR VGND sg13g2_fill_1
X_4681_ _0155_ _0705_ _0706_ _3426_ net1593 VPWR VGND sg13g2_a22oi_1
X_6420_ _2251_ _2253_ _2278_ VPWR VGND sg13g2_nor2b_1
X_6351_ _2209_ net485 net1360 VPWR VGND sg13g2_nand2b_1
X_5302_ _1268_ VPWR _1269_ VGND net1199 _1267_ sg13g2_o21ai_1
XFILLER_45_0 VPWR VGND sg13g2_fill_2
X_6282_ VPWR VGND _2158_ _2080_ _2153_ _2134_ _2159_ _2136_ sg13g2_a221oi_1
X_5233_ VGND VPWR net1463 _1203_ _1206_ _1205_ sg13g2_a21oi_1
X_5164_ net1198 _3456_ _1147_ VPWR VGND sg13g2_nor2_1
X_4115_ _3491_ net513 VPWR VGND sg13g2_inv_2
X_5095_ _1080_ _3392_ s0.data_out\[19\]\[1\] VPWR VGND sg13g2_nand2_1
X_4046_ VPWR _3422_ net501 VGND sg13g2_inv_1
X_7805_ net211 VGND VPWR _0283_ s0.data_out\[13\]\[2\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_5997_ VGND VPWR net1392 _1895_ _1898_ _1897_ sg13g2_a21oi_1
XFILLER_13_919 VPWR VGND sg13g2_fill_2
XFILLER_24_278 VPWR VGND sg13g2_fill_2
X_7736_ net286 VGND VPWR _0214_ s0.data_out\[19\]\[5\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_4948_ _0948_ _0945_ _0947_ VPWR VGND sg13g2_nand2_1
X_7667_ net361 VGND VPWR _0145_ s0.was_valid_out\[24\][0] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_4879_ net1482 net1340 _0888_ VPWR VGND sg13g2_nor2b_1
X_6618_ VGND VPWR net1282 _2450_ _2452_ _2451_ sg13g2_a21oi_1
X_7598_ net1696 _3335_ _3336_ VPWR VGND sg13g2_nor2_1
X_6549_ _2312_ _2393_ _2394_ _2395_ VPWR VGND sg13g2_nor3_1
XFILLER_3_116 VPWR VGND sg13g2_fill_1
XFILLER_0_845 VPWR VGND sg13g2_decap_8
XFILLER_48_816 VPWR VGND sg13g2_decap_8
XFILLER_16_724 VPWR VGND sg13g2_fill_1
XFILLER_28_573 VPWR VGND sg13g2_fill_2
X_7935__71 VPWR VGND net71 sg13g2_tiehi
XFILLER_12_996 VPWR VGND sg13g2_decap_8
XFILLER_8_989 VPWR VGND sg13g2_decap_8
XFILLER_23_92 VPWR VGND sg13g2_fill_2
XFILLER_39_827 VPWR VGND sg13g2_fill_1
XFILLER_38_304 VPWR VGND sg13g2_fill_1
Xfanout1440 net1441 net1440 VPWR VGND sg13g2_buf_8
Xfanout1451 net1452 net1451 VPWR VGND sg13g2_buf_8
Xfanout1484 net1485 net1484 VPWR VGND sg13g2_buf_1
Xfanout1473 net1476 net1473 VPWR VGND sg13g2_buf_8
Xfanout1462 net1463 net1462 VPWR VGND sg13g2_buf_1
Xfanout1495 net1497 net1495 VPWR VGND sg13g2_buf_8
XFILLER_19_540 VPWR VGND sg13g2_decap_4
XFILLER_47_871 VPWR VGND sg13g2_decap_8
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
X_5920_ net1627 _1751_ _1830_ VPWR VGND sg13g2_nor2_1
XFILLER_46_392 VPWR VGND sg13g2_fill_2
X_5851_ _1764_ net1402 _1763_ VPWR VGND sg13g2_nand2b_1
X_4802_ _0816_ VPWR _0817_ VGND net1727 net610 sg13g2_o21ai_1
X_5782_ VGND VPWR _1707_ net1568 net396 sg13g2_or2_1
X_7521_ net1211 net1343 _3271_ VPWR VGND sg13g2_nor2b_1
X_4733_ s0.data_out\[23\]\[7\] s0.data_out\[22\]\[7\] net1503 _0754_ VPWR VGND sg13g2_mux2_1
X_7452_ _0083_ _3204_ _3205_ _3538_ net1584 VPWR VGND sg13g2_a22oi_1
X_4664_ net1589 _0617_ _0694_ VPWR VGND sg13g2_nor2_1
X_6403_ _2261_ _2260_ net1320 VPWR VGND sg13g2_nand2b_1
X_4595_ net1510 net1357 _0628_ VPWR VGND sg13g2_nor2b_1
X_7383_ s0.data_out\[2\]\[7\] s0.data_out\[1\]\[7\] net1224 _3145_ VPWR VGND sg13g2_mux2_1
X_6334_ net1638 net1352 _2199_ VPWR VGND sg13g2_nor2_1
X_6265_ VGND VPWR _2033_ _2141_ _2142_ net1366 sg13g2_a21oi_1
X_5216_ _1189_ s0.data_out\[18\]\[1\] net1465 VPWR VGND sg13g2_nand2b_1
X_6196_ _0300_ _2075_ _2076_ _3487_ net1613 VPWR VGND sg13g2_a22oi_1
X_5147_ net1673 _1131_ _1132_ VPWR VGND sg13g2_nor2_1
XFILLER_29_304 VPWR VGND sg13g2_fill_1
X_5078_ _1064_ _1065_ _1066_ VPWR VGND sg13g2_nor2_1
X_4029_ VPWR _3405_ net461 VGND sg13g2_inv_1
XFILLER_13_716 VPWR VGND sg13g2_fill_2
X_7719_ net304 VGND VPWR _0197_ s0.data_out\[20\]\[0\] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_20_281 VPWR VGND sg13g2_fill_1
X_7932__74 VPWR VGND net74 sg13g2_tiehi
XFILLER_5_937 VPWR VGND sg13g2_decap_8
XFILLER_0_631 VPWR VGND sg13g2_decap_8
XFILLER_48_624 VPWR VGND sg13g2_fill_1
XFILLER_48_613 VPWR VGND sg13g2_decap_8
XFILLER_16_510 VPWR VGND sg13g2_fill_1
X_7782__236 VPWR VGND net236 sg13g2_tiehi
XFILLER_31_513 VPWR VGND sg13g2_decap_4
XFILLER_15_1024 VPWR VGND sg13g2_decap_4
Xhold208 s0.data_out\[13\]\[1\] VPWR VGND net577 sg13g2_dlygate4sd3_1
X_4380_ s0.data_out\[26\]\[4\] s0.data_out\[25\]\[4\] net1540 _0437_ VPWR VGND sg13g2_mux2_1
Xhold219 s0.data_out\[14\]\[4\] VPWR VGND net588 sg13g2_dlygate4sd3_1
X_6050_ net1385 net597 _1947_ VPWR VGND sg13g2_and2_1
X_5001_ net1663 _0997_ _0999_ VPWR VGND sg13g2_nor2_1
Xfanout1292 s0.valid_out\[7\][0] net1292 VPWR VGND sg13g2_buf_8
Xfanout1281 s0.valid_out\[6\][0] net1281 VPWR VGND sg13g2_buf_8
XFILLER_38_145 VPWR VGND sg13g2_fill_1
Xfanout1270 net1272 net1270 VPWR VGND sg13g2_buf_8
X_6952_ net1263 net584 _2755_ VPWR VGND sg13g2_and2_1
XFILLER_35_841 VPWR VGND sg13g2_decap_4
X_6883_ _2693_ net584 net1280 VPWR VGND sg13g2_nand2b_1
XFILLER_34_340 VPWR VGND sg13g2_fill_2
X_5903_ _3406_ _1803_ _1812_ _1816_ VPWR VGND sg13g2_or3_1
X_5834_ s0.data_out\[14\]\[2\] s0.data_out\[13\]\[2\] net1398 _1747_ VPWR VGND sg13g2_mux2_1
XFILLER_34_395 VPWR VGND sg13g2_fill_2
X_5765_ net1404 net1345 _1690_ VPWR VGND sg13g2_nor2b_1
X_7504_ net1220 _3250_ _3254_ VPWR VGND sg13g2_nor2_1
X_4716_ _0737_ net1183 _0736_ VPWR VGND sg13g2_nand2_1
X_5696_ net1405 _1619_ _1624_ VPWR VGND sg13g2_nor2_1
X_7435_ net1221 s0.data_out\[1\]\[4\] _3192_ VPWR VGND sg13g2_and2_1
X_4647_ _0643_ _0661_ _0679_ _0680_ VPWR VGND sg13g2_or3_1
X_7366_ VPWR VGND _3126_ _3127_ _3119_ net1571 _3128_ _3111_ sg13g2_a221oi_1
X_6317_ net1612 _2131_ _2186_ VPWR VGND sg13g2_nor2_1
X_4578_ net1592 _0606_ _0146_ VPWR VGND sg13g2_nor2_1
XFILLER_1_439 VPWR VGND sg13g2_fill_2
X_7297_ _3069_ VPWR _3070_ VGND net1190 _3068_ sg13g2_o21ai_1
X_6248_ VGND VPWR net1369 _2122_ _2125_ _2124_ sg13g2_a21oi_1
XFILLER_39_69 VPWR VGND sg13g2_fill_2
X_6179_ _3383_ _3497_ _2063_ VPWR VGND sg13g2_nor2_1
XFILLER_17_318 VPWR VGND sg13g2_fill_1
XFILLER_9_506 VPWR VGND sg13g2_decap_4
XFILLER_40_398 VPWR VGND sg13g2_decap_4
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_955 VPWR VGND sg13g2_decap_8
XFILLER_36_605 VPWR VGND sg13g2_fill_1
Xhold80 _3589_ VPWR VGND net449 sg13g2_dlygate4sd3_1
Xhold91 s0.shift_out\[17\][0] VPWR VGND net460 sg13g2_dlygate4sd3_1
XFILLER_17_885 VPWR VGND sg13g2_decap_4
X_5550_ VGND VPWR net1207 _1466_ _1494_ net1622 sg13g2_a21oi_1
XFILLER_8_583 VPWR VGND sg13g2_fill_2
X_4501_ VGND VPWR _0546_ _0536_ net1647 sg13g2_or2_1
X_5481_ net1692 _1429_ _1430_ VPWR VGND sg13g2_nor2_1
X_4432_ VPWR _0131_ _0481_ VGND sg13g2_inv_1
X_7220_ net1228 net1352 _2994_ VPWR VGND sg13g2_nor2b_1
X_4363_ _0418_ net1533 _0419_ _0420_ VPWR VGND sg13g2_a21o_1
X_7151_ s0.data_out\[4\]\[6\] s0.data_out\[3\]\[6\] net1246 _2937_ VPWR VGND sg13g2_mux2_1
X_4294_ _0115_ _0358_ _0359_ _3413_ net1576 VPWR VGND sg13g2_a22oi_1
X_7082_ net1249 _2762_ _2871_ VPWR VGND sg13g2_nor2_1
X_6102_ VGND VPWR net1367 _1989_ _1991_ _1990_ sg13g2_a21oi_1
X_6033_ VPWR VGND _1929_ _1933_ _1932_ _1891_ _1934_ _1931_ sg13g2_a221oi_1
XFILLER_6_1022 VPWR VGND sg13g2_decap_8
X_6935_ _2741_ VPWR _2742_ VGND net1175 _2740_ sg13g2_o21ai_1
XFILLER_25_49 VPWR VGND sg13g2_fill_1
X_6866_ _2676_ net1572 _2674_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_505 VPWR VGND sg13g2_decap_8
X_6797_ VGND VPWR net1271 s0.data_out\[6\]\[0\] _2618_ _2559_ sg13g2_a21oi_1
X_5817_ net1195 _3476_ _1734_ VPWR VGND sg13g2_nor2_1
X_5748_ _1671_ net1405 _1672_ _1673_ VPWR VGND sg13g2_a21o_1
X_5679_ net1427 VPWR _1610_ VGND _1577_ _1609_ sg13g2_o21ai_1
X_7418_ _3178_ VPWR _3179_ VGND net1187 _3177_ sg13g2_o21ai_1
X_7349_ _3110_ VPWR _3111_ VGND net1189 _3108_ sg13g2_o21ai_1
XFILLER_49_229 VPWR VGND sg13g2_fill_1
XFILLER_46_925 VPWR VGND sg13g2_decap_8
XFILLER_18_638 VPWR VGND sg13g2_fill_2
XFILLER_41_630 VPWR VGND sg13g2_fill_1
XFILLER_13_376 VPWR VGND sg13g2_fill_1
XFILLER_14_888 VPWR VGND sg13g2_fill_2
XFILLER_49_7 VPWR VGND sg13g2_decap_8
Xoutput2 net2 uio_out[2] VPWR VGND sg13g2_buf_1
XFILLER_49_752 VPWR VGND sg13g2_decap_8
XFILLER_45_991 VPWR VGND sg13g2_decap_8
X_4981_ VGND VPWR _0859_ _0978_ _0979_ net1486 sg13g2_a21oi_1
X_6720_ net1729 net386 _0014_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_43_clk clknet_3_0__leaf_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
X_6651_ s0.data_out\[8\]\[4\] s0.data_out\[7\]\[4\] net1292 _2485_ VPWR VGND sg13g2_mux2_1
X_6582_ _2420_ VPWR _2421_ VGND net1731 net731 sg13g2_o21ai_1
X_5602_ _1539_ _1538_ net1424 VPWR VGND sg13g2_nand2b_1
X_5533_ _1480_ VPWR _1481_ VGND net1206 _1479_ sg13g2_o21ai_1
X_5464_ _1413_ net1435 net655 VPWR VGND sg13g2_nand2_1
X_5395_ _1335_ _1354_ _1355_ _1356_ VPWR VGND sg13g2_or3_1
X_4415_ _0127_ _0467_ _0468_ _3412_ net1578 VPWR VGND sg13g2_a22oi_1
X_7203_ net1248 VPWR _2981_ VGND _2932_ _2980_ sg13g2_o21ai_1
X_4346_ _0403_ net1552 _0402_ VPWR VGND sg13g2_nand2b_1
X_7134_ net1242 net1343 _2920_ VPWR VGND sg13g2_nor2b_1
X_4277_ VGND VPWR _3625_ _0345_ _0346_ _3616_ sg13g2_a21oi_1
X_7065_ net1596 _2824_ _2858_ VPWR VGND sg13g2_nor2_1
X_6016_ VGND VPWR net1392 _1914_ _1917_ _1916_ sg13g2_a21oi_1
XFILLER_36_15 VPWR VGND sg13g2_fill_2
XFILLER_27_457 VPWR VGND sg13g2_decap_4
XFILLER_43_928 VPWR VGND sg13g2_decap_8
X_7967_ net132 VGND VPWR _0101_ s0.data_out\[0\]\[1\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_6918_ _2727_ VPWR _2728_ VGND _2686_ _2688_ sg13g2_o21ai_1
X_7898_ net111 VGND VPWR _0032_ s0.data_out\[6\]\[4\] clknet_leaf_16_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_34_clk clknet_3_4__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
X_6849_ VGND VPWR _2551_ _2658_ _2659_ net1270 sg13g2_a21oi_1
Xhold380 _0000_ VPWR VGND net749 sg13g2_dlygate4sd3_1
Xhold391 s0.data_out\[11\]\[3\] VPWR VGND net760 sg13g2_dlygate4sd3_1
XFILLER_46_744 VPWR VGND sg13g2_decap_8
XFILLER_26_70 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_25_clk clknet_3_7__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_42_961 VPWR VGND sg13g2_decap_8
XFILLER_13_151 VPWR VGND sg13g2_fill_2
XFILLER_9_155 VPWR VGND sg13g2_fill_2
X_4200_ _3564_ net1555 net464 VPWR VGND sg13g2_nand2_1
X_5180_ net1457 s0.data_out\[19\]\[5\] _1159_ VPWR VGND sg13g2_and2_1
X_4131_ VPWR _3507_ net561 VGND sg13g2_inv_1
X_4062_ VPWR _3438_ net552 VGND sg13g2_inv_1
X_7821_ net194 VGND VPWR _0299_ s0.data_out\[12\]\[6\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_7752_ net268 VGND VPWR _0230_ s0.valid_out\[17\][0] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_4964_ _0843_ VPWR _0962_ VGND net1492 _3450_ sg13g2_o21ai_1
Xclkbuf_leaf_16_clk clknet_3_3__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_6703_ _0010_ _2528_ _2529_ _3508_ net1600 VPWR VGND sg13g2_a22oi_1
X_4895_ VGND VPWR _0890_ _0892_ _0904_ net1673 sg13g2_a21oi_1
X_7683_ net343 VGND VPWR _0161_ s0.data_out\[23\]\[0\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_6634_ s0.data_out\[8\]\[6\] s0.data_out\[7\]\[6\] net1292 _2468_ VPWR VGND sg13g2_mux2_1
XFILLER_20_666 VPWR VGND sg13g2_fill_2
X_6565_ _3394_ _3511_ _2407_ VPWR VGND sg13g2_nor2_1
X_5516_ _1465_ net1442 _1464_ VPWR VGND sg13g2_nand2b_1
X_6496_ _2326_ _2340_ _2341_ _2342_ VPWR VGND sg13g2_nor3_1
X_5447_ VGND VPWR _3366_ _1393_ _0229_ _1398_ sg13g2_a21oi_1
X_5378_ _1337_ net1439 _1338_ _1339_ VPWR VGND sg13g2_a21o_1
X_4329_ s0.data_out\[26\]\[2\] s0.data_out\[25\]\[2\] net1541 _0386_ VPWR VGND sg13g2_mux2_1
X_7117_ _2901_ net1242 _2902_ _2903_ VPWR VGND sg13g2_a21o_1
X_7048_ _2790_ _2844_ net1726 _2845_ VPWR VGND sg13g2_nand3_1
XFILLER_47_58 VPWR VGND sg13g2_fill_1
XFILLER_28_755 VPWR VGND sg13g2_fill_1
XFILLER_15_438 VPWR VGND sg13g2_fill_2
XFILLER_24_972 VPWR VGND sg13g2_decap_8
XFILLER_11_655 VPWR VGND sg13g2_fill_1
XFILLER_3_865 VPWR VGND sg13g2_decap_8
XFILLER_2_331 VPWR VGND sg13g2_fill_2
Xfanout1600 net1601 net1600 VPWR VGND sg13g2_buf_8
Xfanout1633 net1636 net1633 VPWR VGND sg13g2_buf_8
Xfanout1622 net1625 net1622 VPWR VGND sg13g2_buf_8
Xfanout1611 net1614 net1611 VPWR VGND sg13g2_buf_8
Xfanout1644 net1646 net1644 VPWR VGND sg13g2_buf_8
Xfanout1666 net1667 net1666 VPWR VGND sg13g2_buf_8
Xfanout1655 net1656 net1655 VPWR VGND sg13g2_buf_8
XFILLER_19_8 VPWR VGND sg13g2_fill_2
Xfanout1699 net1700 net1699 VPWR VGND sg13g2_buf_8
Xfanout1688 net1689 net1688 VPWR VGND sg13g2_buf_8
Xfanout1677 net1681 net1677 VPWR VGND sg13g2_buf_8
XFILLER_46_530 VPWR VGND sg13g2_fill_2
X_4680_ net1593 _0656_ _0706_ VPWR VGND sg13g2_nor2_1
XFILLER_14_493 VPWR VGND sg13g2_decap_4
XFILLER_30_986 VPWR VGND sg13g2_decap_8
X_6350_ _2206_ net1307 _2207_ _2208_ VPWR VGND sg13g2_a21o_1
X_5301_ VGND VPWR net1199 _1232_ _1268_ net1618 sg13g2_a21oi_1
X_6281_ _2137_ _2152_ _2158_ VPWR VGND sg13g2_nor2b_1
X_5232_ VGND VPWR _1091_ _1204_ _1205_ net1463 sg13g2_a21oi_1
Xclkbuf_leaf_5_clk clknet_3_1__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
XFILLER_38_0 VPWR VGND sg13g2_decap_4
X_5163_ VPWR _0197_ _1146_ VGND sg13g2_inv_1
XFILLER_29_508 VPWR VGND sg13g2_fill_2
X_4114_ VPWR _3490_ net789 VGND sg13g2_inv_1
X_5094_ _1077_ net1458 _1078_ _1079_ VPWR VGND sg13g2_a21o_1
XFILLER_49_390 VPWR VGND sg13g2_decap_4
X_4045_ VPWR _3421_ net707 VGND sg13g2_inv_1
XFILLER_13_909 VPWR VGND sg13g2_fill_1
X_7804_ net212 VGND VPWR _0282_ s0.data_out\[13\]\[1\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_5996_ VGND VPWR _1797_ _1896_ _1897_ net1391 sg13g2_a21oi_1
X_7944__61 VPWR VGND net61 sg13g2_tiehi
X_4947_ net1180 VPWR _0947_ VGND s0.was_valid_out\[20\][0] net1489 sg13g2_o21ai_1
X_7735_ net287 VGND VPWR net500 s0.data_out\[19\]\[4\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_4878_ s0.data_out\[22\]\[5\] s0.data_out\[21\]\[5\] net1490 _0887_ VPWR VGND sg13g2_mux2_1
X_7666_ net362 VGND VPWR _0144_ s0.data_out\[25\]\[7\] clknet_leaf_44_clk sg13g2_dfrbpq_2
X_6617_ net1283 net1359 _2451_ VPWR VGND sg13g2_nor2b_1
X_7597_ _3334_ VPWR _3335_ VGND _3393_ net1348 sg13g2_o21ai_1
X_7701__324 VPWR VGND net324 sg13g2_tiehi
X_6548_ _2365_ _2366_ _2394_ VPWR VGND sg13g2_nor2b_1
X_6479_ VGND VPWR net1305 _2322_ _2325_ _2324_ sg13g2_a21oi_1
XFILLER_0_824 VPWR VGND sg13g2_decap_8
XFILLER_28_585 VPWR VGND sg13g2_fill_2
XFILLER_15_268 VPWR VGND sg13g2_decap_8
XFILLER_8_913 VPWR VGND sg13g2_fill_2
X_7950__42 VPWR VGND net42 sg13g2_tiehi
XFILLER_7_412 VPWR VGND sg13g2_fill_1
XFILLER_23_82 VPWR VGND sg13g2_fill_2
X_7821__194 VPWR VGND net194 sg13g2_tiehi
XFILLER_8_968 VPWR VGND sg13g2_decap_8
XFILLER_7_467 VPWR VGND sg13g2_fill_2
XFILLER_7_434 VPWR VGND sg13g2_fill_1
XFILLER_48_1026 VPWR VGND sg13g2_fill_2
XFILLER_39_817 VPWR VGND sg13g2_fill_2
Xfanout1441 net1442 net1441 VPWR VGND sg13g2_buf_8
Xfanout1430 net1431 net1430 VPWR VGND sg13g2_buf_8
Xfanout1474 net1476 net1474 VPWR VGND sg13g2_buf_1
Xfanout1452 net475 net1452 VPWR VGND sg13g2_buf_8
Xfanout1463 s0.shift_out\[19\][0] net1463 VPWR VGND sg13g2_buf_8
XFILLER_47_850 VPWR VGND sg13g2_decap_8
XFILLER_38_349 VPWR VGND sg13g2_decap_4
Xfanout1485 net477 net1485 VPWR VGND sg13g2_buf_2
Xfanout1496 net1497 net1496 VPWR VGND sg13g2_buf_1
XFILLER_0_1006 VPWR VGND sg13g2_decap_8
XFILLER_0_64 VPWR VGND sg13g2_fill_2
XFILLER_19_585 VPWR VGND sg13g2_fill_2
X_5850_ VGND VPWR net1390 _1761_ _1763_ _1762_ sg13g2_a21oi_1
X_4801_ _0815_ VPWR _0816_ VGND net1183 _0814_ sg13g2_o21ai_1
X_5781_ VGND VPWR _1700_ _1704_ _1706_ _1705_ sg13g2_a21oi_1
X_7520_ s0.data_out\[1\]\[4\] s0.data_out\[0\]\[4\] net1215 _3270_ VPWR VGND sg13g2_mux2_1
X_4732_ _0753_ net1505 net558 VPWR VGND sg13g2_nand2_1
XFILLER_30_750 VPWR VGND sg13g2_fill_2
X_4663_ net1525 VPWR _0693_ VGND _0614_ _0692_ sg13g2_o21ai_1
X_7451_ net1582 _3149_ _3205_ VPWR VGND sg13g2_nor2_1
X_7941__64 VPWR VGND net64 sg13g2_tiehi
X_6402_ s0.data_out\[9\]\[4\] s0.data_out\[10\]\[4\] net1360 _2260_ VPWR VGND sg13g2_mux2_1
X_4594_ s0.data_out\[24\]\[0\] s0.data_out\[23\]\[0\] net1515 _0627_ VPWR VGND sg13g2_mux2_1
X_7382_ VGND VPWR net1230 _3141_ _3144_ _3143_ sg13g2_a21oi_1
XFILLER_7_990 VPWR VGND sg13g2_decap_8
X_6333_ VGND VPWR net1638 net1570 _0315_ _2198_ sg13g2_a21oi_1
X_6264_ _2141_ net747 net1372 VPWR VGND sg13g2_nand2b_1
X_5215_ _1186_ net1447 _1187_ _1188_ VPWR VGND sg13g2_a21o_1
X_6195_ net1613 _2018_ _2076_ VPWR VGND sg13g2_nor2_1
X_5146_ VGND VPWR net1473 _1128_ _1131_ _1130_ sg13g2_a21oi_1
X_5077_ VGND VPWR _3367_ _3392_ _1065_ net1473 sg13g2_a21oi_1
X_4028_ VPWR _3404_ net491 VGND sg13g2_inv_1
X_7768__251 VPWR VGND net251 sg13g2_tiehi
X_5979_ VGND VPWR _1869_ _1871_ _1880_ net1708 sg13g2_a21oi_1
X_7718_ net305 VGND VPWR _0196_ s0.shift_out\[20\][0] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_7649_ net36 VGND VPWR net465 s0.data_out\[26\]\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_2
XFILLER_5_916 VPWR VGND sg13g2_decap_8
X_7775__244 VPWR VGND net244 sg13g2_tiehi
XFILLER_0_610 VPWR VGND sg13g2_decap_8
XFILLER_0_698 VPWR VGND sg13g2_decap_8
XFILLER_48_669 VPWR VGND sg13g2_decap_8
XFILLER_43_330 VPWR VGND sg13g2_fill_1
XFILLER_44_897 VPWR VGND sg13g2_decap_8
XFILLER_15_1003 VPWR VGND sg13g2_decap_8
Xhold209 s0.was_valid_out\[24\][0] VPWR VGND net578 sg13g2_dlygate4sd3_1
X_5000_ _0998_ _0997_ net1663 _0990_ net1653 VPWR VGND sg13g2_a22oi_1
Xfanout1260 net1261 net1260 VPWR VGND sg13g2_buf_2
Xfanout1282 net1283 net1282 VPWR VGND sg13g2_buf_8
Xfanout1271 net1272 net1271 VPWR VGND sg13g2_buf_1
Xfanout1293 net1294 net1293 VPWR VGND sg13g2_buf_2
X_6951_ VPWR _0033_ _2754_ VGND sg13g2_inv_1
XFILLER_19_393 VPWR VGND sg13g2_decap_4
X_6882_ _2690_ net1264 _2691_ _2692_ VPWR VGND sg13g2_a21o_1
X_5902_ _1796_ _1812_ _1813_ _1814_ _1815_ VPWR VGND sg13g2_nor4_1
X_5833_ _1746_ net1397 s0.data_out\[13\]\[2\] VPWR VGND sg13g2_nand2_1
X_7503_ VGND VPWR net1209 _3251_ _3253_ _3252_ sg13g2_a21oi_1
X_5764_ _1686_ _1688_ net1675 _1689_ VPWR VGND sg13g2_nand3_1
X_4715_ s0.data_out\[22\]\[2\] s0.data_out\[23\]\[2\] net1517 _0736_ VPWR VGND sg13g2_mux2_1
X_5695_ _1621_ VPWR _1623_ VGND s0.was_valid_out\[14\][0] net1410 sg13g2_o21ai_1
X_7434_ _0079_ _3190_ _3191_ _3540_ net1587 VPWR VGND sg13g2_a22oi_1
X_4646_ _0679_ _0674_ _0678_ VPWR VGND sg13g2_nand2_1
X_4577_ VGND VPWR _0608_ _0611_ _0145_ _0612_ sg13g2_a21oi_1
X_7365_ VGND VPWR _3116_ _3118_ _3127_ net1702 sg13g2_a21oi_1
X_6316_ net1368 VPWR _2185_ VGND _2128_ _2184_ sg13g2_o21ai_1
X_7296_ VGND VPWR net1190 _3003_ _3069_ net1582 sg13g2_a21oi_1
X_6247_ VGND VPWR _2006_ _2123_ _2124_ net1368 sg13g2_a21oi_1
X_6178_ _0296_ _2061_ _2062_ _3489_ net1613 VPWR VGND sg13g2_a22oi_1
X_5129_ _1114_ _1113_ net1654 _1106_ net1664 VPWR VGND sg13g2_a22oi_1
XFILLER_44_138 VPWR VGND sg13g2_fill_2
XFILLER_41_801 VPWR VGND sg13g2_fill_1
XFILLER_38_1014 VPWR VGND sg13g2_decap_8
XFILLER_26_875 VPWR VGND sg13g2_fill_1
XFILLER_25_385 VPWR VGND sg13g2_fill_2
XFILLER_4_212 VPWR VGND sg13g2_fill_2
XFILLER_4_245 VPWR VGND sg13g2_fill_2
XFILLER_49_934 VPWR VGND sg13g2_decap_8
XFILLER_1_985 VPWR VGND sg13g2_decap_8
XFILLER_0_495 VPWR VGND sg13g2_decap_4
Xhold70 s0.data_out\[0\]\[5\] VPWR VGND net439 sg13g2_dlygate4sd3_1
Xhold81 s0.was_valid_out\[12\][0] VPWR VGND net450 sg13g2_dlygate4sd3_1
Xhold92 s0.data_out\[27\]\[5\] VPWR VGND net461 sg13g2_dlygate4sd3_1
XFILLER_45_91 VPWR VGND sg13g2_fill_2
XFILLER_44_683 VPWR VGND sg13g2_decap_4
XFILLER_43_182 VPWR VGND sg13g2_fill_1
XFILLER_31_355 VPWR VGND sg13g2_fill_1
XFILLER_32_889 VPWR VGND sg13g2_fill_2
XFILLER_8_551 VPWR VGND sg13g2_fill_1
X_4500_ net1658 _0543_ _0545_ VPWR VGND sg13g2_nor2_1
X_5480_ VGND VPWR net1438 _1426_ _1429_ _1428_ sg13g2_a21oi_1
X_4431_ _0480_ VPWR _0481_ VGND net1714 net706 sg13g2_o21ai_1
X_4362_ net1533 net1333 _0419_ VPWR VGND sg13g2_nor2b_1
X_7150_ VGND VPWR net1248 _2933_ _2936_ _2935_ sg13g2_a21oi_1
X_4293_ net1576 _3563_ _0359_ VPWR VGND sg13g2_nor2_1
X_7081_ VGND VPWR net1633 net1246 _2870_ _2868_ sg13g2_a21oi_1
X_6101_ net1367 s0.data_new_delayed\[0\] _1990_ VPWR VGND sg13g2_nor2b_1
X_6032_ _1852_ VPWR _1933_ VGND _1925_ _1927_ sg13g2_o21ai_1
XFILLER_6_1001 VPWR VGND sg13g2_decap_8
XFILLER_39_444 VPWR VGND sg13g2_decap_4
XFILLER_20_0 VPWR VGND sg13g2_fill_2
X_6934_ VGND VPWR net1175 _2672_ _2741_ net1590 sg13g2_a21oi_1
XFILLER_26_149 VPWR VGND sg13g2_fill_1
X_7765__254 VPWR VGND net254 sg13g2_tiehi
XFILLER_34_160 VPWR VGND sg13g2_fill_2
X_6865_ VGND VPWR _2675_ _2674_ net1571 sg13g2_or2_1
XFILLER_34_193 VPWR VGND sg13g2_fill_1
X_6796_ VGND VPWR _2615_ _2616_ _0015_ _2617_ sg13g2_a21oi_1
X_5816_ VPWR _0263_ net773 VGND sg13g2_inv_1
X_5747_ net1405 net1335 _1672_ VPWR VGND sg13g2_nor2b_1
X_5678_ net1415 net644 _1609_ VPWR VGND sg13g2_and2_1
X_7417_ VGND VPWR net1187 _3123_ _3178_ net1582 sg13g2_a21oi_1
X_4629_ s0.data_out\[24\]\[4\] s0.data_out\[23\]\[4\] net1515 _0662_ VPWR VGND sg13g2_mux2_1
X_7956__295 VPWR VGND net295 sg13g2_tiehi
X_7348_ _3110_ net1188 _3109_ VPWR VGND sg13g2_nand2_1
XFILLER_2_749 VPWR VGND sg13g2_decap_8
X_7279_ _3052_ VPWR _3053_ VGND net1237 _3537_ sg13g2_o21ai_1
X_7772__247 VPWR VGND net247 sg13g2_tiehi
XFILLER_46_904 VPWR VGND sg13g2_decap_8
XFILLER_17_105 VPWR VGND sg13g2_fill_2
XFILLER_9_348 VPWR VGND sg13g2_decap_4
XFILLER_12_1017 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
Xoutput3 net3 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_49_731 VPWR VGND sg13g2_decap_8
XFILLER_1_782 VPWR VGND sg13g2_decap_8
XFILLER_45_970 VPWR VGND sg13g2_decap_8
X_4980_ _0978_ s0.data_out\[20\]\[3\] net1492 VPWR VGND sg13g2_nand2b_1
XFILLER_23_119 VPWR VGND sg13g2_fill_1
X_6650_ _2482_ _2483_ _2481_ _2484_ VPWR VGND sg13g2_nand3_1
XFILLER_32_664 VPWR VGND sg13g2_fill_2
X_6581_ _2419_ net1731 _2420_ VPWR VGND _2363_ sg13g2_nand3b_1
X_5601_ s0.data_out\[15\]\[0\] s0.data_out\[16\]\[0\] net1432 _1538_ VPWR VGND sg13g2_mux2_1
X_5532_ VGND VPWR net1206 _1406_ _1480_ net1620 sg13g2_a21oi_1
X_5463_ VPWR VGND _1411_ net1711 _1407_ net1706 _1412_ _1405_ sg13g2_a221oi_1
X_4414_ net1578 _0390_ _0468_ VPWR VGND sg13g2_nor2_1
X_5394_ _1353_ VPWR _1355_ VGND _1308_ _1317_ sg13g2_o21ai_1
X_7202_ net1191 _3535_ _2980_ VPWR VGND sg13g2_nor2_1
X_4345_ VGND VPWR net1535 _0400_ _0402_ _0401_ sg13g2_a21oi_1
X_7133_ _2915_ _2913_ net1668 _2919_ VPWR VGND sg13g2_a21o_1
XFILLER_28_1013 VPWR VGND sg13g2_decap_8
X_7064_ net1263 VPWR _2857_ VGND _2821_ _2856_ sg13g2_o21ai_1
X_4276_ _0345_ _3634_ _3635_ VPWR VGND sg13g2_nand2_1
X_6015_ VGND VPWR _1785_ _1915_ _1916_ net1392 sg13g2_a21oi_1
XFILLER_43_907 VPWR VGND sg13g2_decap_8
X_7966_ net145 VGND VPWR _0100_ s0.data_out\[0\]\[0\] clknet_leaf_10_clk sg13g2_dfrbpq_2
XFILLER_42_439 VPWR VGND sg13g2_fill_1
X_6917_ _2706_ _2723_ _2724_ _2725_ _2727_ VPWR VGND sg13g2_nor4_1
X_7897_ net112 VGND VPWR _0031_ s0.data_out\[6\]\[3\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_6848_ _2658_ s0.data_out\[5\]\[1\] net1278 VPWR VGND sg13g2_nand2b_1
XFILLER_11_848 VPWR VGND sg13g2_fill_2
X_6779_ _2601_ net1280 s0.data_out\[6\]\[5\] VPWR VGND sg13g2_nand2_1
Xhold370 _1959_ VPWR VGND net739 sg13g2_dlygate4sd3_1
Xhold381 s0.data_out\[2\]\[1\] VPWR VGND net750 sg13g2_dlygate4sd3_1
Xhold392 _0308_ VPWR VGND net761 sg13g2_dlygate4sd3_1
XFILLER_46_723 VPWR VGND sg13g2_decap_8
XFILLER_18_425 VPWR VGND sg13g2_fill_2
XFILLER_42_940 VPWR VGND sg13g2_decap_8
XFILLER_26_491 VPWR VGND sg13g2_fill_2
XFILLER_27_992 VPWR VGND sg13g2_decap_8
XFILLER_9_112 VPWR VGND sg13g2_decap_8
XFILLER_13_163 VPWR VGND sg13g2_fill_2
XFILLER_5_373 VPWR VGND sg13g2_decap_4
X_4130_ VPWR _3506_ net549 VGND sg13g2_inv_1
X_4061_ VPWR _3437_ net558 VGND sg13g2_inv_1
XFILLER_3_1026 VPWR VGND sg13g2_fill_2
X_7820_ net195 VGND VPWR _0298_ s0.data_out\[12\]\[5\] clknet_leaf_20_clk sg13g2_dfrbpq_2
XFILLER_36_233 VPWR VGND sg13g2_fill_1
XFILLER_25_907 VPWR VGND sg13g2_fill_2
XFILLER_18_981 VPWR VGND sg13g2_decap_8
XFILLER_25_929 VPWR VGND sg13g2_fill_2
X_7751_ net270 VGND VPWR net429 s0.was_valid_out\[17\][0] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_4963_ _0961_ net1488 _0960_ VPWR VGND sg13g2_nand2b_1
X_6702_ net1600 _2472_ _2529_ VPWR VGND sg13g2_nor2_1
X_7682_ net344 VGND VPWR _0160_ s0.shift_out\[23\][0] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_6633_ _2467_ net1291 net801 VPWR VGND sg13g2_nand2_1
X_4894_ VGND VPWR _0898_ _0900_ _0903_ net1682 sg13g2_a21oi_1
XFILLER_33_995 VPWR VGND sg13g2_decap_8
X_6564_ _0338_ _2405_ _2406_ _3505_ net1608 VPWR VGND sg13g2_a22oi_1
X_5515_ VGND VPWR net1426 _1463_ _1464_ _1461_ sg13g2_a21oi_1
X_6495_ VPWR VGND _2339_ net1711 _2337_ net1709 _2341_ _2333_ sg13g2_a221oi_1
X_5446_ net1744 VPWR _1398_ VGND _1395_ _1397_ sg13g2_o21ai_1
X_5377_ net1439 net1345 _1338_ VPWR VGND sg13g2_nor2b_1
X_4328_ _0385_ net1543 s0.data_out\[25\]\[2\] VPWR VGND sg13g2_nand2_1
X_7116_ net1242 net1347 _2902_ VPWR VGND sg13g2_nor2b_1
XFILLER_47_509 VPWR VGND sg13g2_fill_2
XFILLER_41_1010 VPWR VGND sg13g2_decap_8
X_4259_ _3621_ net1545 _3622_ _3623_ VPWR VGND sg13g2_a21o_1
X_7047_ net1261 VPWR _2844_ VGND _2786_ _2843_ sg13g2_o21ai_1
XFILLER_27_277 VPWR VGND sg13g2_fill_1
XFILLER_43_748 VPWR VGND sg13g2_fill_2
X_7949_ net55 VGND VPWR net569 s0.data_out\[2\]\[7\] clknet_leaf_8_clk sg13g2_dfrbpq_2
XFILLER_30_409 VPWR VGND sg13g2_fill_2
XFILLER_7_627 VPWR VGND sg13g2_fill_1
XFILLER_6_137 VPWR VGND sg13g2_fill_2
XFILLER_3_844 VPWR VGND sg13g2_decap_8
XFILLER_3_833 VPWR VGND sg13g2_decap_8
Xfanout1601 net1602 net1601 VPWR VGND sg13g2_buf_8
Xfanout1623 net1625 net1623 VPWR VGND sg13g2_buf_2
Xfanout1612 net1614 net1612 VPWR VGND sg13g2_buf_8
Xfanout1645 net1646 net1645 VPWR VGND sg13g2_buf_2
Xfanout1656 net1657 net1656 VPWR VGND sg13g2_buf_8
Xfanout1667 ui_in[6] net1667 VPWR VGND sg13g2_buf_8
Xfanout1634 net1636 net1634 VPWR VGND sg13g2_buf_8
Xfanout1678 net1681 net1678 VPWR VGND sg13g2_buf_1
Xfanout1689 ui_in[3] net1689 VPWR VGND sg13g2_buf_8
X_7965__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_37_70 VPWR VGND sg13g2_fill_1
XFILLER_19_789 VPWR VGND sg13g2_fill_2
XFILLER_18_1023 VPWR VGND sg13g2_decap_4
X_5300_ VGND VPWR net1450 net700 _1267_ _1229_ sg13g2_a21oi_1
X_6280_ _2157_ _2118_ _2156_ VPWR VGND sg13g2_nand2_1
X_5231_ _1204_ net487 net1467 VPWR VGND sg13g2_nand2b_1
X_5162_ _1145_ VPWR _1146_ VGND net1737 net691 sg13g2_o21ai_1
XFILLER_25_1016 VPWR VGND sg13g2_decap_8
X_4113_ VPWR _3489_ net597 VGND sg13g2_inv_1
X_5093_ net1458 net1354 _1078_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_1027 VPWR VGND sg13g2_fill_2
X_4044_ _3420_ net637 VPWR VGND sg13g2_inv_2
XFILLER_37_564 VPWR VGND sg13g2_fill_1
X_7803_ net213 VGND VPWR _0281_ s0.data_out\[13\]\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_2
XFILLER_24_203 VPWR VGND sg13g2_fill_2
X_5995_ _1896_ net418 net1398 VPWR VGND sg13g2_nand2b_1
X_7734_ net288 VGND VPWR net815 s0.data_out\[19\]\[3\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_4946_ net1468 _0940_ _0946_ VPWR VGND sg13g2_nor2_1
X_4877_ _0886_ net1489 net797 VPWR VGND sg13g2_nand2_1
X_7665_ net363 VGND VPWR _0143_ s0.data_out\[25\]\[6\] clknet_leaf_43_clk sg13g2_dfrbpq_2
X_7596_ net459 net1215 net1212 _3334_ VPWR VGND sg13g2_a21o_1
XFILLER_21_998 VPWR VGND sg13g2_decap_8
X_6616_ s0.data_out\[8\]\[0\] s0.data_out\[7\]\[0\] net1289 _2450_ VPWR VGND sg13g2_mux2_1
X_6547_ VGND VPWR _2377_ _2392_ _2393_ _2368_ sg13g2_a21oi_1
X_6478_ VGND VPWR _2205_ _2323_ _2324_ net1305 sg13g2_a21oi_1
XFILLER_0_803 VPWR VGND sg13g2_decap_8
X_5429_ net1451 VPWR _1383_ VGND _1320_ _1382_ sg13g2_o21ai_1
XFILLER_16_759 VPWR VGND sg13g2_decap_4
XFILLER_43_545 VPWR VGND sg13g2_fill_1
XFILLER_15_236 VPWR VGND sg13g2_fill_1
XFILLER_48_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_663 VPWR VGND sg13g2_fill_2
Xfanout1431 s0.shift_out\[16\][0] net1431 VPWR VGND sg13g2_buf_2
Xfanout1420 net1421 net1420 VPWR VGND sg13g2_buf_8
XFILLER_38_328 VPWR VGND sg13g2_fill_2
Xfanout1453 net1454 net1453 VPWR VGND sg13g2_buf_8
Xfanout1464 net1467 net1464 VPWR VGND sg13g2_buf_8
Xfanout1475 net1476 net1475 VPWR VGND sg13g2_buf_8
Xfanout1442 net460 net1442 VPWR VGND sg13g2_buf_2
Xfanout1497 s0.shift_out\[22\][0] net1497 VPWR VGND sg13g2_buf_2
Xfanout1486 net1488 net1486 VPWR VGND sg13g2_buf_8
XFILLER_46_394 VPWR VGND sg13g2_fill_1
XFILLER_34_534 VPWR VGND sg13g2_fill_1
X_4800_ VGND VPWR net1183 _0776_ _0815_ net1594 sg13g2_a21oi_1
XFILLER_15_770 VPWR VGND sg13g2_fill_2
X_5780_ _1622_ VPWR _1705_ VGND _1677_ _1680_ sg13g2_o21ai_1
X_4731_ _0751_ VPWR _0752_ VGND _0739_ _0749_ sg13g2_o21ai_1
X_4662_ net1182 _3435_ _0692_ VPWR VGND sg13g2_nor2_1
X_7450_ net1231 VPWR _3204_ VGND _3146_ _3203_ sg13g2_o21ai_1
XFILLER_31_1020 VPWR VGND sg13g2_decap_8
X_6401_ _2259_ net1320 _2258_ VPWR VGND sg13g2_nand2b_1
X_4593_ VGND VPWR net1525 _0623_ _0626_ _0625_ sg13g2_a21oi_1
X_7381_ VGND VPWR _3024_ _3142_ _3143_ net1230 sg13g2_a21oi_1
X_6332_ net1638 net1356 _2198_ VPWR VGND sg13g2_nor2_1
X_6263_ _2138_ net1325 _2139_ _2140_ VPWR VGND sg13g2_a21o_1
X_5214_ net1447 net1354 _1187_ VPWR VGND sg13g2_nor2b_1
X_6194_ net1379 VPWR _2075_ VGND _2015_ _2074_ sg13g2_o21ai_1
X_5145_ VGND VPWR _1002_ _1129_ _1130_ net1469 sg13g2_a21oi_1
X_5076_ net1460 _1058_ _1064_ VPWR VGND sg13g2_nor2_1
XFILLER_38_851 VPWR VGND sg13g2_fill_2
X_4027_ net1671 _3403_ VPWR VGND sg13g2_inv_4
XFILLER_37_394 VPWR VGND sg13g2_fill_1
XFILLER_25_545 VPWR VGND sg13g2_fill_2
X_5978_ _3418_ _1878_ _1879_ VPWR VGND sg13g2_and2_1
X_7717_ net306 VGND VPWR _0195_ s0.genblk1\[1\].modules.bubble clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
X_4929_ _0892_ _0931_ net1734 _0932_ VPWR VGND sg13g2_nand3_1
X_7648_ net37 VGND VPWR net622 s0.data_out\[26\]\[1\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_7579_ net1741 net394 _0098_ VPWR VGND sg13g2_and2_1
XFILLER_0_677 VPWR VGND sg13g2_decap_8
XFILLER_48_648 VPWR VGND sg13g2_decap_8
XFILLER_47_125 VPWR VGND sg13g2_fill_1
XFILLER_29_851 VPWR VGND sg13g2_fill_2
XFILLER_44_876 VPWR VGND sg13g2_decap_8
XFILLER_34_93 VPWR VGND sg13g2_decap_4
XFILLER_7_265 VPWR VGND sg13g2_fill_1
XFILLER_4_983 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_fill_2
Xfanout1250 net1251 net1250 VPWR VGND sg13g2_buf_2
XFILLER_22_1008 VPWR VGND sg13g2_decap_8
Xfanout1261 net1262 net1261 VPWR VGND sg13g2_buf_8
Xfanout1283 net1284 net1283 VPWR VGND sg13g2_buf_8
Xfanout1272 net1273 net1272 VPWR VGND sg13g2_buf_1
X_6950_ _2753_ VPWR _2754_ VGND net1729 net807 sg13g2_o21ai_1
Xfanout1294 net1300 net1294 VPWR VGND sg13g2_buf_8
X_5901_ _1811_ VPWR _1814_ VGND net1694 _1775_ sg13g2_o21ai_1
X_6881_ net1263 net1333 _2691_ VPWR VGND sg13g2_nor2b_1
X_5832_ net1749 net373 _0267_ VPWR VGND sg13g2_and2_1
XFILLER_14_19 VPWR VGND sg13g2_fill_2
XFILLER_22_559 VPWR VGND sg13g2_decap_4
X_5763_ _1688_ net1196 _1687_ VPWR VGND sg13g2_nand2_1
X_7502_ net1209 net1334 _3252_ VPWR VGND sg13g2_nor2b_1
X_4714_ VGND VPWR net1495 _0733_ _0735_ _0734_ sg13g2_a21oi_1
X_5694_ VGND VPWR net1196 _1509_ _1622_ _1621_ sg13g2_a21oi_1
X_7433_ net1587 _3135_ _3191_ VPWR VGND sg13g2_nor2_1
X_4645_ _0675_ _0676_ _0677_ _0678_ VPWR VGND sg13g2_nor3_1
XFILLER_30_29 VPWR VGND sg13g2_fill_2
X_4576_ net1725 VPWR _0612_ VGND net578 _0606_ sg13g2_o21ai_1
X_7364_ net1570 _3125_ _3126_ VPWR VGND sg13g2_and2_1
X_6315_ net1326 net522 _2184_ VPWR VGND sg13g2_and2_1
X_7295_ VGND VPWR net1228 net721 _3068_ _3001_ sg13g2_a21oi_1
X_6246_ _2123_ s0.data_out\[10\]\[6\] net1374 VPWR VGND sg13g2_nand2b_1
X_6177_ net1613 _2002_ _2062_ VPWR VGND sg13g2_nor2_1
X_5128_ VGND VPWR net1474 _1110_ _1113_ _1112_ sg13g2_a21oi_1
X_5059_ _0189_ _1049_ _1050_ _3442_ net1604 VPWR VGND sg13g2_a22oi_1
XFILLER_41_824 VPWR VGND sg13g2_fill_2
XFILLER_40_301 VPWR VGND sg13g2_fill_1
XFILLER_40_334 VPWR VGND sg13g2_fill_2
XFILLER_45_1019 VPWR VGND sg13g2_decap_8
XFILLER_49_913 VPWR VGND sg13g2_decap_8
XFILLER_1_964 VPWR VGND sg13g2_decap_8
XFILLER_0_474 VPWR VGND sg13g2_fill_2
Xhold82 _0289_ VPWR VGND net451 sg13g2_dlygate4sd3_1
Xhold60 _0229_ VPWR VGND net429 sg13g2_dlygate4sd3_1
Xhold71 s0.shift_out\[3\][0] VPWR VGND net440 sg13g2_dlygate4sd3_1
Xhold93 _0118_ VPWR VGND net462 sg13g2_dlygate4sd3_1
XFILLER_32_835 VPWR VGND sg13g2_decap_4
X_4430_ _0479_ net1714 _0480_ VPWR VGND _0422_ sg13g2_nand3b_1
X_4361_ s0.data_out\[26\]\[6\] s0.data_out\[25\]\[6\] net1540 _0418_ VPWR VGND sg13g2_mux2_1
X_7758__262 VPWR VGND net262 sg13g2_tiehi
X_6100_ s0.data_out\[12\]\[0\] s0.data_out\[11\]\[0\] net1373 _1989_ VPWR VGND sg13g2_mux2_1
X_4292_ net1561 VPWR _0358_ VGND _3566_ _0357_ sg13g2_o21ai_1
X_7080_ _2869_ net1633 net1247 VPWR VGND sg13g2_nand2_1
X_6031_ _1908_ VPWR _1932_ VGND _1899_ _1907_ sg13g2_o21ai_1
XFILLER_26_128 VPWR VGND sg13g2_fill_1
X_6933_ VGND VPWR net1261 s0.data_out\[5\]\[2\] _2740_ _2670_ sg13g2_a21oi_1
X_6864_ _2673_ VPWR _2674_ VGND net1175 _2671_ sg13g2_o21ai_1
XFILLER_25_29 VPWR VGND sg13g2_fill_2
X_5815_ _1732_ VPWR _1733_ VGND net1748 net772 sg13g2_o21ai_1
X_6795_ VGND VPWR _2617_ net1566 net383 sg13g2_or2_1
X_5746_ s0.data_out\[15\]\[6\] s0.data_out\[14\]\[6\] net1410 _1671_ VPWR VGND sg13g2_mux2_1
X_5677_ _0249_ _1607_ _1608_ _3468_ net1622 VPWR VGND sg13g2_a22oi_1
X_4628_ _0659_ _0660_ _0658_ _0661_ VPWR VGND sg13g2_nand3_1
X_7416_ VGND VPWR net1217 s0.data_out\[1\]\[0\] _3177_ _3121_ sg13g2_a21oi_1
X_7347_ s0.data_out\[1\]\[2\] s0.data_out\[2\]\[2\] net1237 _3109_ VPWR VGND sg13g2_mux2_1
X_4559_ net1538 VPWR _0597_ VGND _0539_ _0596_ sg13g2_o21ai_1
XFILLER_2_728 VPWR VGND sg13g2_decap_8
X_7278_ _3052_ net1237 net520 VPWR VGND sg13g2_nand2_1
X_6229_ s0.data_out\[10\]\[0\] s0.data_out\[11\]\[0\] net1372 _2106_ VPWR VGND sg13g2_mux2_1
XFILLER_17_117 VPWR VGND sg13g2_fill_1
XFILLER_13_334 VPWR VGND sg13g2_fill_2
XFILLER_5_544 VPWR VGND sg13g2_fill_2
Xoutput4 net4 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_761 VPWR VGND sg13g2_decap_8
XFILLER_49_710 VPWR VGND sg13g2_decap_8
XFILLER_49_787 VPWR VGND sg13g2_decap_8
XFILLER_36_459 VPWR VGND sg13g2_fill_2
X_6580_ net1310 VPWR _2419_ VGND _2360_ _2418_ sg13g2_o21ai_1
X_5600_ _1537_ net1424 _1536_ VPWR VGND sg13g2_nand2b_1
X_5531_ VGND VPWR net1423 s0.data_out\[16\]\[0\] _1479_ _1408_ sg13g2_a21oi_1
XFILLER_8_382 VPWR VGND sg13g2_fill_1
X_5462_ _1411_ net1437 _1410_ VPWR VGND sg13g2_nand2b_1
X_7201_ _0058_ _2978_ _2979_ _3532_ net1580 VPWR VGND sg13g2_a22oi_1
X_5393_ _1350_ VPWR _1354_ VGND net1684 _1342_ sg13g2_o21ai_1
X_4413_ net1551 VPWR _0467_ VGND _0387_ _0466_ sg13g2_o21ai_1
X_4344_ net1535 net1356 _0401_ VPWR VGND sg13g2_nor2b_1
X_7132_ _2916_ _2917_ _2918_ VPWR VGND sg13g2_nor2_1
X_7063_ net454 s0.data_out\[4\]\[4\] _2856_ VPWR VGND sg13g2_and2_1
X_6014_ _1915_ net723 net1398 VPWR VGND sg13g2_nand2b_1
X_4275_ _3638_ VPWR _0344_ VGND _3587_ _3596_ sg13g2_o21ai_1
XFILLER_27_415 VPWR VGND sg13g2_fill_1
X_7965_ net158 VGND VPWR _0099_ s0.shift_out\[0\][0] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_6916_ _2713_ _2711_ net1670 _2726_ VPWR VGND sg13g2_a21o_1
XFILLER_36_993 VPWR VGND sg13g2_decap_8
X_7896_ net113 VGND VPWR _0030_ s0.data_out\[6\]\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_6847_ _2655_ net1261 _2656_ _2657_ VPWR VGND sg13g2_a21o_1
XFILLER_35_1018 VPWR VGND sg13g2_decap_8
X_6778_ VGND VPWR _2600_ _2599_ _3406_ sg13g2_or2_1
X_5729_ net1403 net1168 _1654_ VPWR VGND sg13g2_nor2_1
Xhold360 s0.shift_out\[13\][0] VPWR VGND net729 sg13g2_dlygate4sd3_1
Xhold371 s0.data_out\[23\]\[0\] VPWR VGND net740 sg13g2_dlygate4sd3_1
Xhold393 s0.data_out\[25\]\[2\] VPWR VGND net762 sg13g2_dlygate4sd3_1
Xhold382 _3184_ VPWR VGND net751 sg13g2_dlygate4sd3_1
XFILLER_46_702 VPWR VGND sg13g2_decap_8
XFILLER_46_779 VPWR VGND sg13g2_decap_8
XFILLER_27_971 VPWR VGND sg13g2_decap_8
XFILLER_42_996 VPWR VGND sg13g2_decap_8
X_7755__265 VPWR VGND net265 sg13g2_tiehi
XFILLER_3_87 VPWR VGND sg13g2_fill_1
X_4060_ VPWR _3436_ net816 VGND sg13g2_inv_1
XFILLER_49_584 VPWR VGND sg13g2_decap_8
XFILLER_36_201 VPWR VGND sg13g2_fill_2
XFILLER_3_1005 VPWR VGND sg13g2_decap_8
XFILLER_45_790 VPWR VGND sg13g2_fill_1
X_7750_ net271 VGND VPWR _0228_ s0.data_out\[18\]\[7\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_4962_ VGND VPWR net1470 _0959_ _0960_ _0957_ sg13g2_a21oi_1
XFILLER_17_481 VPWR VGND sg13g2_fill_2
X_6701_ net1297 VPWR _2528_ VGND _2469_ _2527_ sg13g2_o21ai_1
X_7681_ net345 VGND VPWR _0159_ s0.genblk1\[22\].modules.bubble clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_4893_ _0902_ _0893_ _0901_ VPWR VGND sg13g2_nand2_1
XFILLER_33_974 VPWR VGND sg13g2_decap_8
X_7762__258 VPWR VGND net258 sg13g2_tiehi
X_6632_ VPWR VGND net1691 _2458_ _2465_ net1699 _2466_ _2441_ sg13g2_a221oi_1
XFILLER_20_668 VPWR VGND sg13g2_fill_1
X_6563_ net1608 _2324_ _2406_ VPWR VGND sg13g2_nor2_1
X_5514_ s0.data_out\[17\]\[4\] s0.data_out\[16\]\[4\] net1433 _1463_ VPWR VGND sg13g2_mux2_1
X_6494_ net1705 _2333_ _2340_ VPWR VGND sg13g2_nor2_1
X_5445_ _1397_ _1394_ _1396_ VPWR VGND sg13g2_nand2_1
X_5376_ _1336_ VPWR _1337_ VGND net1445 _3459_ sg13g2_o21ai_1
X_7115_ s0.data_out\[4\]\[3\] s0.data_out\[3\]\[3\] net1245 _2901_ VPWR VGND sg13g2_mux2_1
X_4327_ net1716 net379 _0123_ VPWR VGND sg13g2_and2_1
XFILLER_47_16 VPWR VGND sg13g2_fill_2
X_4258_ net1545 net1338 _3622_ VPWR VGND sg13g2_nor2b_1
X_7046_ net1251 s0.data_out\[4\]\[0\] _2843_ VPWR VGND sg13g2_and2_1
X_4189_ VGND VPWR _3556_ _3555_ _3554_ sg13g2_or2_1
X_7948_ net57 VGND VPWR _0082_ s0.data_out\[2\]\[6\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_7879_ net131 VGND VPWR _0013_ s0.valid_out\[7\][0] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_11_613 VPWR VGND sg13g2_fill_2
XFILLER_23_495 VPWR VGND sg13g2_fill_1
XFILLER_6_105 VPWR VGND sg13g2_fill_1
XFILLER_3_812 VPWR VGND sg13g2_decap_8
XFILLER_12_85 VPWR VGND sg13g2_fill_2
Xfanout1624 net1625 net1624 VPWR VGND sg13g2_buf_8
Xhold190 s0.data_out\[27\]\[1\] VPWR VGND net559 sg13g2_dlygate4sd3_1
Xfanout1602 net1603 net1602 VPWR VGND sg13g2_buf_8
Xfanout1613 net1614 net1613 VPWR VGND sg13g2_buf_1
Xfanout1646 uio_in[0] net1646 VPWR VGND sg13g2_buf_8
Xfanout1657 ui_in[7] net1657 VPWR VGND sg13g2_buf_8
Xfanout1635 net1636 net1635 VPWR VGND sg13g2_buf_8
Xfanout1668 net1672 net1668 VPWR VGND sg13g2_buf_8
Xfanout1679 net1681 net1679 VPWR VGND sg13g2_buf_8
XFILLER_46_532 VPWR VGND sg13g2_fill_1
XFILLER_18_1002 VPWR VGND sg13g2_decap_8
XFILLER_15_996 VPWR VGND sg13g2_decap_8
X_5230_ _1201_ net1452 _1202_ _1203_ VPWR VGND sg13g2_a21o_1
X_5161_ _1088_ _1144_ net1736 _1145_ VPWR VGND sg13g2_nand3_1
X_4112_ VPWR _3488_ net746 VGND sg13g2_inv_1
X_5092_ _1076_ VPWR _1077_ VGND net1465 _3450_ sg13g2_o21ai_1
X_4043_ VPWR _3419_ net572 VGND sg13g2_inv_1
XFILLER_37_532 VPWR VGND sg13g2_fill_2
X_7802_ net214 VGND VPWR _0280_ s0.shift_out\[13\][0] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5994_ _1893_ net1382 _1894_ _1895_ VPWR VGND sg13g2_a21o_1
XFILLER_25_738 VPWR VGND sg13g2_fill_2
X_4945_ _0942_ VPWR _0945_ VGND s0.was_valid_out\[20\][0] net1478 sg13g2_o21ai_1
X_7733_ net289 VGND VPWR net635 s0.data_out\[19\]\[2\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_4876_ _0882_ _0883_ _0884_ _0885_ VPWR VGND sg13g2_nor3_1
X_7664_ net364 VGND VPWR _0142_ s0.data_out\[25\]\[5\] clknet_leaf_43_clk sg13g2_dfrbpq_2
X_7595_ net1702 _3329_ _3333_ VPWR VGND sg13g2_nor2_1
XFILLER_21_977 VPWR VGND sg13g2_decap_8
X_6615_ VGND VPWR net1293 _2446_ _2449_ _2448_ sg13g2_a21oi_1
X_6546_ _2376_ _3403_ _2385_ _2392_ VPWR VGND sg13g2_a21o_1
X_6477_ _2323_ s0.data_out\[8\]\[2\] net1314 VPWR VGND sg13g2_nand2b_1
X_5428_ net1441 s0.data_out\[17\]\[6\] _1382_ VPWR VGND sg13g2_and2_1
X_5359_ net1441 net1336 _1320_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_859 VPWR VGND sg13g2_decap_8
X_7029_ s0.data_out\[5\]\[5\] s0.data_out\[4\]\[5\] net1256 _2827_ VPWR VGND sg13g2_mux2_1
XFILLER_15_259 VPWR VGND sg13g2_decap_4
XFILLER_7_469 VPWR VGND sg13g2_fill_1
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
Xfanout1410 s0.valid_out\[14\][0] net1410 VPWR VGND sg13g2_buf_8
Xfanout1432 net1435 net1432 VPWR VGND sg13g2_buf_8
Xfanout1421 net1422 net1421 VPWR VGND sg13g2_buf_8
X_7752__268 VPWR VGND net268 sg13g2_tiehi
Xfanout1454 net1456 net1454 VPWR VGND sg13g2_buf_8
Xfanout1465 net1467 net1465 VPWR VGND sg13g2_buf_8
Xfanout1443 net1446 net1443 VPWR VGND sg13g2_buf_8
XFILLER_24_8 VPWR VGND sg13g2_decap_4
Xfanout1498 net1499 net1498 VPWR VGND sg13g2_buf_8
Xfanout1476 net1477 net1476 VPWR VGND sg13g2_buf_2
Xfanout1487 net1488 net1487 VPWR VGND sg13g2_buf_1
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_47_885 VPWR VGND sg13g2_decap_8
XFILLER_0_55 VPWR VGND sg13g2_fill_1
XFILLER_9_53 VPWR VGND sg13g2_fill_2
X_4730_ _0751_ net1690 _0748_ VPWR VGND sg13g2_nand2_1
X_4661_ _0150_ _0690_ _0691_ _3431_ net1590 VPWR VGND sg13g2_a22oi_1
XFILLER_30_752 VPWR VGND sg13g2_fill_1
X_7380_ _3142_ s0.data_out\[1\]\[6\] net1236 VPWR VGND sg13g2_nand2b_1
X_6400_ VGND VPWR net1312 _2256_ _2258_ _2257_ sg13g2_a21oi_1
X_6331_ net1610 _2195_ _0314_ VPWR VGND sg13g2_nor2_1
X_4592_ VGND VPWR _0494_ _0624_ _0625_ net1525 sg13g2_a21oi_1
X_6262_ net1325 net1346 _2139_ VPWR VGND sg13g2_nor2b_1
X_6193_ _3383_ _3495_ _2074_ VPWR VGND sg13g2_nor2_1
X_5213_ _1185_ VPWR _1186_ VGND net1453 _3456_ sg13g2_o21ai_1
X_5144_ _1129_ s0.data_out\[19\]\[5\] net1480 VPWR VGND sg13g2_nand2b_1
XFILLER_29_318 VPWR VGND sg13g2_fill_1
X_5075_ VGND VPWR _1063_ _1062_ _1060_ sg13g2_or2_1
XFILLER_29_329 VPWR VGND sg13g2_fill_1
X_4026_ _3402_ net1658 VPWR VGND sg13g2_inv_2
X_5977_ _1877_ VPWR _1878_ VGND net1192 _1875_ sg13g2_o21ai_1
X_4928_ net1499 VPWR _0931_ VGND _0888_ _0930_ sg13g2_o21ai_1
X_7716_ net307 VGND VPWR _0194_ s0.valid_out\[20\][0] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_7647_ net38 VGND VPWR _0125_ s0.data_out\[26\]\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_2
XFILLER_20_240 VPWR VGND sg13g2_fill_2
X_4859_ s0.data_out\[22\]\[7\] s0.data_out\[21\]\[7\] net1490 _0868_ VPWR VGND sg13g2_mux2_1
X_7578_ net1639 _3317_ _0097_ VPWR VGND sg13g2_nor2_1
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
X_6529_ _2375_ _2374_ VPWR VGND net1309 sg13g2_nand2b_2
XFILLER_0_645 VPWR VGND sg13g2_decap_8
XFILLER_44_855 VPWR VGND sg13g2_decap_8
XFILLER_4_962 VPWR VGND sg13g2_decap_8
Xfanout1240 net1241 net1240 VPWR VGND sg13g2_buf_8
Xfanout1251 net1252 net1251 VPWR VGND sg13g2_buf_8
Xfanout1262 net480 net1262 VPWR VGND sg13g2_buf_8
Xfanout1273 net445 net1273 VPWR VGND sg13g2_buf_1
Xfanout1284 s0.shift_out\[7\][0] net1284 VPWR VGND sg13g2_buf_8
Xfanout1295 net1300 net1295 VPWR VGND sg13g2_buf_2
XFILLER_47_682 VPWR VGND sg13g2_decap_8
X_5900_ _1813_ _3406_ _1803_ VPWR VGND sg13g2_xnor2_1
X_6880_ s0.data_out\[6\]\[6\] s0.data_out\[5\]\[6\] net1268 _2690_ VPWR VGND sg13g2_mux2_1
X_5831_ net1629 _1740_ _0266_ VPWR VGND sg13g2_nor2_1
X_5762_ _1575_ VPWR _1687_ VGND net1420 _3477_ sg13g2_o21ai_1
X_7501_ s0.data_out\[1\]\[6\] s0.data_out\[0\]\[6\] net1214 _3251_ VPWR VGND sg13g2_mux2_1
X_4713_ net1495 net1349 _0734_ VPWR VGND sg13g2_nor2b_1
X_5693_ _1619_ _1620_ _1621_ VPWR VGND sg13g2_nor2_1
X_7432_ net1233 VPWR _3190_ VGND _3132_ _3189_ sg13g2_o21ai_1
X_4644_ net1679 _0667_ _0677_ VPWR VGND sg13g2_nor2_1
X_4575_ _0609_ _0610_ _0611_ VPWR VGND sg13g2_nor2_1
X_7363_ _3124_ VPWR _3125_ VGND net1187 _3122_ sg13g2_o21ai_1
X_6314_ VPWR _0311_ net688 VGND sg13g2_inv_1
X_7294_ VGND VPWR _3063_ _3066_ _0063_ _3067_ sg13g2_a21oi_1
X_6245_ _2120_ net1325 _2121_ _2122_ VPWR VGND sg13g2_a21o_1
X_6176_ net1377 VPWR _2061_ VGND _1999_ _2060_ sg13g2_o21ai_1
X_5127_ VGND VPWR _0984_ _1111_ _1112_ net1474 sg13g2_a21oi_1
XFILLER_29_104 VPWR VGND sg13g2_fill_2
X_5058_ net1604 _1007_ _1050_ VPWR VGND sg13g2_nor2_1
X_4009_ VPWR _3385_ s0.valid_out\[27\][0] VGND sg13g2_inv_1
XFILLER_25_332 VPWR VGND sg13g2_fill_2
X_7807__209 VPWR VGND net209 sg13g2_tiehi
XFILLER_40_313 VPWR VGND sg13g2_fill_1
XFILLER_4_247 VPWR VGND sg13g2_fill_1
XFILLER_1_943 VPWR VGND sg13g2_decap_8
Xhold50 s0.was_valid_out\[25\][0] VPWR VGND net419 sg13g2_dlygate4sd3_1
XFILLER_49_969 VPWR VGND sg13g2_decap_8
Xhold72 s0.was_valid_out\[10\][0] VPWR VGND net441 sg13g2_dlygate4sd3_1
Xhold61 s0.data_out\[0\]\[1\] VPWR VGND net430 sg13g2_dlygate4sd3_1
Xhold83 s0.data_out\[26\]\[3\] VPWR VGND net452 sg13g2_dlygate4sd3_1
Xhold94 s0.was_valid_out\[11\][0] VPWR VGND net463 sg13g2_dlygate4sd3_1
XFILLER_44_652 VPWR VGND sg13g2_fill_2
XFILLER_32_858 VPWR VGND sg13g2_decap_4
X_7897__112 VPWR VGND net112 sg13g2_tiehi
X_4360_ _0417_ net1542 net775 VPWR VGND sg13g2_nand2_1
X_4291_ net1546 net464 _0357_ VPWR VGND sg13g2_and2_1
X_6030_ _1907_ _1909_ _1910_ _1930_ _1931_ VPWR VGND sg13g2_nor4_1
XFILLER_20_2 VPWR VGND sg13g2_fill_1
XFILLER_48_991 VPWR VGND sg13g2_decap_8
XFILLER_26_107 VPWR VGND sg13g2_fill_1
X_6932_ _0029_ _2738_ _2739_ _3523_ net1590 VPWR VGND sg13g2_a22oi_1
X_6863_ _2673_ net1175 _2672_ VPWR VGND sg13g2_nand2_1
XFILLER_35_663 VPWR VGND sg13g2_fill_1
XFILLER_23_836 VPWR VGND sg13g2_fill_2
X_5814_ _1731_ net1748 _1732_ VPWR VGND _1675_ sg13g2_nand3b_1
XFILLER_34_162 VPWR VGND sg13g2_fill_1
X_6794_ VPWR VGND _2592_ _2536_ _2614_ _2574_ _2616_ _2613_ sg13g2_a221oi_1
X_5745_ _1670_ net1411 net696 VPWR VGND sg13g2_nand2_1
XFILLER_10_519 VPWR VGND sg13g2_decap_8
X_5676_ net1622 _1573_ _1608_ VPWR VGND sg13g2_nor2_1
X_7415_ net371 net1565 _3176_ _0075_ VPWR VGND sg13g2_nor3_1
X_4627_ VGND VPWR _0660_ _0650_ net1650 sg13g2_or2_1
X_7346_ VGND VPWR net1222 _3106_ _3108_ _3107_ sg13g2_a21oi_1
X_4558_ net1519 s0.data_out\[24\]\[6\] _0596_ VPWR VGND sg13g2_and2_1
X_4489_ _0534_ net525 net1542 VPWR VGND sg13g2_nand2b_1
X_7277_ _3039_ _3050_ _3051_ VPWR VGND sg13g2_and2_1
X_7813__202 VPWR VGND net202 sg13g2_tiehi
X_6228_ _2105_ net1365 _2104_ VPWR VGND sg13g2_nand2b_1
X_6159_ _1967_ _2046_ _2047_ _2048_ VPWR VGND sg13g2_nor3_1
XFILLER_46_939 VPWR VGND sg13g2_decap_8
XFILLER_45_438 VPWR VGND sg13g2_fill_1
XFILLER_38_490 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_37_clk clknet_3_4__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_41_600 VPWR VGND sg13g2_fill_1
XFILLER_15_85 VPWR VGND sg13g2_fill_2
Xoutput5 net5 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_740 VPWR VGND sg13g2_decap_8
XFILLER_49_766 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_28_clk clknet_3_6__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_32_666 VPWR VGND sg13g2_fill_1
XFILLER_13_891 VPWR VGND sg13g2_fill_2
X_5530_ VGND VPWR _1474_ _1477_ _0232_ _1478_ sg13g2_a21oi_1
X_5461_ VGND VPWR net1423 _1409_ _1410_ _1408_ sg13g2_a21oi_1
X_4412_ net1186 _3423_ _0466_ VPWR VGND sg13g2_nor2_1
X_7200_ net1580 _2941_ _2979_ VPWR VGND sg13g2_nor2_1
X_5392_ _1351_ _1352_ _1353_ VPWR VGND sg13g2_nor2_1
X_4343_ s0.data_out\[26\]\[0\] s0.data_out\[25\]\[0\] net1541 _0400_ VPWR VGND sg13g2_mux2_1
X_7131_ net1686 _2906_ _2917_ VPWR VGND sg13g2_nor2_1
X_4274_ _3616_ _3634_ _3636_ _3637_ _3638_ VPWR VGND sg13g2_nor4_1
X_7062_ _0043_ _2854_ _2855_ _3528_ net1596 VPWR VGND sg13g2_a22oi_1
X_6013_ _1912_ net1382 _1913_ _1914_ VPWR VGND sg13g2_a21o_1
X_7964_ net178 VGND VPWR _0098_ s0.genblk1\[9\].modules.bubble clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_19_clk clknet_3_6__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
X_6915_ VGND VPWR _2711_ _2713_ _2725_ net1670 sg13g2_a21oi_1
XFILLER_36_972 VPWR VGND sg13g2_decap_8
X_7895_ net114 VGND VPWR net695 s0.data_out\[6\]\[1\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_35_482 VPWR VGND sg13g2_fill_2
X_6846_ net1261 net1353 _2656_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_666 VPWR VGND sg13g2_decap_4
X_6777_ _2598_ VPWR _2599_ VGND net1176 _2596_ sg13g2_o21ai_1
XFILLER_22_176 VPWR VGND sg13g2_decap_8
X_3989_ VPWR _3365_ net405 VGND sg13g2_inv_1
X_5728_ _1652_ VPWR _1653_ VGND net1409 _3473_ sg13g2_o21ai_1
XFILLER_6_309 VPWR VGND sg13g2_fill_1
X_5659_ _1539_ _1594_ net1742 _1595_ VPWR VGND sg13g2_nand3_1
Xhold350 s0.data_out\[6\]\[6\] VPWR VGND net719 sg13g2_dlygate4sd3_1
X_7329_ net1582 _3037_ _3095_ VPWR VGND sg13g2_nor2_1
Xhold361 s0.data_out\[14\]\[2\] VPWR VGND net730 sg13g2_dlygate4sd3_1
Xhold394 _0584_ VPWR VGND net763 sg13g2_dlygate4sd3_1
Xhold372 _0799_ VPWR VGND net741 sg13g2_dlygate4sd3_1
Xhold383 s0.data_out\[5\]\[1\] VPWR VGND net752 sg13g2_dlygate4sd3_1
XFILLER_19_917 VPWR VGND sg13g2_fill_2
XFILLER_46_758 VPWR VGND sg13g2_decap_8
X_7748__273 VPWR VGND net273 sg13g2_tiehi
XFILLER_42_975 VPWR VGND sg13g2_decap_8
X_7894__115 VPWR VGND net115 sg13g2_tiehi
XFILLER_3_22 VPWR VGND sg13g2_fill_2
XFILLER_3_33 VPWR VGND sg13g2_fill_1
XFILLER_49_563 VPWR VGND sg13g2_decap_8
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
XFILLER_36_279 VPWR VGND sg13g2_fill_2
X_4961_ s0.data_out\[21\]\[1\] s0.data_out\[20\]\[1\] net1478 _0959_ VPWR VGND sg13g2_mux2_1
X_6700_ net1287 s0.data_out\[7\]\[6\] _2527_ VPWR VGND sg13g2_and2_1
X_7680_ net346 VGND VPWR _0158_ s0.valid_out\[23\][0] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_4892_ _0898_ _0900_ net1682 _0901_ VPWR VGND sg13g2_nand3_1
XFILLER_32_474 VPWR VGND sg13g2_fill_1
X_6631_ VGND VPWR net1294 _2462_ _2465_ _2464_ sg13g2_a21oi_1
X_6562_ net1305 VPWR _2405_ VGND _2321_ _2404_ sg13g2_o21ai_1
X_5513_ _1462_ net1433 net791 VPWR VGND sg13g2_nand2_1
X_6493_ _2339_ _2338_ net1307 VPWR VGND sg13g2_nand2b_1
X_5444_ net1207 VPWR _1396_ VGND s0.was_valid_out\[16\][0] net1444 sg13g2_o21ai_1
Xclkbuf_leaf_8_clk clknet_3_2__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_5375_ _1336_ net1445 s0.data_out\[17\]\[4\] VPWR VGND sg13g2_nand2_1
X_7114_ _2900_ net1245 net794 VPWR VGND sg13g2_nand2_1
X_4326_ net1577 _0377_ _0378_ _0122_ VPWR VGND sg13g2_nor3_1
X_4257_ s0.data_out\[27\]\[5\] s0.data_out\[26\]\[5\] net1554 _3621_ VPWR VGND sg13g2_mux2_1
X_7045_ VGND VPWR _2838_ _2841_ _0039_ _2842_ sg13g2_a21oi_1
X_4188_ VGND VPWR net1633 net1563 _3555_ net1559 sg13g2_a21oi_1
X_7947_ net58 VGND VPWR _0081_ s0.data_out\[2\]\[5\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_7878_ net133 VGND VPWR _0012_ s0.was_valid_out\[7\][0] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6829_ _3396_ _3519_ _2643_ VPWR VGND sg13g2_nor2_1
XFILLER_24_986 VPWR VGND sg13g2_decap_8
XFILLER_10_135 VPWR VGND sg13g2_fill_2
XFILLER_12_97 VPWR VGND sg13g2_fill_2
XFILLER_3_879 VPWR VGND sg13g2_decap_8
Xhold180 s0.data_out\[9\]\[1\] VPWR VGND net549 sg13g2_dlygate4sd3_1
Xhold191 _0114_ VPWR VGND net560 sg13g2_dlygate4sd3_1
Xfanout1603 net1632 net1603 VPWR VGND sg13g2_buf_8
Xfanout1614 net1615 net1614 VPWR VGND sg13g2_buf_8
Xfanout1658 net1662 net1658 VPWR VGND sg13g2_buf_8
Xfanout1636 _3373_ net1636 VPWR VGND sg13g2_buf_8
Xfanout1647 net1652 net1647 VPWR VGND sg13g2_buf_8
Xfanout1625 net1632 net1625 VPWR VGND sg13g2_buf_8
Xfanout1669 net1672 net1669 VPWR VGND sg13g2_buf_1
XFILLER_33_249 VPWR VGND sg13g2_fill_2
XFILLER_15_975 VPWR VGND sg13g2_decap_8
XFILLER_10_680 VPWR VGND sg13g2_fill_1
XFILLER_6_640 VPWR VGND sg13g2_fill_2
X_5160_ net1475 VPWR _1144_ VGND _1084_ _1143_ sg13g2_o21ai_1
X_4111_ VPWR _3487_ net540 VGND sg13g2_inv_1
X_5091_ _1076_ net1465 net709 VPWR VGND sg13g2_nand2_1
X_4042_ VPWR _3418_ net1710 VGND sg13g2_inv_1
X_5993_ net1382 net1346 _1894_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_205 VPWR VGND sg13g2_fill_1
XFILLER_25_728 VPWR VGND sg13g2_fill_1
X_7801_ net215 VGND VPWR _0279_ s0.genblk1\[12\].modules.bubble clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_4944_ _0942_ _0943_ _0944_ VPWR VGND sg13g2_nor2_1
X_7732_ net290 VGND VPWR net710 s0.data_out\[19\]\[1\] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_21_901 VPWR VGND sg13g2_fill_1
X_4875_ net1653 _0873_ _0884_ VPWR VGND sg13g2_nor2_1
X_7663_ net365 VGND VPWR _0141_ s0.data_out\[25\]\[4\] clknet_leaf_42_clk sg13g2_dfrbpq_2
XFILLER_32_282 VPWR VGND sg13g2_fill_2
X_7594_ VPWR VGND _3331_ net1710 _3330_ net1702 _3332_ _3329_ sg13g2_a221oi_1
XFILLER_20_455 VPWR VGND sg13g2_fill_2
X_6614_ VGND VPWR _2327_ _2447_ _2448_ net1293 sg13g2_a21oi_1
X_6545_ _2350_ _2368_ _2386_ _2390_ _2391_ VPWR VGND sg13g2_or4_1
X_6476_ _2320_ net1295 _2321_ _2322_ VPWR VGND sg13g2_a21o_1
X_5427_ _0226_ _1380_ _1381_ _3458_ net1624 VPWR VGND sg13g2_a22oi_1
X_5358_ s0.data_out\[18\]\[6\] s0.data_out\[17\]\[6\] net1444 _1319_ VPWR VGND sg13g2_mux2_1
XFILLER_0_838 VPWR VGND sg13g2_decap_8
XFILLER_48_809 VPWR VGND sg13g2_decap_8
X_4309_ net1575 _3607_ _0371_ VPWR VGND sg13g2_nor2_1
X_5289_ net1463 VPWR _1259_ VGND _1179_ _1258_ sg13g2_o21ai_1
X_7028_ _2826_ net1254 s0.data_out\[4\]\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_43_536 VPWR VGND sg13g2_fill_2
X_7745__276 VPWR VGND net276 sg13g2_tiehi
XFILLER_12_989 VPWR VGND sg13g2_decap_8
XFILLER_8_949 VPWR VGND sg13g2_fill_1
X_7891__118 VPWR VGND net118 sg13g2_tiehi
XFILLER_3_621 VPWR VGND sg13g2_fill_2
Xfanout1400 net831 net1400 VPWR VGND sg13g2_buf_8
Xfanout1411 s0.valid_out\[14\][0] net1411 VPWR VGND sg13g2_buf_1
Xfanout1422 s0.valid_out\[15\][0] net1422 VPWR VGND sg13g2_buf_8
Xfanout1455 net1456 net1455 VPWR VGND sg13g2_buf_8
Xfanout1466 net1467 net1466 VPWR VGND sg13g2_buf_2
Xfanout1444 net1445 net1444 VPWR VGND sg13g2_buf_8
Xfanout1433 net1435 net1433 VPWR VGND sg13g2_buf_8
Xfanout1499 net424 net1499 VPWR VGND sg13g2_buf_2
Xfanout1477 s0.shift_out\[20\][0] net1477 VPWR VGND sg13g2_buf_1
Xfanout1488 net477 net1488 VPWR VGND sg13g2_buf_8
XFILLER_47_864 VPWR VGND sg13g2_decap_8
XFILLER_0_45 VPWR VGND sg13g2_fill_1
XFILLER_19_577 VPWR VGND sg13g2_decap_4
XFILLER_21_208 VPWR VGND sg13g2_fill_2
XFILLER_42_591 VPWR VGND sg13g2_fill_1
X_4660_ net1590 _0625_ _0691_ VPWR VGND sg13g2_nor2_1
X_6330_ _2196_ _2197_ _0313_ VPWR VGND sg13g2_nor2_1
X_4591_ _0624_ s0.data_out\[23\]\[1\] net1531 VPWR VGND sg13g2_nand2b_1
X_6261_ s0.data_out\[11\]\[4\] s0.data_out\[10\]\[4\] net1363 _2138_ VPWR VGND sg13g2_mux2_1
X_6192_ VPWR _0299_ net724 VGND sg13g2_inv_1
X_5212_ _1185_ net1453 s0.data_out\[18\]\[1\] VPWR VGND sg13g2_nand2_1
X_5143_ _1126_ net1457 _1127_ _1128_ VPWR VGND sg13g2_a21o_1
XFILLER_9_1023 VPWR VGND sg13g2_decap_4
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_5074_ net437 net1464 _1062_ VPWR VGND sg13g2_nor2_1
X_4025_ VPWR _3401_ net1333 VGND sg13g2_inv_1
XFILLER_38_864 VPWR VGND sg13g2_fill_2
XFILLER_38_853 VPWR VGND sg13g2_fill_1
XFILLER_25_547 VPWR VGND sg13g2_fill_1
X_5976_ _1877_ net1192 _1876_ VPWR VGND sg13g2_nand2_1
XFILLER_40_528 VPWR VGND sg13g2_fill_2
X_7715_ net309 VGND VPWR net652 s0.was_valid_out\[20\][0] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_4927_ net1180 _3442_ _0930_ VPWR VGND sg13g2_nor2_1
X_7646_ net39 VGND VPWR _0124_ s0.shift_out\[26\][0] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_4858_ _0867_ net1489 net538 VPWR VGND sg13g2_nand2_1
X_7699__326 VPWR VGND net326 sg13g2_tiehi
X_7577_ _3316_ _3317_ _0096_ VPWR VGND sg13g2_nor2_1
X_4789_ VPWR _0163_ net620 VGND sg13g2_inv_1
X_6528_ _2263_ VPWR _2374_ VGND net1316 _3509_ sg13g2_o21ai_1
X_6459_ net1310 VPWR _2308_ VGND net1646 net1298 sg13g2_o21ai_1
XFILLER_0_624 VPWR VGND sg13g2_decap_8
XFILLER_48_606 VPWR VGND sg13g2_decap_8
XFILLER_34_62 VPWR VGND sg13g2_decap_8
XFILLER_15_1017 VPWR VGND sg13g2_decap_8
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
XFILLER_4_941 VPWR VGND sg13g2_decap_8
Xfanout1241 net1244 net1241 VPWR VGND sg13g2_buf_8
Xfanout1230 net1231 net1230 VPWR VGND sg13g2_buf_8
Xfanout1274 net1275 net1274 VPWR VGND sg13g2_buf_8
Xfanout1263 net1265 net1263 VPWR VGND sg13g2_buf_8
Xfanout1252 net454 net1252 VPWR VGND sg13g2_buf_8
Xfanout1285 net1288 net1285 VPWR VGND sg13g2_buf_8
Xfanout1296 net1299 net1296 VPWR VGND sg13g2_buf_8
XFILLER_47_661 VPWR VGND sg13g2_decap_8
XFILLER_35_845 VPWR VGND sg13g2_fill_1
X_5830_ VGND VPWR _1741_ _1744_ _0265_ _1745_ sg13g2_a21oi_1
X_5761_ _1686_ net1417 _1685_ VPWR VGND sg13g2_nand2b_1
X_7500_ s0.data_out\[0\]\[6\] s0.data_out\[1\]\[6\] net1225 _3250_ VPWR VGND sg13g2_mux2_1
X_4712_ _0732_ VPWR _0733_ VGND net1504 _3435_ sg13g2_o21ai_1
X_7431_ net1221 net614 _3189_ VPWR VGND sg13g2_and2_1
X_5692_ net1645 net1410 _1620_ VPWR VGND sg13g2_nor2b_1
X_4643_ net1671 _0673_ _0676_ VPWR VGND sg13g2_nor2_1
X_4574_ VGND VPWR _3370_ _3389_ _0610_ net1523 sg13g2_a21oi_1
X_7362_ _3124_ net1187 _3123_ VPWR VGND sg13g2_nand2_1
X_6313_ _2182_ VPWR _2183_ VGND net1739 net687 sg13g2_o21ai_1
X_7293_ VGND VPWR _3067_ net1565 net381 sg13g2_or2_1
X_6244_ net1326 net1335 _2121_ VPWR VGND sg13g2_nor2b_1
X_6175_ _3383_ _3493_ _2060_ VPWR VGND sg13g2_nor2_1
X_5126_ _1111_ s0.data_out\[19\]\[7\] net1480 VPWR VGND sg13g2_nand2b_1
X_5057_ net1484 VPWR _1049_ VGND _1004_ _1048_ sg13g2_o21ai_1
X_4008_ VPWR _3384_ net1239 VGND sg13g2_inv_1
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
X_5959_ net1378 net1351 _1860_ VPWR VGND sg13g2_nor2b_1
X_7629_ VGND VPWR net1721 _3321_ _0107_ _3358_ sg13g2_a21oi_1
X_7742__279 VPWR VGND net279 sg13g2_tiehi
XFILLER_20_31 VPWR VGND sg13g2_fill_1
XFILLER_0_410 VPWR VGND sg13g2_decap_8
XFILLER_1_922 VPWR VGND sg13g2_decap_8
XFILLER_49_948 VPWR VGND sg13g2_decap_8
Xhold40 s0.was_valid_out\[23\][0] VPWR VGND net409 sg13g2_dlygate4sd3_1
XFILLER_1_999 VPWR VGND sg13g2_decap_8
Xhold73 _0313_ VPWR VGND net442 sg13g2_dlygate4sd3_1
Xhold51 _0133_ VPWR VGND net420 sg13g2_dlygate4sd3_1
Xhold62 s0.data_out\[25\]\[4\] VPWR VGND net431 sg13g2_dlygate4sd3_1
Xhold84 _0361_ VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold95 s0.data_out\[26\]\[2\] VPWR VGND net464 sg13g2_dlygate4sd3_1
XFILLER_29_694 VPWR VGND sg13g2_decap_8
XFILLER_17_878 VPWR VGND sg13g2_decap_8
XFILLER_17_889 VPWR VGND sg13g2_fill_2
XFILLER_8_543 VPWR VGND sg13g2_fill_2
XFILLER_4_793 VPWR VGND sg13g2_decap_8
X_4290_ _0114_ _0355_ _0356_ _3417_ net1578 VPWR VGND sg13g2_a22oi_1
XFILLER_39_414 VPWR VGND sg13g2_fill_1
XFILLER_6_1015 VPWR VGND sg13g2_decap_8
XFILLER_27_609 VPWR VGND sg13g2_fill_1
XFILLER_48_970 VPWR VGND sg13g2_decap_8
X_6931_ net1590 _2659_ _2739_ VPWR VGND sg13g2_nor2_1
X_6862_ _2543_ VPWR _2672_ VGND net1278 _3529_ sg13g2_o21ai_1
XFILLER_23_815 VPWR VGND sg13g2_fill_1
X_5813_ net1417 VPWR _1731_ VGND _1672_ _1730_ sg13g2_o21ai_1
X_7806__210 VPWR VGND net210 sg13g2_tiehi
X_6793_ _2615_ _2590_ _2589_ VPWR VGND sg13g2_nand2b_1
X_5744_ VGND VPWR net1417 _1666_ _1669_ _1668_ sg13g2_a21oi_1
X_5675_ net1427 VPWR _1607_ VGND _1570_ _1606_ sg13g2_o21ai_1
X_4626_ VGND VPWR _0659_ _0657_ net1660 sg13g2_or2_1
X_7414_ VPWR VGND _3138_ _3175_ _3174_ _3163_ _3176_ _3171_ sg13g2_a221oi_1
X_7345_ net1222 net1348 _3107_ VPWR VGND sg13g2_nor2b_1
X_7696__329 VPWR VGND net329 sg13g2_tiehi
X_4557_ VPWR _0142_ _0595_ VGND sg13g2_inv_1
X_4488_ _0531_ net1520 _0532_ _0533_ VPWR VGND sg13g2_a21o_1
X_7276_ _3040_ _3041_ _3050_ VPWR VGND sg13g2_nor2_1
X_6227_ VGND VPWR net1321 _2102_ _2104_ _2103_ sg13g2_a21oi_1
X_6158_ _2020_ _2022_ _2047_ VPWR VGND sg13g2_nor2b_1
XFILLER_46_918 VPWR VGND sg13g2_decap_8
X_5109_ _1092_ net1459 _1093_ _1094_ VPWR VGND sg13g2_a21o_1
X_6089_ _1978_ net551 net1386 VPWR VGND sg13g2_nand2b_1
XFILLER_39_992 VPWR VGND sg13g2_decap_8
XFILLER_26_620 VPWR VGND sg13g2_fill_2
XFILLER_41_623 VPWR VGND sg13g2_fill_1
XFILLER_41_612 VPWR VGND sg13g2_fill_2
XFILLER_41_667 VPWR VGND sg13g2_fill_2
Xoutput6 net6 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_796 VPWR VGND sg13g2_decap_8
XFILLER_49_745 VPWR VGND sg13g2_decap_8
XFILLER_17_642 VPWR VGND sg13g2_fill_2
XFILLER_17_664 VPWR VGND sg13g2_fill_1
XFILLER_45_984 VPWR VGND sg13g2_decap_8
XFILLER_12_380 VPWR VGND sg13g2_fill_2
X_5460_ s0.data_out\[17\]\[0\] s0.data_out\[16\]\[0\] net1432 _1409_ VPWR VGND sg13g2_mux2_1
X_4411_ _0126_ _0464_ _0465_ _3416_ net1579 VPWR VGND sg13g2_a22oi_1
X_5391_ net1693 _1315_ _1352_ VPWR VGND sg13g2_nor2_1
X_4342_ VGND VPWR net1552 _0396_ _0399_ _0398_ sg13g2_a21oi_1
X_7130_ _2916_ net1668 _2913_ _2915_ VPWR VGND sg13g2_and3_1
X_4273_ _3625_ VPWR _3637_ VGND net1687 _3594_ sg13g2_o21ai_1
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
X_7061_ net1596 _2798_ _2855_ VPWR VGND sg13g2_nor2_1
X_6012_ net1382 net1336 _1913_ VPWR VGND sg13g2_nor2b_1
.ends

