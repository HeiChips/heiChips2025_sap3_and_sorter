module heichips25_top_sorter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire \s0.data_new_delayed[0] ;
 wire \s0.data_new_delayed[1] ;
 wire \s0.data_new_delayed[2] ;
 wire \s0.data_new_delayed[3] ;
 wire \s0.data_new_delayed[4] ;
 wire \s0.data_new_delayed[5] ;
 wire \s0.data_new_delayed[6] ;
 wire \s0.data_new_delayed[7] ;
 wire \s0.data_out[0][0] ;
 wire \s0.data_out[0][1] ;
 wire \s0.data_out[0][2] ;
 wire \s0.data_out[0][3] ;
 wire \s0.data_out[0][4] ;
 wire \s0.data_out[0][5] ;
 wire \s0.data_out[0][6] ;
 wire \s0.data_out[0][7] ;
 wire \s0.data_out[10][0] ;
 wire \s0.data_out[10][1] ;
 wire \s0.data_out[10][2] ;
 wire \s0.data_out[10][3] ;
 wire \s0.data_out[10][4] ;
 wire \s0.data_out[10][5] ;
 wire \s0.data_out[10][6] ;
 wire \s0.data_out[10][7] ;
 wire \s0.data_out[11][0] ;
 wire \s0.data_out[11][1] ;
 wire \s0.data_out[11][2] ;
 wire \s0.data_out[11][3] ;
 wire \s0.data_out[11][4] ;
 wire \s0.data_out[11][5] ;
 wire \s0.data_out[11][6] ;
 wire \s0.data_out[11][7] ;
 wire \s0.data_out[12][0] ;
 wire \s0.data_out[12][1] ;
 wire \s0.data_out[12][2] ;
 wire \s0.data_out[12][3] ;
 wire \s0.data_out[12][4] ;
 wire \s0.data_out[12][5] ;
 wire \s0.data_out[12][6] ;
 wire \s0.data_out[12][7] ;
 wire \s0.data_out[13][0] ;
 wire \s0.data_out[13][1] ;
 wire \s0.data_out[13][2] ;
 wire \s0.data_out[13][3] ;
 wire \s0.data_out[13][4] ;
 wire \s0.data_out[13][5] ;
 wire \s0.data_out[13][6] ;
 wire \s0.data_out[13][7] ;
 wire \s0.data_out[14][0] ;
 wire \s0.data_out[14][1] ;
 wire \s0.data_out[14][2] ;
 wire \s0.data_out[14][3] ;
 wire \s0.data_out[14][4] ;
 wire \s0.data_out[14][5] ;
 wire \s0.data_out[14][6] ;
 wire \s0.data_out[14][7] ;
 wire \s0.data_out[15][0] ;
 wire \s0.data_out[15][1] ;
 wire \s0.data_out[15][2] ;
 wire \s0.data_out[15][3] ;
 wire \s0.data_out[15][4] ;
 wire \s0.data_out[15][5] ;
 wire \s0.data_out[15][6] ;
 wire \s0.data_out[15][7] ;
 wire \s0.data_out[16][0] ;
 wire \s0.data_out[16][1] ;
 wire \s0.data_out[16][2] ;
 wire \s0.data_out[16][3] ;
 wire \s0.data_out[16][4] ;
 wire \s0.data_out[16][5] ;
 wire \s0.data_out[16][6] ;
 wire \s0.data_out[16][7] ;
 wire \s0.data_out[17][0] ;
 wire \s0.data_out[17][1] ;
 wire \s0.data_out[17][2] ;
 wire \s0.data_out[17][3] ;
 wire \s0.data_out[17][4] ;
 wire \s0.data_out[17][5] ;
 wire \s0.data_out[17][6] ;
 wire \s0.data_out[17][7] ;
 wire \s0.data_out[18][0] ;
 wire \s0.data_out[18][1] ;
 wire \s0.data_out[18][2] ;
 wire \s0.data_out[18][3] ;
 wire \s0.data_out[18][4] ;
 wire \s0.data_out[18][5] ;
 wire \s0.data_out[18][6] ;
 wire \s0.data_out[18][7] ;
 wire \s0.data_out[19][0] ;
 wire \s0.data_out[19][1] ;
 wire \s0.data_out[19][2] ;
 wire \s0.data_out[19][3] ;
 wire \s0.data_out[19][4] ;
 wire \s0.data_out[19][5] ;
 wire \s0.data_out[19][6] ;
 wire \s0.data_out[19][7] ;
 wire \s0.data_out[1][0] ;
 wire \s0.data_out[1][1] ;
 wire \s0.data_out[1][2] ;
 wire \s0.data_out[1][3] ;
 wire \s0.data_out[1][4] ;
 wire \s0.data_out[1][5] ;
 wire \s0.data_out[1][6] ;
 wire \s0.data_out[1][7] ;
 wire \s0.data_out[20][0] ;
 wire \s0.data_out[20][1] ;
 wire \s0.data_out[20][2] ;
 wire \s0.data_out[20][3] ;
 wire \s0.data_out[20][4] ;
 wire \s0.data_out[20][5] ;
 wire \s0.data_out[20][6] ;
 wire \s0.data_out[20][7] ;
 wire \s0.data_out[21][0] ;
 wire \s0.data_out[21][1] ;
 wire \s0.data_out[21][2] ;
 wire \s0.data_out[21][3] ;
 wire \s0.data_out[21][4] ;
 wire \s0.data_out[21][5] ;
 wire \s0.data_out[21][6] ;
 wire \s0.data_out[21][7] ;
 wire \s0.data_out[22][0] ;
 wire \s0.data_out[22][1] ;
 wire \s0.data_out[22][2] ;
 wire \s0.data_out[22][3] ;
 wire \s0.data_out[22][4] ;
 wire \s0.data_out[22][5] ;
 wire \s0.data_out[22][6] ;
 wire \s0.data_out[22][7] ;
 wire \s0.data_out[23][0] ;
 wire \s0.data_out[23][1] ;
 wire \s0.data_out[23][2] ;
 wire \s0.data_out[23][3] ;
 wire \s0.data_out[23][4] ;
 wire \s0.data_out[23][5] ;
 wire \s0.data_out[23][6] ;
 wire \s0.data_out[23][7] ;
 wire \s0.data_out[24][0] ;
 wire \s0.data_out[24][1] ;
 wire \s0.data_out[24][2] ;
 wire \s0.data_out[24][3] ;
 wire \s0.data_out[24][4] ;
 wire \s0.data_out[24][5] ;
 wire \s0.data_out[24][6] ;
 wire \s0.data_out[24][7] ;
 wire \s0.data_out[25][0] ;
 wire \s0.data_out[25][1] ;
 wire \s0.data_out[25][2] ;
 wire \s0.data_out[25][3] ;
 wire \s0.data_out[25][4] ;
 wire \s0.data_out[25][5] ;
 wire \s0.data_out[25][6] ;
 wire \s0.data_out[25][7] ;
 wire \s0.data_out[26][0] ;
 wire \s0.data_out[26][1] ;
 wire \s0.data_out[26][2] ;
 wire \s0.data_out[26][3] ;
 wire \s0.data_out[26][4] ;
 wire \s0.data_out[26][5] ;
 wire \s0.data_out[26][6] ;
 wire \s0.data_out[26][7] ;
 wire \s0.data_out[27][0] ;
 wire \s0.data_out[27][1] ;
 wire \s0.data_out[27][2] ;
 wire \s0.data_out[27][3] ;
 wire \s0.data_out[27][4] ;
 wire \s0.data_out[27][5] ;
 wire \s0.data_out[27][6] ;
 wire \s0.data_out[27][7] ;
 wire \s0.data_out[2][0] ;
 wire \s0.data_out[2][1] ;
 wire \s0.data_out[2][2] ;
 wire \s0.data_out[2][3] ;
 wire \s0.data_out[2][4] ;
 wire \s0.data_out[2][5] ;
 wire \s0.data_out[2][6] ;
 wire \s0.data_out[2][7] ;
 wire \s0.data_out[3][0] ;
 wire \s0.data_out[3][1] ;
 wire \s0.data_out[3][2] ;
 wire \s0.data_out[3][3] ;
 wire \s0.data_out[3][4] ;
 wire \s0.data_out[3][5] ;
 wire \s0.data_out[3][6] ;
 wire \s0.data_out[3][7] ;
 wire \s0.data_out[4][0] ;
 wire \s0.data_out[4][1] ;
 wire \s0.data_out[4][2] ;
 wire \s0.data_out[4][3] ;
 wire \s0.data_out[4][4] ;
 wire \s0.data_out[4][5] ;
 wire \s0.data_out[4][6] ;
 wire \s0.data_out[4][7] ;
 wire \s0.data_out[5][0] ;
 wire \s0.data_out[5][1] ;
 wire \s0.data_out[5][2] ;
 wire \s0.data_out[5][3] ;
 wire \s0.data_out[5][4] ;
 wire \s0.data_out[5][5] ;
 wire \s0.data_out[5][6] ;
 wire \s0.data_out[5][7] ;
 wire \s0.data_out[6][0] ;
 wire \s0.data_out[6][1] ;
 wire \s0.data_out[6][2] ;
 wire \s0.data_out[6][3] ;
 wire \s0.data_out[6][4] ;
 wire \s0.data_out[6][5] ;
 wire \s0.data_out[6][6] ;
 wire \s0.data_out[6][7] ;
 wire \s0.data_out[7][0] ;
 wire \s0.data_out[7][1] ;
 wire \s0.data_out[7][2] ;
 wire \s0.data_out[7][3] ;
 wire \s0.data_out[7][4] ;
 wire \s0.data_out[7][5] ;
 wire \s0.data_out[7][6] ;
 wire \s0.data_out[7][7] ;
 wire \s0.data_out[8][0] ;
 wire \s0.data_out[8][1] ;
 wire \s0.data_out[8][2] ;
 wire \s0.data_out[8][3] ;
 wire \s0.data_out[8][4] ;
 wire \s0.data_out[8][5] ;
 wire \s0.data_out[8][6] ;
 wire \s0.data_out[8][7] ;
 wire \s0.data_out[9][0] ;
 wire \s0.data_out[9][1] ;
 wire \s0.data_out[9][2] ;
 wire \s0.data_out[9][3] ;
 wire \s0.data_out[9][4] ;
 wire \s0.data_out[9][5] ;
 wire \s0.data_out[9][6] ;
 wire \s0.data_out[9][7] ;
 wire \s0.genblk1[10].modules.bubble ;
 wire \s0.genblk1[11].modules.bubble ;
 wire \s0.genblk1[12].modules.bubble ;
 wire \s0.genblk1[13].modules.bubble ;
 wire \s0.genblk1[14].modules.bubble ;
 wire \s0.genblk1[15].modules.bubble ;
 wire \s0.genblk1[16].modules.bubble ;
 wire \s0.genblk1[17].modules.bubble ;
 wire \s0.genblk1[18].modules.bubble ;
 wire \s0.genblk1[19].modules.bubble ;
 wire \s0.genblk1[1].modules.bubble ;
 wire \s0.genblk1[20].modules.bubble ;
 wire \s0.genblk1[21].modules.bubble ;
 wire \s0.genblk1[22].modules.bubble ;
 wire \s0.genblk1[23].modules.bubble ;
 wire \s0.genblk1[24].modules.bubble ;
 wire \s0.genblk1[25].modules.bubble ;
 wire \s0.genblk1[26].modules.bubble ;
 wire \s0.genblk1[27].modules.bubble ;
 wire \s0.genblk1[2].modules.bubble ;
 wire \s0.genblk1[3].modules.bubble ;
 wire \s0.genblk1[4].modules.bubble ;
 wire \s0.genblk1[5].modules.bubble ;
 wire \s0.genblk1[6].modules.bubble ;
 wire \s0.genblk1[7].modules.bubble ;
 wire \s0.genblk1[8].modules.bubble ;
 wire \s0.genblk1[9].modules.bubble ;
 wire \s0.module0.bubble ;
 wire net12;
 wire net13;
 wire net369;
 wire net14;
 wire net15;
 wire clknet_leaf_0_clk;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1;
 wire net11;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire [0:0] \s0.shift_out[0] ;
 wire [0:0] \s0.shift_out[10] ;
 wire [0:0] \s0.shift_out[11] ;
 wire [0:0] \s0.shift_out[12] ;
 wire [0:0] \s0.shift_out[13] ;
 wire [0:0] \s0.shift_out[14] ;
 wire [0:0] \s0.shift_out[15] ;
 wire [0:0] \s0.shift_out[16] ;
 wire [0:0] \s0.shift_out[17] ;
 wire [0:0] \s0.shift_out[18] ;
 wire [0:0] \s0.shift_out[19] ;
 wire [0:0] \s0.shift_out[1] ;
 wire [0:0] \s0.shift_out[20] ;
 wire [0:0] \s0.shift_out[21] ;
 wire [0:0] \s0.shift_out[22] ;
 wire [0:0] \s0.shift_out[23] ;
 wire [0:0] \s0.shift_out[24] ;
 wire [0:0] \s0.shift_out[25] ;
 wire [0:0] \s0.shift_out[26] ;
 wire [0:0] \s0.shift_out[27] ;
 wire [0:0] \s0.shift_out[2] ;
 wire [0:0] \s0.shift_out[3] ;
 wire [0:0] \s0.shift_out[4] ;
 wire [0:0] \s0.shift_out[5] ;
 wire [0:0] \s0.shift_out[6] ;
 wire [0:0] \s0.shift_out[7] ;
 wire [0:0] \s0.shift_out[8] ;
 wire [0:0] \s0.shift_out[9] ;
 wire [0:0] \s0.valid_out[0] ;
 wire [0:0] \s0.valid_out[10] ;
 wire [0:0] \s0.valid_out[11] ;
 wire [0:0] \s0.valid_out[12] ;
 wire [0:0] \s0.valid_out[13] ;
 wire [0:0] \s0.valid_out[14] ;
 wire [0:0] \s0.valid_out[15] ;
 wire [0:0] \s0.valid_out[16] ;
 wire [0:0] \s0.valid_out[17] ;
 wire [0:0] \s0.valid_out[18] ;
 wire [0:0] \s0.valid_out[19] ;
 wire [0:0] \s0.valid_out[1] ;
 wire [0:0] \s0.valid_out[20] ;
 wire [0:0] \s0.valid_out[21] ;
 wire [0:0] \s0.valid_out[22] ;
 wire [0:0] \s0.valid_out[23] ;
 wire [0:0] \s0.valid_out[24] ;
 wire [0:0] \s0.valid_out[25] ;
 wire [0:0] \s0.valid_out[26] ;
 wire [0:0] \s0.valid_out[27] ;
 wire [0:0] \s0.valid_out[2] ;
 wire [0:0] \s0.valid_out[3] ;
 wire [0:0] \s0.valid_out[4] ;
 wire [0:0] \s0.valid_out[5] ;
 wire [0:0] \s0.valid_out[6] ;
 wire [0:0] \s0.valid_out[7] ;
 wire [0:0] \s0.valid_out[8] ;
 wire [0:0] \s0.valid_out[9] ;
 wire [0:0] \s0.was_valid_out[0] ;
 wire [0:0] \s0.was_valid_out[10] ;
 wire [0:0] \s0.was_valid_out[11] ;
 wire [0:0] \s0.was_valid_out[12] ;
 wire [0:0] \s0.was_valid_out[13] ;
 wire [0:0] \s0.was_valid_out[14] ;
 wire [0:0] \s0.was_valid_out[15] ;
 wire [0:0] \s0.was_valid_out[16] ;
 wire [0:0] \s0.was_valid_out[17] ;
 wire [0:0] \s0.was_valid_out[18] ;
 wire [0:0] \s0.was_valid_out[19] ;
 wire [0:0] \s0.was_valid_out[1] ;
 wire [0:0] \s0.was_valid_out[20] ;
 wire [0:0] \s0.was_valid_out[21] ;
 wire [0:0] \s0.was_valid_out[22] ;
 wire [0:0] \s0.was_valid_out[23] ;
 wire [0:0] \s0.was_valid_out[24] ;
 wire [0:0] \s0.was_valid_out[25] ;
 wire [0:0] \s0.was_valid_out[26] ;
 wire [0:0] \s0.was_valid_out[27] ;
 wire [0:0] \s0.was_valid_out[2] ;
 wire [0:0] \s0.was_valid_out[3] ;
 wire [0:0] \s0.was_valid_out[4] ;
 wire [0:0] \s0.was_valid_out[5] ;
 wire [0:0] \s0.was_valid_out[6] ;
 wire [0:0] \s0.was_valid_out[7] ;
 wire [0:0] \s0.was_valid_out[8] ;
 wire [0:0] \s0.was_valid_out[9] ;

 sg13g2_inv_1 _3983_ (.Y(_3359_),
    .A(net432));
 sg13g2_inv_1 _3984_ (.Y(_3360_),
    .A(net406));
 sg13g2_inv_1 _3985_ (.Y(_3361_),
    .A(net416));
 sg13g2_inv_1 _3986_ (.Y(_3362_),
    .A(net434));
 sg13g2_inv_1 _3987_ (.Y(_3363_),
    .A(net422));
 sg13g2_inv_1 _3988_ (.Y(_3364_),
    .A(net439));
 sg13g2_inv_1 _3989_ (.Y(_3365_),
    .A(net398));
 sg13g2_inv_1 _3990_ (.Y(_3366_),
    .A(net420));
 sg13g2_inv_1 _3991_ (.Y(_3367_),
    .A(net409));
 sg13g2_inv_1 _3992_ (.Y(_3368_),
    .A(net400));
 sg13g2_inv_1 _3993_ (.Y(_3369_),
    .A(net411));
 sg13g2_inv_1 _3994_ (.Y(_3370_),
    .A(net412));
 sg13g2_inv_1 _3995_ (.Y(_3371_),
    .A(net418));
 sg13g2_inv_1 _3996_ (.Y(_3372_),
    .A(net506));
 sg13g2_inv_1 _3997_ (.Y(_3373_),
    .A(net1630));
 sg13g2_inv_1 _3998_ (.Y(_3374_),
    .A(net1723));
 sg13g2_inv_2 _3999_ (.Y(_3375_),
    .A(net1434));
 sg13g2_inv_1 _4000_ (.Y(_3376_),
    .A(net1425));
 sg13g2_inv_1 _4001_ (.Y(_3377_),
    .A(net1445));
 sg13g2_inv_1 _4002_ (.Y(_3378_),
    .A(net1212));
 sg13g2_inv_1 _4003_ (.Y(_3379_),
    .A(net1455));
 sg13g2_inv_2 _4004_ (.Y(_3380_),
    .A(net1408));
 sg13g2_inv_2 _4005_ (.Y(_3381_),
    .A(net1396));
 sg13g2_inv_1 _4006_ (.Y(_3382_),
    .A(net1384));
 sg13g2_inv_4 _4007_ (.A(net1358),
    .Y(_3383_));
 sg13g2_inv_1 _4008_ (.Y(_3384_),
    .A(net1235));
 sg13g2_inv_1 _4009_ (.Y(_3385_),
    .A(net454));
 sg13g2_inv_1 _4010_ (.Y(_3386_),
    .A(net1552));
 sg13g2_inv_1 _4011_ (.Y(_3387_),
    .A(net1222));
 sg13g2_inv_1 _4012_ (.Y(_3388_),
    .A(net1524));
 sg13g2_inv_2 _4013_ (.Y(_3389_),
    .A(net1521));
 sg13g2_inv_1 _4014_ (.Y(_3390_),
    .A(net1504));
 sg13g2_inv_1 _4015_ (.Y(_3391_),
    .A(net1480));
 sg13g2_inv_2 _4016_ (.Y(_3392_),
    .A(net1472));
 sg13g2_inv_4 _4017_ (.A(net1202),
    .Y(_3393_));
 sg13g2_inv_4 _4018_ (.A(net1289),
    .Y(_3394_));
 sg13g2_inv_2 _4019_ (.Y(_3395_),
    .A(net1278));
 sg13g2_inv_4 _4020_ (.A(net1268),
    .Y(_3396_));
 sg13g2_inv_1 _4021_ (.Y(_3397_),
    .A(net1239));
 sg13g2_inv_1 _4022_ (.Y(_3398_),
    .A(net536));
 sg13g2_inv_1 _4023_ (.Y(_3399_),
    .A(net612));
 sg13g2_inv_1 _4024_ (.Y(_3400_),
    .A(net486));
 sg13g2_inv_1 _4025_ (.Y(_3401_),
    .A(net1325));
 sg13g2_inv_2 _4026_ (.Y(_3402_),
    .A(net1646));
 sg13g2_inv_4 _4027_ (.A(net1658),
    .Y(_3403_));
 sg13g2_inv_1 _4028_ (.Y(_3404_),
    .A(net512));
 sg13g2_inv_1 _4029_ (.Y(_3405_),
    .A(net467));
 sg13g2_inv_8 _4030_ (.Y(_3406_),
    .A(net1665));
 sg13g2_inv_1 _4031_ (.Y(_3407_),
    .A(net511));
 sg13g2_inv_1 _4032_ (.Y(_3408_),
    .A(net463));
 sg13g2_inv_2 _4033_ (.Y(_3409_),
    .A(net824));
 sg13g2_inv_2 _4034_ (.Y(_3410_),
    .A(net456));
 sg13g2_inv_1 _4035_ (.Y(_3411_),
    .A(net1339));
 sg13g2_inv_1 _4036_ (.Y(_3412_),
    .A(net477));
 sg13g2_inv_1 _4037_ (.Y(_3413_),
    .A(net507));
 sg13g2_inv_1 _4038_ (.Y(_3414_),
    .A(net1684));
 sg13g2_inv_2 _4039_ (.Y(_3415_),
    .A(net1690));
 sg13g2_inv_1 _4040_ (.Y(_3416_),
    .A(net670));
 sg13g2_inv_1 _4041_ (.Y(_3417_),
    .A(net600));
 sg13g2_inv_1 _4042_ (.Y(_3418_),
    .A(net1700));
 sg13g2_inv_1 _4043_ (.Y(_3419_),
    .A(net524));
 sg13g2_inv_2 _4044_ (.Y(_3420_),
    .A(net556));
 sg13g2_inv_1 _4045_ (.Y(_3421_),
    .A(net767));
 sg13g2_inv_1 _4046_ (.Y(_3422_),
    .A(net775));
 sg13g2_inv_1 _4047_ (.Y(_3423_),
    .A(\s0.data_out[25][2] ));
 sg13g2_inv_1 _4048_ (.Y(_3424_),
    .A(net548));
 sg13g2_inv_1 _4049_ (.Y(_3425_),
    .A(net540));
 sg13g2_inv_1 _4050_ (.Y(_3426_),
    .A(net554));
 sg13g2_inv_1 _4051_ (.Y(_3427_),
    .A(net429));
 sg13g2_inv_1 _4052_ (.Y(_3428_),
    .A(net592));
 sg13g2_inv_1 _4053_ (.Y(_3429_),
    .A(net502));
 sg13g2_inv_1 _4054_ (.Y(_3430_),
    .A(net631));
 sg13g2_inv_1 _4055_ (.Y(_3431_),
    .A(net509));
 sg13g2_inv_1 _4056_ (.Y(_3432_),
    .A(net727));
 sg13g2_inv_1 _4057_ (.Y(_3433_),
    .A(net570));
 sg13g2_inv_1 _4058_ (.Y(_3434_),
    .A(net802));
 sg13g2_inv_1 _4059_ (.Y(_3435_),
    .A(\s0.data_out[23][2] ));
 sg13g2_inv_1 _4060_ (.Y(_3436_),
    .A(net817));
 sg13g2_inv_1 _4061_ (.Y(_3437_),
    .A(net526));
 sg13g2_inv_1 _4062_ (.Y(_3438_),
    .A(net488));
 sg13g2_inv_1 _4063_ (.Y(_3439_),
    .A(net611));
 sg13g2_inv_1 _4064_ (.Y(_3440_),
    .A(net658));
 sg13g2_inv_1 _4065_ (.Y(_3441_),
    .A(net544));
 sg13g2_inv_1 _4066_ (.Y(_3442_),
    .A(net449));
 sg13g2_inv_1 _4067_ (.Y(_3443_),
    .A(net499));
 sg13g2_inv_2 _4068_ (.Y(_3444_),
    .A(\s0.data_out[21][2] ));
 sg13g2_inv_1 _4069_ (.Y(_3445_),
    .A(net694));
 sg13g2_inv_1 _4070_ (.Y(_3446_),
    .A(net492));
 sg13g2_inv_2 _4071_ (.Y(_3447_),
    .A(net516));
 sg13g2_inv_1 _4072_ (.Y(_3448_),
    .A(net644));
 sg13g2_inv_1 _4073_ (.Y(_3449_),
    .A(net691));
 sg13g2_inv_2 _4074_ (.Y(_3450_),
    .A(net560));
 sg13g2_inv_1 _4075_ (.Y(_3451_),
    .A(net755));
 sg13g2_inv_1 _4076_ (.Y(_3452_),
    .A(net764));
 sg13g2_inv_1 _4077_ (.Y(_3453_),
    .A(net790));
 sg13g2_inv_2 _4078_ (.Y(_3454_),
    .A(net656));
 sg13g2_inv_1 _4079_ (.Y(_3455_),
    .A(net662));
 sg13g2_inv_1 _4080_ (.Y(_3456_),
    .A(net725));
 sg13g2_inv_1 _4081_ (.Y(_3457_),
    .A(net805));
 sg13g2_inv_1 _4082_ (.Y(_3458_),
    .A(net574));
 sg13g2_inv_2 _4083_ (.Y(_3459_),
    .A(net598));
 sg13g2_inv_1 _4084_ (.Y(_3460_),
    .A(net482));
 sg13g2_inv_1 _4085_ (.Y(_3461_),
    .A(net627));
 sg13g2_inv_1 _4086_ (.Y(_3462_),
    .A(net582));
 sg13g2_inv_1 _4087_ (.Y(_3463_),
    .A(net819));
 sg13g2_inv_2 _4088_ (.Y(_3464_),
    .A(\s0.data_out[17][2] ));
 sg13g2_inv_1 _4089_ (.Y(_3465_),
    .A(net823));
 sg13g2_inv_1 _4090_ (.Y(_3466_),
    .A(net538));
 sg13g2_inv_1 _4091_ (.Y(_3467_),
    .A(net465));
 sg13g2_inv_1 _4092_ (.Y(_3468_),
    .A(net716));
 sg13g2_inv_1 _4093_ (.Y(_3469_),
    .A(net471));
 sg13g2_inv_1 _4094_ (.Y(_3470_),
    .A(net564));
 sg13g2_inv_1 _4095_ (.Y(_3471_),
    .A(net484));
 sg13g2_inv_1 _4096_ (.Y(_3472_),
    .A(net578));
 sg13g2_inv_1 _4097_ (.Y(_3473_),
    .A(net786));
 sg13g2_inv_1 _4098_ (.Y(_3474_),
    .A(\s0.data_out[15][2] ));
 sg13g2_inv_1 _4099_ (.Y(_3475_),
    .A(net814));
 sg13g2_inv_1 _4100_ (.Y(_3476_),
    .A(net712));
 sg13g2_inv_1 _4101_ (.Y(_3477_),
    .A(net783));
 sg13g2_inv_1 _4102_ (.Y(_3478_),
    .A(\s0.data_out[14][4] ));
 sg13g2_inv_1 _4103_ (.Y(_3479_),
    .A(net730));
 sg13g2_inv_1 _4104_ (.Y(_3480_),
    .A(net648));
 sg13g2_inv_1 _4105_ (.Y(_3481_),
    .A(net729));
 sg13g2_inv_1 _4106_ (.Y(_3482_),
    .A(net608));
 sg13g2_inv_1 _4107_ (.Y(_3483_),
    .A(net583));
 sg13g2_inv_2 _4108_ (.Y(_3484_),
    .A(net518));
 sg13g2_inv_1 _4109_ (.Y(_3485_),
    .A(net692));
 sg13g2_inv_1 _4110_ (.Y(_3486_),
    .A(\s0.data_out[13][2] ));
 sg13g2_inv_1 _4111_ (.Y(_3487_),
    .A(net522));
 sg13g2_inv_1 _4112_ (.Y(_3488_),
    .A(net660));
 sg13g2_inv_1 _4113_ (.Y(_3489_),
    .A(net580));
 sg13g2_inv_1 _4114_ (.Y(_3490_),
    .A(net749));
 sg13g2_inv_1 _4115_ (.Y(_3491_),
    .A(net820));
 sg13g2_inv_1 _4116_ (.Y(_3492_),
    .A(net753));
 sg13g2_inv_1 _4117_ (.Y(_3493_),
    .A(net746));
 sg13g2_inv_1 _4118_ (.Y(_3494_),
    .A(net571));
 sg13g2_inv_1 _4119_ (.Y(_3495_),
    .A(net568));
 sg13g2_inv_1 _4120_ (.Y(_3496_),
    .A(net605));
 sg13g2_inv_1 _4121_ (.Y(_3497_),
    .A(net788));
 sg13g2_inv_1 _4122_ (.Y(_3498_),
    .A(net659));
 sg13g2_inv_1 _4123_ (.Y(_3499_),
    .A(net436));
 sg13g2_inv_1 _4124_ (.Y(_3500_),
    .A(net479));
 sg13g2_inv_1 _4125_ (.Y(_3501_),
    .A(net514));
 sg13g2_inv_1 _4126_ (.Y(_3502_),
    .A(net497));
 sg13g2_inv_1 _4127_ (.Y(_3503_),
    .A(net534));
 sg13g2_inv_1 _4128_ (.Y(_3504_),
    .A(net664));
 sg13g2_inv_1 _4129_ (.Y(_3505_),
    .A(net490));
 sg13g2_inv_1 _4130_ (.Y(_3506_),
    .A(net475));
 sg13g2_inv_1 _4131_ (.Y(_3507_),
    .A(net553));
 sg13g2_inv_1 _4132_ (.Y(_3508_),
    .A(net640));
 sg13g2_inv_1 _4133_ (.Y(_3509_),
    .A(net813));
 sg13g2_inv_1 _4134_ (.Y(_3510_),
    .A(net773));
 sg13g2_inv_1 _4135_ (.Y(_3511_),
    .A(net610));
 sg13g2_inv_1 _4136_ (.Y(_3512_),
    .A(net562));
 sg13g2_inv_1 _4137_ (.Y(_3513_),
    .A(net594));
 sg13g2_inv_1 _4138_ (.Y(_3514_),
    .A(net796));
 sg13g2_inv_1 _4139_ (.Y(_3515_),
    .A(net576));
 sg13g2_inv_1 _4140_ (.Y(_3516_),
    .A(net590));
 sg13g2_inv_1 _4141_ (.Y(_3517_),
    .A(net460));
 sg13g2_inv_1 _4142_ (.Y(_3518_),
    .A(net740));
 sg13g2_inv_1 _4143_ (.Y(_3519_),
    .A(net668));
 sg13g2_inv_1 _4144_ (.Y(_3520_),
    .A(net779));
 sg13g2_inv_1 _4145_ (.Y(_3521_),
    .A(\s0.data_out[6][3] ));
 sg13g2_inv_1 _4146_ (.Y(_3522_),
    .A(net549));
 sg13g2_inv_1 _4147_ (.Y(_3523_),
    .A(net737));
 sg13g2_inv_1 _4148_ (.Y(_3524_),
    .A(net528));
 sg13g2_inv_1 _4149_ (.Y(_3525_),
    .A(net596));
 sg13g2_inv_1 _4150_ (.Y(_3526_),
    .A(net651));
 sg13g2_inv_1 _4151_ (.Y(_3527_),
    .A(net751));
 sg13g2_inv_1 _4152_ (.Y(_3528_),
    .A(net572));
 sg13g2_inv_1 _4153_ (.Y(_3529_),
    .A(net646));
 sg13g2_inv_1 _4154_ (.Y(_3530_),
    .A(net546));
 sg13g2_inv_1 _4155_ (.Y(_3531_),
    .A(net624));
 sg13g2_inv_1 _4156_ (.Y(_3532_),
    .A(net558));
 sg13g2_inv_1 _4157_ (.Y(_3533_),
    .A(net495));
 sg13g2_inv_1 _4158_ (.Y(_3534_),
    .A(net501));
 sg13g2_inv_1 _4159_ (.Y(_3535_),
    .A(net634));
 sg13g2_inv_1 _4160_ (.Y(_3536_),
    .A(net812));
 sg13g2_inv_1 _4161_ (.Y(_3537_),
    .A(net700));
 sg13g2_inv_1 _4162_ (.Y(_3538_),
    .A(net542));
 sg13g2_inv_1 _4163_ (.Y(_3539_),
    .A(net424));
 sg13g2_inv_1 _4164_ (.Y(_3540_),
    .A(net784));
 sg13g2_inv_1 _4165_ (.Y(_3541_),
    .A(\s0.data_out[1][5] ));
 sg13g2_inv_1 _4166_ (.Y(_3542_),
    .A(net736));
 sg13g2_inv_1 _4167_ (.Y(_3543_),
    .A(\s0.data_out[0][3] ));
 sg13g2_nor2_2 _4168_ (.A(\s0.was_valid_out[27] [0]),
    .B(net1551),
    .Y(_3544_));
 sg13g2_nor2_1 _4169_ (.A(\s0.data_out[27][0] ),
    .B(net1159),
    .Y(_3545_));
 sg13g2_a21oi_1 _4170_ (.A1(net1559),
    .A2(net1158),
    .Y(net3),
    .B1(_3545_));
 sg13g2_nor2_1 _4171_ (.A(\s0.data_out[27][1] ),
    .B(net1159),
    .Y(_3546_));
 sg13g2_a21oi_1 _4172_ (.A1(_3415_),
    .A2(net1158),
    .Y(net4),
    .B1(_3546_));
 sg13g2_nor2_1 _4173_ (.A(\s0.data_out[27][2] ),
    .B(net1159),
    .Y(_3547_));
 sg13g2_a21oi_1 _4174_ (.A1(net1560),
    .A2(net1159),
    .Y(net5),
    .B1(_3547_));
 sg13g2_nand2_1 _4175_ (.Y(_3548_),
    .A(net1675),
    .B(net1158));
 sg13g2_o21ai_1 _4176_ (.B1(_3548_),
    .Y(net6),
    .A1(_3410_),
    .A2(net1158));
 sg13g2_nor2_1 _4177_ (.A(\s0.data_out[27][4] ),
    .B(_3544_),
    .Y(_3549_));
 sg13g2_a21oi_1 _4178_ (.A1(_3406_),
    .A2(net1159),
    .Y(net7),
    .B1(_3549_));
 sg13g2_nor2_1 _4179_ (.A(\s0.data_out[27][5] ),
    .B(net1159),
    .Y(_3550_));
 sg13g2_a21oi_1 _4180_ (.A1(_3403_),
    .A2(net1159),
    .Y(net8),
    .B1(_3550_));
 sg13g2_nor2_1 _4181_ (.A(\s0.data_out[27][6] ),
    .B(net1158),
    .Y(_3551_));
 sg13g2_a21oi_1 _4182_ (.A1(_3402_),
    .A2(net1158),
    .Y(net9),
    .B1(_3551_));
 sg13g2_nand2_1 _4183_ (.Y(_3552_),
    .A(net1637),
    .B(net1158));
 sg13g2_o21ai_1 _4184_ (.B1(_3552_),
    .Y(net10),
    .A1(_3399_),
    .A2(net1158));
 sg13g2_and2_1 _4185_ (.A(net1709),
    .B(net384),
    .X(_0108_));
 sg13g2_o21ai_1 _4186_ (.B1(net1549),
    .Y(_3553_),
    .A1(net1627),
    .A2(net1535));
 sg13g2_a21oi_1 _4187_ (.A1(net1621),
    .A2(net1545),
    .Y(_3554_),
    .B1(_3553_));
 sg13g2_a21oi_1 _4188_ (.A1(net1621),
    .A2(net1553),
    .Y(_3555_),
    .B1(net1549));
 sg13g2_or2_1 _4189_ (.X(_3556_),
    .B(_3555_),
    .A(_3554_));
 sg13g2_o21ai_1 _4190_ (.B1(_3554_),
    .Y(_3557_),
    .A1(net506),
    .A2(net1545));
 sg13g2_nor2_1 _4191_ (.A(net1535),
    .B(_3553_),
    .Y(_3558_));
 sg13g2_a21oi_1 _4192_ (.A1(_3372_),
    .A2(_3385_),
    .Y(_3559_),
    .B1(net1549));
 sg13g2_nor2_1 _4193_ (.A(_3558_),
    .B(_3559_),
    .Y(_3560_));
 sg13g2_o21ai_1 _4194_ (.B1(net1704),
    .Y(_3561_),
    .A1(net769),
    .A2(_3556_));
 sg13g2_a21oi_1 _4195_ (.A1(_3557_),
    .A2(_3560_),
    .Y(_0109_),
    .B1(_3561_));
 sg13g2_nor2_1 _4196_ (.A(net1564),
    .B(_3556_),
    .Y(_0110_));
 sg13g2_and2_1 _4197_ (.A(net1704),
    .B(net371),
    .X(_0111_));
 sg13g2_o21ai_1 _4198_ (.B1(_3386_),
    .Y(_3562_),
    .A1(net1554),
    .A2(net477));
 sg13g2_a21oi_1 _4199_ (.A1(net1554),
    .A2(_3413_),
    .Y(_3563_),
    .B1(_3562_));
 sg13g2_nand2_1 _4200_ (.Y(_3564_),
    .A(net1546),
    .B(net477));
 sg13g2_o21ai_1 _4201_ (.B1(_3564_),
    .Y(_3565_),
    .A1(net1546),
    .A2(_3413_));
 sg13g2_nor2b_1 _4202_ (.A(net1537),
    .B_N(net1340),
    .Y(_3566_));
 sg13g2_a21o_1 _4203_ (.A2(_3565_),
    .A1(net1538),
    .B1(_3566_),
    .X(_3567_));
 sg13g2_a21oi_1 _4204_ (.A1(net1551),
    .A2(_3567_),
    .Y(_3568_),
    .B1(_3563_));
 sg13g2_nor2_1 _4205_ (.A(net1684),
    .B(_3568_),
    .Y(_3569_));
 sg13g2_o21ai_1 _4206_ (.B1(_3386_),
    .Y(_3570_),
    .A1(net1554),
    .A2(\s0.data_out[26][1] ));
 sg13g2_a21oi_1 _4207_ (.A1(net454),
    .A2(_3417_),
    .Y(_3571_),
    .B1(_3570_));
 sg13g2_nand2_1 _4208_ (.Y(_3572_),
    .A(net1546),
    .B(net670));
 sg13g2_o21ai_1 _4209_ (.B1(_3572_),
    .Y(_3573_),
    .A1(net1545),
    .A2(_3417_));
 sg13g2_nor2b_1 _4210_ (.A(net1537),
    .B_N(net1344),
    .Y(_3574_));
 sg13g2_a21o_1 _4211_ (.A2(_3573_),
    .A1(net1537),
    .B1(_3574_),
    .X(_3575_));
 sg13g2_a21oi_1 _4212_ (.A1(net1551),
    .A2(_3575_),
    .Y(_3576_),
    .B1(_3571_));
 sg13g2_nand2_1 _4213_ (.Y(_3577_),
    .A(net1690),
    .B(_3576_));
 sg13g2_o21ai_1 _4214_ (.B1(_3386_),
    .Y(_3578_),
    .A1(net1554),
    .A2(\s0.data_out[26][0] ));
 sg13g2_a21oi_1 _4215_ (.A1(net1554),
    .A2(_3419_),
    .Y(_3579_),
    .B1(_3578_));
 sg13g2_nor2b_1 _4216_ (.A(net1537),
    .B_N(net1348),
    .Y(_3580_));
 sg13g2_nand2_1 _4217_ (.Y(_3581_),
    .A(net1548),
    .B(\s0.data_out[26][0] ));
 sg13g2_mux2_1 _4218_ (.A0(\s0.data_out[27][0] ),
    .A1(\s0.data_out[26][0] ),
    .S(net1546),
    .X(_3582_));
 sg13g2_a21oi_1 _4219_ (.A1(net1537),
    .A2(_3582_),
    .Y(_3583_),
    .B1(_3580_));
 sg13g2_nor2b_1 _4220_ (.A(_3583_),
    .B_N(net1551),
    .Y(_3584_));
 sg13g2_o21ai_1 _4221_ (.B1(net1559),
    .Y(_3585_),
    .A1(_3579_),
    .A2(_3584_));
 sg13g2_o21ai_1 _4222_ (.B1(_3585_),
    .Y(_3586_),
    .A1(net1690),
    .A2(_3576_));
 sg13g2_a21oi_1 _4223_ (.A1(_3577_),
    .A2(_3586_),
    .Y(_3587_),
    .B1(_3569_));
 sg13g2_a21o_1 _4224_ (.A2(_3409_),
    .A1(_3385_),
    .B1(net1552),
    .X(_3588_));
 sg13g2_a21oi_1 _4225_ (.A1(net1554),
    .A2(_3410_),
    .Y(_3589_),
    .B1(_3588_));
 sg13g2_nand2_1 _4226_ (.Y(_3590_),
    .A(net1545),
    .B(net824));
 sg13g2_o21ai_1 _4227_ (.B1(_3590_),
    .Y(_3591_),
    .A1(net1546),
    .A2(_3410_));
 sg13g2_nor2_1 _4228_ (.A(net1538),
    .B(net1160),
    .Y(_3592_));
 sg13g2_a21o_1 _4229_ (.A2(_3591_),
    .A1(net1537),
    .B1(_3592_),
    .X(_3593_));
 sg13g2_a21oi_1 _4230_ (.A1(net1551),
    .A2(_3593_),
    .Y(_3594_),
    .B1(_3589_));
 sg13g2_a22oi_1 _4231_ (.Y(_3595_),
    .B1(_3594_),
    .B2(net1675),
    .A2(_3568_),
    .A1(net1684));
 sg13g2_inv_1 _4232_ (.Y(_3596_),
    .A(_3595_));
 sg13g2_nor2b_1 _4233_ (.A(net612),
    .B_N(net1553),
    .Y(_3597_));
 sg13g2_nor2_1 _4234_ (.A(net1553),
    .B(net536),
    .Y(_3598_));
 sg13g2_nor3_1 _4235_ (.A(net1550),
    .B(_3597_),
    .C(_3598_),
    .Y(_3599_));
 sg13g2_nand2_1 _4236_ (.Y(_3600_),
    .A(net1547),
    .B(net536));
 sg13g2_mux2_1 _4237_ (.A0(\s0.data_out[27][7] ),
    .A1(\s0.data_out[26][7] ),
    .S(net1545),
    .X(_3601_));
 sg13g2_nor2b_1 _4238_ (.A(net1535),
    .B_N(net1320),
    .Y(_3602_));
 sg13g2_a21o_1 _4239_ (.A2(_3601_),
    .A1(net1535),
    .B1(_3602_),
    .X(_3603_));
 sg13g2_a21oi_1 _4240_ (.A1(net1550),
    .A2(_3603_),
    .Y(_3604_),
    .B1(_3599_));
 sg13g2_nor2b_1 _4241_ (.A(net486),
    .B_N(net1553),
    .Y(_3605_));
 sg13g2_nor2_1 _4242_ (.A(net1553),
    .B(\s0.data_out[26][6] ),
    .Y(_3606_));
 sg13g2_nor3_1 _4243_ (.A(net1550),
    .B(_3605_),
    .C(_3606_),
    .Y(_3607_));
 sg13g2_nand2_1 _4244_ (.Y(_3608_),
    .A(net1547),
    .B(net680));
 sg13g2_mux2_1 _4245_ (.A0(\s0.data_out[27][6] ),
    .A1(\s0.data_out[26][6] ),
    .S(net1545),
    .X(_3609_));
 sg13g2_nor2b_1 _4246_ (.A(net1535),
    .B_N(net1325),
    .Y(_3610_));
 sg13g2_a21o_1 _4247_ (.A2(_3609_),
    .A1(net1535),
    .B1(_3610_),
    .X(_3611_));
 sg13g2_a21oi_1 _4248_ (.A1(net1550),
    .A2(_3611_),
    .Y(_3612_),
    .B1(_3607_));
 sg13g2_a22oi_1 _4249_ (.Y(_3613_),
    .B1(_3612_),
    .B2(net1646),
    .A2(_3604_),
    .A1(net1637));
 sg13g2_nor2_1 _4250_ (.A(net1637),
    .B(_3604_),
    .Y(_3614_));
 sg13g2_or2_1 _4251_ (.X(_3615_),
    .B(_3612_),
    .A(net1646));
 sg13g2_nand3b_1 _4252_ (.B(_3615_),
    .C(_3613_),
    .Y(_3616_),
    .A_N(_3614_));
 sg13g2_nor2b_1 _4253_ (.A(net467),
    .B_N(net1553),
    .Y(_3617_));
 sg13g2_nor2_1 _4254_ (.A(net1554),
    .B(\s0.data_out[26][5] ),
    .Y(_3618_));
 sg13g2_nor3_1 _4255_ (.A(net1549),
    .B(_3617_),
    .C(_3618_),
    .Y(_3619_));
 sg13g2_nand2_1 _4256_ (.Y(_3620_),
    .A(net1547),
    .B(net512));
 sg13g2_mux2_1 _4257_ (.A0(\s0.data_out[27][5] ),
    .A1(\s0.data_out[26][5] ),
    .S(net1545),
    .X(_3621_));
 sg13g2_nor2b_1 _4258_ (.A(net1536),
    .B_N(net1330),
    .Y(_3622_));
 sg13g2_a21o_1 _4259_ (.A2(_3621_),
    .A1(net1536),
    .B1(_3622_),
    .X(_3623_));
 sg13g2_a21oi_1 _4260_ (.A1(net1549),
    .A2(_3623_),
    .Y(_3624_),
    .B1(_3619_));
 sg13g2_nand2_1 _4261_ (.Y(_3625_),
    .A(net1655),
    .B(_3624_));
 sg13g2_nor2b_1 _4262_ (.A(net463),
    .B_N(net1553),
    .Y(_3626_));
 sg13g2_nor2_1 _4263_ (.A(net1553),
    .B(\s0.data_out[26][4] ),
    .Y(_3627_));
 sg13g2_nor3_1 _4264_ (.A(net1550),
    .B(_3626_),
    .C(_3627_),
    .Y(_3628_));
 sg13g2_nand2_1 _4265_ (.Y(_3629_),
    .A(net1547),
    .B(net511));
 sg13g2_mux2_1 _4266_ (.A0(\s0.data_out[27][4] ),
    .A1(\s0.data_out[26][4] ),
    .S(net1545),
    .X(_3630_));
 sg13g2_nor2b_1 _4267_ (.A(net1542),
    .B_N(net1335),
    .Y(_3631_));
 sg13g2_a21o_1 _4268_ (.A2(_3630_),
    .A1(net1536),
    .B1(_3631_),
    .X(_3632_));
 sg13g2_a21oi_1 _4269_ (.A1(net1549),
    .A2(_3632_),
    .Y(_3633_),
    .B1(_3628_));
 sg13g2_and2_1 _4270_ (.A(net1665),
    .B(_3633_),
    .X(_3634_));
 sg13g2_or2_1 _4271_ (.X(_3635_),
    .B(_3624_),
    .A(net1655));
 sg13g2_o21ai_1 _4272_ (.B1(_3635_),
    .Y(_3636_),
    .A1(net1665),
    .A2(_3633_));
 sg13g2_o21ai_1 _4273_ (.B1(_3625_),
    .Y(_3637_),
    .A1(net1675),
    .A2(_3594_));
 sg13g2_nor4_1 _4274_ (.A(_3616_),
    .B(_3634_),
    .C(_3636_),
    .D(_3637_),
    .Y(_3638_));
 sg13g2_o21ai_1 _4275_ (.B1(_3638_),
    .Y(_0344_),
    .A1(_3587_),
    .A2(_3596_));
 sg13g2_nand2_1 _4276_ (.Y(_0345_),
    .A(_3634_),
    .B(_3635_));
 sg13g2_a21oi_1 _4277_ (.A1(_3625_),
    .A2(_0345_),
    .Y(_0346_),
    .B1(_3616_));
 sg13g2_nor2_1 _4278_ (.A(_3613_),
    .B(_3614_),
    .Y(_0347_));
 sg13g2_nor3_1 _4279_ (.A(_3556_),
    .B(_0346_),
    .C(_0347_),
    .Y(_0348_));
 sg13g2_nand2_2 _4280_ (.Y(_0349_),
    .A(net1626),
    .B(net1705));
 sg13g2_or2_1 _4281_ (.X(_0350_),
    .B(net1555),
    .A(net383));
 sg13g2_a21oi_1 _4282_ (.A1(_0344_),
    .A2(_0348_),
    .Y(_0112_),
    .B1(_0350_));
 sg13g2_and2_1 _4283_ (.A(net1537),
    .B(\s0.data_out[26][0] ),
    .X(_0351_));
 sg13g2_o21ai_1 _4284_ (.B1(net1551),
    .Y(_0352_),
    .A1(_3580_),
    .A2(_0351_));
 sg13g2_nor2_1 _4285_ (.A(net1566),
    .B(_3579_),
    .Y(_0353_));
 sg13g2_a22oi_1 _4286_ (.Y(_0113_),
    .B1(_0352_),
    .B2(_0353_),
    .A2(_3419_),
    .A1(net1566));
 sg13g2_and2_1 _4287_ (.A(net1537),
    .B(\s0.data_out[26][1] ),
    .X(_0354_));
 sg13g2_o21ai_1 _4288_ (.B1(net1551),
    .Y(_0355_),
    .A1(_3574_),
    .A2(_0354_));
 sg13g2_nor2_1 _4289_ (.A(net1566),
    .B(net455),
    .Y(_0356_));
 sg13g2_a22oi_1 _4290_ (.Y(_0114_),
    .B1(_0355_),
    .B2(_0356_),
    .A2(_3417_),
    .A1(net1566));
 sg13g2_and2_1 _4291_ (.A(net1538),
    .B(net477),
    .X(_0357_));
 sg13g2_o21ai_1 _4292_ (.B1(net1552),
    .Y(_0358_),
    .A1(_3566_),
    .A2(_0357_));
 sg13g2_nor2_1 _4293_ (.A(net1566),
    .B(_3563_),
    .Y(_0359_));
 sg13g2_a22oi_1 _4294_ (.Y(_0115_),
    .B1(_0358_),
    .B2(_0359_),
    .A2(_3413_),
    .A1(net1566));
 sg13g2_and2_1 _4295_ (.A(net1538),
    .B(\s0.data_out[26][3] ),
    .X(_0360_));
 sg13g2_o21ai_1 _4296_ (.B1(net1551),
    .Y(_0361_),
    .A1(_3592_),
    .A2(_0360_));
 sg13g2_nor2_1 _4297_ (.A(net1565),
    .B(_3589_),
    .Y(_0362_));
 sg13g2_a22oi_1 _4298_ (.Y(_0116_),
    .B1(_0361_),
    .B2(_0362_),
    .A2(_3410_),
    .A1(net1564));
 sg13g2_and2_1 _4299_ (.A(net1536),
    .B(\s0.data_out[26][4] ),
    .X(_0363_));
 sg13g2_o21ai_1 _4300_ (.B1(net1549),
    .Y(_0364_),
    .A1(_3631_),
    .A2(_0363_));
 sg13g2_nor2_1 _4301_ (.A(net1565),
    .B(_3628_),
    .Y(_0365_));
 sg13g2_a22oi_1 _4302_ (.Y(_0117_),
    .B1(_0364_),
    .B2(_0365_),
    .A2(_3408_),
    .A1(net1565));
 sg13g2_and2_1 _4303_ (.A(net1536),
    .B(\s0.data_out[26][5] ),
    .X(_0366_));
 sg13g2_o21ai_1 _4304_ (.B1(net1549),
    .Y(_0367_),
    .A1(_3622_),
    .A2(_0366_));
 sg13g2_nor2_1 _4305_ (.A(net1564),
    .B(_3619_),
    .Y(_0368_));
 sg13g2_a22oi_1 _4306_ (.Y(_0118_),
    .B1(_0367_),
    .B2(_0368_),
    .A2(_3405_),
    .A1(net1564));
 sg13g2_and2_1 _4307_ (.A(net1535),
    .B(\s0.data_out[26][6] ),
    .X(_0369_));
 sg13g2_o21ai_1 _4308_ (.B1(net1550),
    .Y(_0370_),
    .A1(_3610_),
    .A2(_0369_));
 sg13g2_nor2_1 _4309_ (.A(net1564),
    .B(_3607_),
    .Y(_0371_));
 sg13g2_a22oi_1 _4310_ (.Y(_0119_),
    .B1(_0370_),
    .B2(_0371_),
    .A2(_3400_),
    .A1(net1564));
 sg13g2_and2_1 _4311_ (.A(net1535),
    .B(net536),
    .X(_0372_));
 sg13g2_o21ai_1 _4312_ (.B1(net1550),
    .Y(_0373_),
    .A1(_3602_),
    .A2(_0372_));
 sg13g2_nor2_1 _4313_ (.A(net1564),
    .B(_3599_),
    .Y(_0374_));
 sg13g2_a22oi_1 _4314_ (.Y(_0120_),
    .B1(_0373_),
    .B2(_0374_),
    .A2(_3399_),
    .A1(net1564));
 sg13g2_o21ai_1 _4315_ (.B1(net1540),
    .Y(_0375_),
    .A1(net1627),
    .A2(net1523));
 sg13g2_nand2_1 _4316_ (.Y(_0376_),
    .A(net1621),
    .B(net1532));
 sg13g2_a21oi_1 _4317_ (.A1(net1621),
    .A2(net1530),
    .Y(_0377_),
    .B1(_0375_));
 sg13g2_a21oi_1 _4318_ (.A1(net1621),
    .A2(net1547),
    .Y(_0378_),
    .B1(net1536));
 sg13g2_nor2_1 _4319_ (.A(_0377_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_o21ai_1 _4320_ (.B1(_0377_),
    .Y(_0380_),
    .A1(net418),
    .A2(net1530));
 sg13g2_nor2_1 _4321_ (.A(net1523),
    .B(_0375_),
    .Y(_0381_));
 sg13g2_nor2_1 _4322_ (.A(net418),
    .B(net1547),
    .Y(_0382_));
 sg13g2_o21ai_1 _4323_ (.B1(_0380_),
    .Y(_0383_),
    .A1(net1540),
    .A2(_0382_));
 sg13g2_o21ai_1 _4324_ (.B1(net1704),
    .Y(_0384_),
    .A1(_0381_),
    .A2(_0383_));
 sg13g2_a21oi_1 _4325_ (.A1(_3372_),
    .A2(_0379_),
    .Y(_0121_),
    .B1(_0384_));
 sg13g2_nor3_1 _4326_ (.A(net1565),
    .B(_0377_),
    .C(_0378_),
    .Y(_0122_));
 sg13g2_and2_1 _4327_ (.A(net1714),
    .B(net379),
    .X(_0123_));
 sg13g2_nand2_1 _4328_ (.Y(_0385_),
    .A(net1533),
    .B(net731));
 sg13g2_mux2_1 _4329_ (.A0(\s0.data_out[26][2] ),
    .A1(\s0.data_out[25][2] ),
    .S(net1531),
    .X(_0386_));
 sg13g2_nor2b_1 _4330_ (.A(net1525),
    .B_N(net1340),
    .Y(_0387_));
 sg13g2_a21o_1 _4331_ (.A2(_0386_),
    .A1(net1525),
    .B1(_0387_),
    .X(_0388_));
 sg13g2_nand2b_1 _4332_ (.Y(_0389_),
    .B(\s0.data_out[25][2] ),
    .A_N(net1548));
 sg13g2_a21oi_1 _4333_ (.A1(_3564_),
    .A2(_0389_),
    .Y(_0390_),
    .B1(net1542));
 sg13g2_a21oi_1 _4334_ (.A1(net1542),
    .A2(_0388_),
    .Y(_0391_),
    .B1(_0390_));
 sg13g2_or2_1 _4335_ (.X(_0392_),
    .B(_0391_),
    .A(net1684));
 sg13g2_nand2_1 _4336_ (.Y(_0393_),
    .A(net1531),
    .B(net767));
 sg13g2_o21ai_1 _4337_ (.B1(_0393_),
    .Y(_0394_),
    .A1(net1531),
    .A2(_3416_));
 sg13g2_nor2b_1 _4338_ (.A(net1525),
    .B_N(net1344),
    .Y(_0395_));
 sg13g2_a21o_1 _4339_ (.A2(_0394_),
    .A1(net1526),
    .B1(_0395_),
    .X(_0396_));
 sg13g2_nand2b_1 _4340_ (.Y(_0397_),
    .B(\s0.data_out[25][1] ),
    .A_N(net1548));
 sg13g2_a21oi_1 _4341_ (.A1(_3572_),
    .A2(_0397_),
    .Y(_0398_),
    .B1(net1543));
 sg13g2_a21oi_1 _4342_ (.A1(net1542),
    .A2(_0396_),
    .Y(_0399_),
    .B1(_0398_));
 sg13g2_mux2_1 _4343_ (.A0(\s0.data_out[26][0] ),
    .A1(\s0.data_out[25][0] ),
    .S(net1531),
    .X(_0400_));
 sg13g2_nor2b_1 _4344_ (.A(net1525),
    .B_N(net1348),
    .Y(_0401_));
 sg13g2_a21oi_1 _4345_ (.A1(net1525),
    .A2(_0400_),
    .Y(_0402_),
    .B1(_0401_));
 sg13g2_nand2b_1 _4346_ (.Y(_0403_),
    .B(net1543),
    .A_N(_0402_));
 sg13g2_o21ai_1 _4347_ (.B1(_3581_),
    .Y(_0404_),
    .A1(net1548),
    .A2(_3420_));
 sg13g2_nand2b_1 _4348_ (.Y(_0405_),
    .B(_0404_),
    .A_N(net1543));
 sg13g2_a221oi_1 _4349_ (.B2(_0405_),
    .C1(net1700),
    .B1(_0403_),
    .A1(net1690),
    .Y(_0406_),
    .A2(_0399_));
 sg13g2_o21ai_1 _4350_ (.B1(_0392_),
    .Y(_0407_),
    .A1(net1690),
    .A2(_0399_));
 sg13g2_nand2_1 _4351_ (.Y(_0408_),
    .A(net1531),
    .B(net775));
 sg13g2_o21ai_1 _4352_ (.B1(_0408_),
    .Y(_0409_),
    .A1(net1531),
    .A2(_3409_));
 sg13g2_nor2_1 _4353_ (.A(net1525),
    .B(net1160),
    .Y(_0410_));
 sg13g2_a21o_1 _4354_ (.A2(_0409_),
    .A1(net1525),
    .B1(_0410_),
    .X(_0411_));
 sg13g2_nand2b_1 _4355_ (.Y(_0412_),
    .B(net775),
    .A_N(net1548));
 sg13g2_a21oi_1 _4356_ (.A1(_3590_),
    .A2(_0412_),
    .Y(_0413_),
    .B1(net1542));
 sg13g2_a21oi_1 _4357_ (.A1(net1542),
    .A2(_0411_),
    .Y(_0414_),
    .B1(_0413_));
 sg13g2_a22oi_1 _4358_ (.Y(_0415_),
    .B1(_0414_),
    .B2(net1675),
    .A2(_0391_),
    .A1(net1684));
 sg13g2_o21ai_1 _4359_ (.B1(_0415_),
    .Y(_0416_),
    .A1(_0406_),
    .A2(_0407_));
 sg13g2_nand2_1 _4360_ (.Y(_0417_),
    .A(net1532),
    .B(\s0.data_out[25][6] ));
 sg13g2_mux2_1 _4361_ (.A0(\s0.data_out[26][6] ),
    .A1(\s0.data_out[25][6] ),
    .S(net1530),
    .X(_0418_));
 sg13g2_nor2b_1 _4362_ (.A(net1523),
    .B_N(net1325),
    .Y(_0419_));
 sg13g2_a21o_1 _4363_ (.A2(_0418_),
    .A1(net1523),
    .B1(_0419_),
    .X(_0420_));
 sg13g2_nand2b_1 _4364_ (.Y(_0421_),
    .B(\s0.data_out[25][6] ),
    .A_N(net1547));
 sg13g2_a21oi_1 _4365_ (.A1(_3608_),
    .A2(_0421_),
    .Y(_0422_),
    .B1(net1540));
 sg13g2_a21oi_1 _4366_ (.A1(net1540),
    .A2(_0420_),
    .Y(_0423_),
    .B1(_0422_));
 sg13g2_nand2_1 _4367_ (.Y(_0424_),
    .A(net1530),
    .B(net548));
 sg13g2_mux2_1 _4368_ (.A0(\s0.data_out[26][7] ),
    .A1(\s0.data_out[25][7] ),
    .S(net1530),
    .X(_0425_));
 sg13g2_nor2b_1 _4369_ (.A(net1524),
    .B_N(net1320),
    .Y(_0426_));
 sg13g2_a21o_1 _4370_ (.A2(_0425_),
    .A1(net1524),
    .B1(_0426_),
    .X(_0427_));
 sg13g2_nand2b_1 _4371_ (.Y(_0428_),
    .B(\s0.data_out[25][7] ),
    .A_N(net1548));
 sg13g2_a21oi_1 _4372_ (.A1(_3600_),
    .A2(_0428_),
    .Y(_0429_),
    .B1(net1541));
 sg13g2_a21oi_1 _4373_ (.A1(net1541),
    .A2(_0427_),
    .Y(_0430_),
    .B1(_0429_));
 sg13g2_a22oi_1 _4374_ (.Y(_0431_),
    .B1(_0430_),
    .B2(net1637),
    .A2(_0423_),
    .A1(net1646));
 sg13g2_nor2_1 _4375_ (.A(net1646),
    .B(_0423_),
    .Y(_0432_));
 sg13g2_nor2_1 _4376_ (.A(net1637),
    .B(_0430_),
    .Y(_0433_));
 sg13g2_or2_1 _4377_ (.X(_0434_),
    .B(_0430_),
    .A(net1637));
 sg13g2_nand3b_1 _4378_ (.B(_0434_),
    .C(_0431_),
    .Y(_0435_),
    .A_N(_0432_));
 sg13g2_nand2_1 _4379_ (.Y(_0436_),
    .A(net1532),
    .B(\s0.data_out[25][4] ));
 sg13g2_mux2_1 _4380_ (.A0(\s0.data_out[26][4] ),
    .A1(\s0.data_out[25][4] ),
    .S(net1531),
    .X(_0437_));
 sg13g2_nor2b_1 _4381_ (.A(net1526),
    .B_N(net1335),
    .Y(_0438_));
 sg13g2_a21o_1 _4382_ (.A2(_0437_),
    .A1(net1526),
    .B1(_0438_),
    .X(_0439_));
 sg13g2_nand2b_1 _4383_ (.Y(_0440_),
    .B(net438),
    .A_N(net1548));
 sg13g2_a21oi_1 _4384_ (.A1(_3629_),
    .A2(_0440_),
    .Y(_0441_),
    .B1(net1541));
 sg13g2_a21oi_1 _4385_ (.A1(net1541),
    .A2(_0439_),
    .Y(_0442_),
    .B1(_0441_));
 sg13g2_nand2_1 _4386_ (.Y(_0443_),
    .A(net1532),
    .B(\s0.data_out[25][5] ));
 sg13g2_mux2_1 _4387_ (.A0(\s0.data_out[26][5] ),
    .A1(\s0.data_out[25][5] ),
    .S(net1530),
    .X(_0444_));
 sg13g2_nor2b_1 _4388_ (.A(net1523),
    .B_N(net1330),
    .Y(_0445_));
 sg13g2_a21o_1 _4389_ (.A2(_0444_),
    .A1(net1523),
    .B1(_0445_),
    .X(_0446_));
 sg13g2_nand2b_1 _4390_ (.Y(_0447_),
    .B(\s0.data_out[25][5] ),
    .A_N(net1547));
 sg13g2_a21oi_1 _4391_ (.A1(_3620_),
    .A2(_0447_),
    .Y(_0448_),
    .B1(net1540));
 sg13g2_a21oi_1 _4392_ (.A1(net1540),
    .A2(_0446_),
    .Y(_0449_),
    .B1(_0448_));
 sg13g2_a22oi_1 _4393_ (.Y(_0450_),
    .B1(_0449_),
    .B2(net1655),
    .A2(_0442_),
    .A1(net1665));
 sg13g2_inv_1 _4394_ (.Y(_0451_),
    .A(_0450_));
 sg13g2_nor2_1 _4395_ (.A(net1675),
    .B(_0414_),
    .Y(_0452_));
 sg13g2_or2_1 _4396_ (.X(_0453_),
    .B(_0449_),
    .A(net1655));
 sg13g2_o21ai_1 _4397_ (.B1(_0453_),
    .Y(_0454_),
    .A1(net1665),
    .A2(_0442_));
 sg13g2_nor4_1 _4398_ (.A(_0435_),
    .B(_0451_),
    .C(_0452_),
    .D(_0454_),
    .Y(_0455_));
 sg13g2_nor2_1 _4399_ (.A(_0435_),
    .B(_0450_),
    .Y(_0456_));
 sg13g2_o21ai_1 _4400_ (.B1(_0379_),
    .Y(_0457_),
    .A1(_0431_),
    .A2(_0433_));
 sg13g2_a221oi_1 _4401_ (.B2(_0453_),
    .C1(_0457_),
    .B1(_0456_),
    .A1(_0416_),
    .Y(_0458_),
    .A2(_0455_));
 sg13g2_nor3_1 _4402_ (.A(net371),
    .B(net1555),
    .C(_0458_),
    .Y(_0124_));
 sg13g2_nor2_1 _4403_ (.A(net1179),
    .B(_3420_),
    .Y(_0459_));
 sg13g2_o21ai_1 _4404_ (.B1(net1543),
    .Y(_0460_),
    .A1(_0401_),
    .A2(_0459_));
 sg13g2_nand3_1 _4405_ (.B(_0405_),
    .C(_0460_),
    .A(net1707),
    .Y(_0461_));
 sg13g2_o21ai_1 _4406_ (.B1(_0461_),
    .Y(_0462_),
    .A1(net1705),
    .A2(net744));
 sg13g2_inv_1 _4407_ (.Y(_0125_),
    .A(_0462_));
 sg13g2_nor2_1 _4408_ (.A(net1179),
    .B(_3421_),
    .Y(_0463_));
 sg13g2_o21ai_1 _4409_ (.B1(net1543),
    .Y(_0464_),
    .A1(_0395_),
    .A2(_0463_));
 sg13g2_nor2_1 _4410_ (.A(net1577),
    .B(_0398_),
    .Y(_0465_));
 sg13g2_a22oi_1 _4411_ (.Y(_0126_),
    .B1(_0464_),
    .B2(_0465_),
    .A2(_3416_),
    .A1(net1570));
 sg13g2_nor2_1 _4412_ (.A(net1179),
    .B(_3423_),
    .Y(_0466_));
 sg13g2_o21ai_1 _4413_ (.B1(net1542),
    .Y(_0467_),
    .A1(_0387_),
    .A2(_0466_));
 sg13g2_nor2_1 _4414_ (.A(net1566),
    .B(_0390_),
    .Y(_0468_));
 sg13g2_a22oi_1 _4415_ (.Y(_0127_),
    .B1(_0467_),
    .B2(_0468_),
    .A2(_3412_),
    .A1(net1567));
 sg13g2_nor2_1 _4416_ (.A(net1179),
    .B(_3422_),
    .Y(_0469_));
 sg13g2_o21ai_1 _4417_ (.B1(net1542),
    .Y(_0470_),
    .A1(_0410_),
    .A2(_0469_));
 sg13g2_nor2_1 _4418_ (.A(net1565),
    .B(_0413_),
    .Y(_0471_));
 sg13g2_a22oi_1 _4419_ (.Y(_0128_),
    .B1(_0470_),
    .B2(_0471_),
    .A2(_3409_),
    .A1(net1567));
 sg13g2_and2_1 _4420_ (.A(net1524),
    .B(net438),
    .X(_0472_));
 sg13g2_o21ai_1 _4421_ (.B1(net1541),
    .Y(_0473_),
    .A1(_0438_),
    .A2(_0472_));
 sg13g2_nor2_1 _4422_ (.A(net1568),
    .B(_0441_),
    .Y(_0474_));
 sg13g2_a22oi_1 _4423_ (.Y(_0129_),
    .B1(_0473_),
    .B2(_0474_),
    .A2(_3407_),
    .A1(net1568));
 sg13g2_and2_1 _4424_ (.A(net1523),
    .B(\s0.data_out[25][5] ),
    .X(_0475_));
 sg13g2_o21ai_1 _4425_ (.B1(net1540),
    .Y(_0476_),
    .A1(_0445_),
    .A2(_0475_));
 sg13g2_nor2_1 _4426_ (.A(net1565),
    .B(_0448_),
    .Y(_0477_));
 sg13g2_a22oi_1 _4427_ (.Y(_0130_),
    .B1(_0476_),
    .B2(_0477_),
    .A2(_3404_),
    .A1(net1565));
 sg13g2_and2_1 _4428_ (.A(net1523),
    .B(\s0.data_out[25][6] ),
    .X(_0478_));
 sg13g2_o21ai_1 _4429_ (.B1(net1540),
    .Y(_0479_),
    .A1(_0419_),
    .A2(_0478_));
 sg13g2_nand3b_1 _4430_ (.B(_0479_),
    .C(net1704),
    .Y(_0480_),
    .A_N(_0422_));
 sg13g2_o21ai_1 _4431_ (.B1(_0480_),
    .Y(_0481_),
    .A1(net1704),
    .A2(net680));
 sg13g2_inv_1 _4432_ (.Y(_0131_),
    .A(_0481_));
 sg13g2_nor2_1 _4433_ (.A(net1179),
    .B(_3424_),
    .Y(_0482_));
 sg13g2_o21ai_1 _4434_ (.B1(net1541),
    .Y(_0483_),
    .A1(_0426_),
    .A2(_0482_));
 sg13g2_nor2_1 _4435_ (.A(net1568),
    .B(_0429_),
    .Y(_0484_));
 sg13g2_a22oi_1 _4436_ (.Y(_0132_),
    .B1(_0483_),
    .B2(_0484_),
    .A2(_3398_),
    .A1(net1568));
 sg13g2_o21ai_1 _4437_ (.B1(net1528),
    .Y(_0485_),
    .A1(net1627),
    .A2(net1510));
 sg13g2_nor2_1 _4438_ (.A(net1629),
    .B(_3389_),
    .Y(_0486_));
 sg13g2_nor2_1 _4439_ (.A(_0485_),
    .B(_0486_),
    .Y(_0487_));
 sg13g2_a21oi_1 _4440_ (.A1(net1177),
    .A2(_0376_),
    .Y(_0488_),
    .B1(_0487_));
 sg13g2_o21ai_1 _4441_ (.B1(_0487_),
    .Y(_0489_),
    .A1(\s0.was_valid_out[24] [0]),
    .A2(net1518));
 sg13g2_nor2_1 _4442_ (.A(net1510),
    .B(_0485_),
    .Y(_0490_));
 sg13g2_o21ai_1 _4443_ (.B1(net1177),
    .Y(_0491_),
    .A1(\s0.was_valid_out[24] [0]),
    .A2(net1532));
 sg13g2_nand2_1 _4444_ (.Y(_0492_),
    .A(_0489_),
    .B(_0491_));
 sg13g2_o21ai_1 _4445_ (.B1(net1714),
    .Y(_0493_),
    .A1(_0490_),
    .A2(_0492_));
 sg13g2_a21oi_1 _4446_ (.A1(_3371_),
    .A2(_0488_),
    .Y(_0133_),
    .B1(_0493_));
 sg13g2_and2_1 _4447_ (.A(net1706),
    .B(_0488_),
    .X(_0134_));
 sg13g2_and2_1 _4448_ (.A(net1716),
    .B(net382),
    .X(_0135_));
 sg13g2_nand2_1 _4449_ (.Y(_0494_),
    .A(net1518),
    .B(net509));
 sg13g2_o21ai_1 _4450_ (.B1(_0494_),
    .Y(_0495_),
    .A1(net1519),
    .A2(_3421_));
 sg13g2_nor2b_1 _4451_ (.A(net1511),
    .B_N(net1344),
    .Y(_0496_));
 sg13g2_a21o_1 _4452_ (.A2(_0495_),
    .A1(net1511),
    .B1(_0496_),
    .X(_0497_));
 sg13g2_nand2b_1 _4453_ (.Y(_0498_),
    .B(net509),
    .A_N(net1533));
 sg13g2_a21oi_1 _4454_ (.A1(_0393_),
    .A2(_0498_),
    .Y(_0499_),
    .B1(net1528));
 sg13g2_a21oi_1 _4455_ (.A1(net1528),
    .A2(_0497_),
    .Y(_0500_),
    .B1(_0499_));
 sg13g2_mux2_1 _4456_ (.A0(\s0.data_out[24][0] ),
    .A1(net556),
    .S(net1533),
    .X(_0501_));
 sg13g2_nand2_1 _4457_ (.Y(_0502_),
    .A(net1178),
    .B(_0501_));
 sg13g2_nor2b_1 _4458_ (.A(net1511),
    .B_N(net1348),
    .Y(_0503_));
 sg13g2_nand2_1 _4459_ (.Y(_0504_),
    .A(net1518),
    .B(\s0.data_out[24][0] ));
 sg13g2_o21ai_1 _4460_ (.B1(_0504_),
    .Y(_0505_),
    .A1(net1519),
    .A2(_3420_));
 sg13g2_a21oi_1 _4461_ (.A1(net1511),
    .A2(_0505_),
    .Y(_0506_),
    .B1(_0503_));
 sg13g2_nand2b_1 _4462_ (.Y(_0507_),
    .B(net1528),
    .A_N(_0506_));
 sg13g2_a221oi_1 _4463_ (.B2(_0507_),
    .C1(net1700),
    .B1(_0502_),
    .A1(net1692),
    .Y(_0508_),
    .A2(_0500_));
 sg13g2_nor2b_1 _4464_ (.A(net1512),
    .B_N(net1340),
    .Y(_0509_));
 sg13g2_nand2_1 _4465_ (.Y(_0510_),
    .A(net1521),
    .B(net631));
 sg13g2_o21ai_1 _4466_ (.B1(_0510_),
    .Y(_0511_),
    .A1(net1519),
    .A2(_3423_));
 sg13g2_a21oi_1 _4467_ (.A1(net1512),
    .A2(_0511_),
    .Y(_0512_),
    .B1(_0509_));
 sg13g2_o21ai_1 _4468_ (.B1(_0385_),
    .Y(_0513_),
    .A1(net1533),
    .A2(_3430_));
 sg13g2_nand2_1 _4469_ (.Y(_0514_),
    .A(net1178),
    .B(_0513_));
 sg13g2_o21ai_1 _4470_ (.B1(_0514_),
    .Y(_0515_),
    .A1(net1178),
    .A2(_0512_));
 sg13g2_or2_1 _4471_ (.X(_0516_),
    .B(_0515_),
    .A(net1560));
 sg13g2_xnor2_1 _4472_ (.Y(_0517_),
    .A(net1560),
    .B(_0515_));
 sg13g2_nor2_1 _4473_ (.A(net1690),
    .B(_0500_),
    .Y(_0518_));
 sg13g2_nand2_1 _4474_ (.Y(_0519_),
    .A(net1518),
    .B(net502));
 sg13g2_o21ai_1 _4475_ (.B1(_0519_),
    .Y(_0520_),
    .A1(net1519),
    .A2(_3422_));
 sg13g2_nor2_1 _4476_ (.A(net1511),
    .B(net1160),
    .Y(_0521_));
 sg13g2_a21o_1 _4477_ (.A2(_0520_),
    .A1(net1511),
    .B1(_0521_),
    .X(_0522_));
 sg13g2_nand2b_1 _4478_ (.Y(_0523_),
    .B(net502),
    .A_N(net1530));
 sg13g2_a21oi_1 _4479_ (.A1(_0408_),
    .A2(_0523_),
    .Y(_0524_),
    .B1(net1525));
 sg13g2_a21oi_1 _4480_ (.A1(net1528),
    .A2(_0522_),
    .Y(_0525_),
    .B1(_0524_));
 sg13g2_nor2_1 _4481_ (.A(net1676),
    .B(_0525_),
    .Y(_0526_));
 sg13g2_nor4_1 _4482_ (.A(_0508_),
    .B(_0517_),
    .C(_0518_),
    .D(_0526_),
    .Y(_0527_));
 sg13g2_nand2_1 _4483_ (.Y(_0528_),
    .A(net1676),
    .B(_0525_));
 sg13g2_o21ai_1 _4484_ (.B1(_0528_),
    .Y(_0529_),
    .A1(_0516_),
    .A2(_0526_));
 sg13g2_nand2_1 _4485_ (.Y(_0530_),
    .A(net1520),
    .B(net540));
 sg13g2_mux2_1 _4486_ (.A0(\s0.data_out[25][7] ),
    .A1(\s0.data_out[24][7] ),
    .S(net1518),
    .X(_0531_));
 sg13g2_nor2b_1 _4487_ (.A(net1509),
    .B_N(net1320),
    .Y(_0532_));
 sg13g2_a21o_1 _4488_ (.A2(_0531_),
    .A1(net1509),
    .B1(_0532_),
    .X(_0533_));
 sg13g2_nand2b_1 _4489_ (.Y(_0534_),
    .B(net540),
    .A_N(net1530));
 sg13g2_a21oi_1 _4490_ (.A1(_0424_),
    .A2(_0534_),
    .Y(_0535_),
    .B1(net1527));
 sg13g2_a21oi_1 _4491_ (.A1(net1527),
    .A2(_0533_),
    .Y(_0536_),
    .B1(_0535_));
 sg13g2_nand2_1 _4492_ (.Y(_0537_),
    .A(net1520),
    .B(net554));
 sg13g2_mux2_1 _4493_ (.A0(\s0.data_out[25][6] ),
    .A1(\s0.data_out[24][6] ),
    .S(net1518),
    .X(_0538_));
 sg13g2_nor2b_1 _4494_ (.A(net1509),
    .B_N(net1325),
    .Y(_0539_));
 sg13g2_a21o_1 _4495_ (.A2(_0538_),
    .A1(net1509),
    .B1(_0539_),
    .X(_0540_));
 sg13g2_nand2b_1 _4496_ (.Y(_0541_),
    .B(\s0.data_out[24][6] ),
    .A_N(net1532));
 sg13g2_a21oi_1 _4497_ (.A1(_0417_),
    .A2(_0541_),
    .Y(_0542_),
    .B1(net1527));
 sg13g2_a21oi_1 _4498_ (.A1(net1527),
    .A2(_0540_),
    .Y(_0543_),
    .B1(_0542_));
 sg13g2_a22oi_1 _4499_ (.Y(_0544_),
    .B1(_0543_),
    .B2(net1646),
    .A2(_0536_),
    .A1(net1637));
 sg13g2_nor2_1 _4500_ (.A(net1646),
    .B(_0543_),
    .Y(_0545_));
 sg13g2_or2_1 _4501_ (.X(_0546_),
    .B(_0536_),
    .A(net1637));
 sg13g2_inv_1 _4502_ (.Y(_0547_),
    .A(_0546_));
 sg13g2_nand3b_1 _4503_ (.B(_0546_),
    .C(_0544_),
    .Y(_0548_),
    .A_N(_0545_));
 sg13g2_nand2_1 _4504_ (.Y(_0549_),
    .A(net1520),
    .B(net429));
 sg13g2_mux2_1 _4505_ (.A0(\s0.data_out[25][5] ),
    .A1(\s0.data_out[24][5] ),
    .S(net1518),
    .X(_0550_));
 sg13g2_nor2b_1 _4506_ (.A(net1509),
    .B_N(net1330),
    .Y(_0551_));
 sg13g2_a21oi_1 _4507_ (.A1(net1510),
    .A2(_0550_),
    .Y(_0552_),
    .B1(_0551_));
 sg13g2_nand2b_1 _4508_ (.Y(_0553_),
    .B(net1527),
    .A_N(_0552_));
 sg13g2_o21ai_1 _4509_ (.B1(_0443_),
    .Y(_0554_),
    .A1(net1532),
    .A2(_3427_));
 sg13g2_nand2_1 _4510_ (.Y(_0555_),
    .A(net1177),
    .B(_0554_));
 sg13g2_nand3_1 _4511_ (.B(_0553_),
    .C(_0555_),
    .A(net1658),
    .Y(_0556_));
 sg13g2_nor2b_1 _4512_ (.A(net1512),
    .B_N(net1335),
    .Y(_0557_));
 sg13g2_nand2_1 _4513_ (.Y(_0558_),
    .A(net1520),
    .B(net592));
 sg13g2_mux2_1 _4514_ (.A0(\s0.data_out[25][4] ),
    .A1(\s0.data_out[24][4] ),
    .S(net1518),
    .X(_0559_));
 sg13g2_a21oi_1 _4515_ (.A1(net1510),
    .A2(_0559_),
    .Y(_0560_),
    .B1(_0557_));
 sg13g2_nand2b_1 _4516_ (.Y(_0561_),
    .B(net1527),
    .A_N(_0560_));
 sg13g2_o21ai_1 _4517_ (.B1(_0436_),
    .Y(_0562_),
    .A1(net1532),
    .A2(_3428_));
 sg13g2_nand2_1 _4518_ (.Y(_0563_),
    .A(net1177),
    .B(_0562_));
 sg13g2_nand3_1 _4519_ (.B(_0561_),
    .C(_0563_),
    .A(net1667),
    .Y(_0564_));
 sg13g2_nand2_1 _4520_ (.Y(_0565_),
    .A(_0556_),
    .B(_0564_));
 sg13g2_a21oi_1 _4521_ (.A1(_0553_),
    .A2(_0555_),
    .Y(_0566_),
    .B1(net1658));
 sg13g2_inv_1 _4522_ (.Y(_0567_),
    .A(_0566_));
 sg13g2_a21oi_1 _4523_ (.A1(_0561_),
    .A2(_0563_),
    .Y(_0568_),
    .B1(net1667));
 sg13g2_nor4_1 _4524_ (.A(_0548_),
    .B(_0565_),
    .C(_0566_),
    .D(_0568_),
    .Y(_0569_));
 sg13g2_o21ai_1 _4525_ (.B1(_0569_),
    .Y(_0570_),
    .A1(_0527_),
    .A2(_0529_));
 sg13g2_a21oi_1 _4526_ (.A1(_0556_),
    .A2(_0564_),
    .Y(_0571_),
    .B1(_0548_));
 sg13g2_o21ai_1 _4527_ (.B1(_0488_),
    .Y(_0572_),
    .A1(_0544_),
    .A2(_0547_));
 sg13g2_a21oi_1 _4528_ (.A1(_0567_),
    .A2(_0571_),
    .Y(_0573_),
    .B1(_0572_));
 sg13g2_or2_1 _4529_ (.X(_0574_),
    .B(net1555),
    .A(net379));
 sg13g2_a21oi_1 _4530_ (.A1(_0570_),
    .A2(_0573_),
    .Y(_0136_),
    .B1(_0574_));
 sg13g2_and2_1 _4531_ (.A(net1511),
    .B(\s0.data_out[24][0] ),
    .X(_0575_));
 sg13g2_o21ai_1 _4532_ (.B1(net1528),
    .Y(_0576_),
    .A1(_0503_),
    .A2(_0575_));
 sg13g2_a21oi_1 _4533_ (.A1(net1178),
    .A2(_0501_),
    .Y(_0577_),
    .B1(net1569));
 sg13g2_a22oi_1 _4534_ (.Y(_0137_),
    .B1(_0576_),
    .B2(_0577_),
    .A2(_3420_),
    .A1(net1569));
 sg13g2_and2_1 _4535_ (.A(net1512),
    .B(net509),
    .X(_0578_));
 sg13g2_o21ai_1 _4536_ (.B1(net1529),
    .Y(_0579_),
    .A1(_0496_),
    .A2(_0578_));
 sg13g2_nor2_1 _4537_ (.A(net1569),
    .B(_0499_),
    .Y(_0580_));
 sg13g2_a22oi_1 _4538_ (.Y(_0138_),
    .B1(_0579_),
    .B2(_0580_),
    .A2(_3421_),
    .A1(net1569));
 sg13g2_and2_1 _4539_ (.A(net1512),
    .B(\s0.data_out[24][2] ),
    .X(_0581_));
 sg13g2_o21ai_1 _4540_ (.B1(net1529),
    .Y(_0582_),
    .A1(_0509_),
    .A2(_0581_));
 sg13g2_nand3_1 _4541_ (.B(_0514_),
    .C(_0582_),
    .A(net1714),
    .Y(_0583_));
 sg13g2_o21ai_1 _4542_ (.B1(_0583_),
    .Y(_0584_),
    .A1(net1714),
    .A2(net731));
 sg13g2_inv_1 _4543_ (.Y(_0139_),
    .A(net732));
 sg13g2_and2_1 _4544_ (.A(net1511),
    .B(net502),
    .X(_0585_));
 sg13g2_o21ai_1 _4545_ (.B1(net1528),
    .Y(_0586_),
    .A1(_0521_),
    .A2(_0585_));
 sg13g2_nor2_1 _4546_ (.A(net1568),
    .B(_0524_),
    .Y(_0587_));
 sg13g2_a22oi_1 _4547_ (.Y(_0140_),
    .B1(_0586_),
    .B2(_0587_),
    .A2(_3422_),
    .A1(net1568));
 sg13g2_a21oi_1 _4548_ (.A1(net1510),
    .A2(net592),
    .Y(_0588_),
    .B1(_0557_));
 sg13g2_a21oi_1 _4549_ (.A1(net1177),
    .A2(_0562_),
    .Y(_0589_),
    .B1(net1578));
 sg13g2_o21ai_1 _4550_ (.B1(_0589_),
    .Y(_0590_),
    .A1(net1177),
    .A2(_0588_));
 sg13g2_o21ai_1 _4551_ (.B1(_0590_),
    .Y(_0591_),
    .A1(net1714),
    .A2(net438));
 sg13g2_inv_1 _4552_ (.Y(_0141_),
    .A(_0591_));
 sg13g2_a21oi_1 _4553_ (.A1(net1509),
    .A2(net429),
    .Y(_0592_),
    .B1(_0551_));
 sg13g2_a21oi_1 _4554_ (.A1(net1177),
    .A2(_0554_),
    .Y(_0593_),
    .B1(net1578));
 sg13g2_o21ai_1 _4555_ (.B1(_0593_),
    .Y(_0594_),
    .A1(net1177),
    .A2(_0592_));
 sg13g2_o21ai_1 _4556_ (.B1(_0594_),
    .Y(_0595_),
    .A1(net1714),
    .A2(net766));
 sg13g2_inv_1 _4557_ (.Y(_0142_),
    .A(_0595_));
 sg13g2_and2_1 _4558_ (.A(net1509),
    .B(\s0.data_out[24][6] ),
    .X(_0596_));
 sg13g2_o21ai_1 _4559_ (.B1(net1527),
    .Y(_0597_),
    .A1(_0539_),
    .A2(_0596_));
 sg13g2_nand3b_1 _4560_ (.B(_0597_),
    .C(net1706),
    .Y(_0598_),
    .A_N(_0542_));
 sg13g2_o21ai_1 _4561_ (.B1(_0598_),
    .Y(_0599_),
    .A1(net1706),
    .A2(net777));
 sg13g2_inv_1 _4562_ (.Y(_0143_),
    .A(net778));
 sg13g2_and2_1 _4563_ (.A(net1509),
    .B(net540),
    .X(_0600_));
 sg13g2_o21ai_1 _4564_ (.B1(net1527),
    .Y(_0601_),
    .A1(_0532_),
    .A2(_0600_));
 sg13g2_nor2_1 _4565_ (.A(net1568),
    .B(_0535_),
    .Y(_0602_));
 sg13g2_a22oi_1 _4566_ (.Y(_0144_),
    .B1(_0601_),
    .B2(_0602_),
    .A2(_3424_),
    .A1(net1568));
 sg13g2_o21ai_1 _4567_ (.B1(net1513),
    .Y(_0603_),
    .A1(net1629),
    .A2(net1500));
 sg13g2_nand2_1 _4568_ (.Y(_0604_),
    .A(net1622),
    .B(net1506));
 sg13g2_nand2b_1 _4569_ (.Y(_0605_),
    .B(_0604_),
    .A_N(_0603_));
 sg13g2_o21ai_1 _4570_ (.B1(_0605_),
    .Y(_0606_),
    .A1(net1514),
    .A2(_0486_));
 sg13g2_nor2_1 _4571_ (.A(net412),
    .B(net1506),
    .Y(_0607_));
 sg13g2_or2_1 _4572_ (.X(_0608_),
    .B(_0607_),
    .A(_0605_));
 sg13g2_nor2_1 _4573_ (.A(net1500),
    .B(_0603_),
    .Y(_0609_));
 sg13g2_a21oi_1 _4574_ (.A1(_3370_),
    .A2(_3389_),
    .Y(_0610_),
    .B1(net1513));
 sg13g2_nor2_1 _4575_ (.A(_0609_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_o21ai_1 _4576_ (.B1(net1714),
    .Y(_0612_),
    .A1(net697),
    .A2(_0606_));
 sg13g2_a21oi_1 _4577_ (.A1(_0608_),
    .A2(_0611_),
    .Y(_0145_),
    .B1(_0612_));
 sg13g2_nor2_1 _4578_ (.A(net1578),
    .B(_0606_),
    .Y(_0146_));
 sg13g2_and2_1 _4579_ (.A(net1716),
    .B(net378),
    .X(_0147_));
 sg13g2_mux2_1 _4580_ (.A0(\s0.data_out[24][2] ),
    .A1(\s0.data_out[23][2] ),
    .S(net1508),
    .X(_0613_));
 sg13g2_nor2b_1 _4581_ (.A(net1501),
    .B_N(net1341),
    .Y(_0614_));
 sg13g2_a21o_1 _4582_ (.A2(_0613_),
    .A1(net1501),
    .B1(_0614_),
    .X(_0615_));
 sg13g2_nand2b_1 _4583_ (.Y(_0616_),
    .B(\s0.data_out[23][2] ),
    .A_N(net1521));
 sg13g2_a21oi_1 _4584_ (.A1(_0510_),
    .A2(_0616_),
    .Y(_0617_),
    .B1(net1515));
 sg13g2_a21oi_1 _4585_ (.A1(net1515),
    .A2(_0615_),
    .Y(_0618_),
    .B1(_0617_));
 sg13g2_nor2_1 _4586_ (.A(net1685),
    .B(_0618_),
    .Y(_0619_));
 sg13g2_nand2_1 _4587_ (.Y(_0620_),
    .A(net1507),
    .B(net817));
 sg13g2_mux2_1 _4588_ (.A0(\s0.data_out[24][1] ),
    .A1(\s0.data_out[23][1] ),
    .S(net1508),
    .X(_0621_));
 sg13g2_nor2b_1 _4589_ (.A(net1501),
    .B_N(net1345),
    .Y(_0622_));
 sg13g2_a21o_1 _4590_ (.A2(_0621_),
    .A1(net1502),
    .B1(_0622_),
    .X(_0623_));
 sg13g2_nand2b_1 _4591_ (.Y(_0624_),
    .B(\s0.data_out[23][1] ),
    .A_N(net1521));
 sg13g2_a21oi_1 _4592_ (.A1(_0494_),
    .A2(_0624_),
    .Y(_0625_),
    .B1(net1516));
 sg13g2_a21oi_1 _4593_ (.A1(net1515),
    .A2(_0623_),
    .Y(_0626_),
    .B1(_0625_));
 sg13g2_mux2_1 _4594_ (.A0(\s0.data_out[24][0] ),
    .A1(\s0.data_out[23][0] ),
    .S(net1508),
    .X(_0627_));
 sg13g2_nor2b_1 _4595_ (.A(net1501),
    .B_N(net1349),
    .Y(_0628_));
 sg13g2_a21oi_1 _4596_ (.A1(net1501),
    .A2(_0627_),
    .Y(_0629_),
    .B1(_0628_));
 sg13g2_nand2b_1 _4597_ (.Y(_0630_),
    .B(net1515),
    .A_N(_0629_));
 sg13g2_nand2_1 _4598_ (.Y(_0631_),
    .A(_3389_),
    .B(\s0.data_out[23][0] ));
 sg13g2_a21o_1 _4599_ (.A2(_0631_),
    .A1(_0504_),
    .B1(net1515),
    .X(_0632_));
 sg13g2_nor2_1 _4600_ (.A(net1692),
    .B(_0626_),
    .Y(_0633_));
 sg13g2_a221oi_1 _4601_ (.B2(_0632_),
    .C1(net1700),
    .B1(_0630_),
    .A1(net1692),
    .Y(_0634_),
    .A2(_0626_));
 sg13g2_nor3_1 _4602_ (.A(_0619_),
    .B(_0633_),
    .C(_0634_),
    .Y(_0635_));
 sg13g2_nand2_1 _4603_ (.Y(_0636_),
    .A(net1507),
    .B(net802));
 sg13g2_mux2_1 _4604_ (.A0(\s0.data_out[24][3] ),
    .A1(\s0.data_out[23][3] ),
    .S(net1508),
    .X(_0637_));
 sg13g2_nor2b_1 _4605_ (.A(net1501),
    .B_N(net1339),
    .Y(_0638_));
 sg13g2_a21o_1 _4606_ (.A2(_0637_),
    .A1(net1501),
    .B1(_0638_),
    .X(_0639_));
 sg13g2_nand2b_1 _4607_ (.Y(_0640_),
    .B(\s0.data_out[23][3] ),
    .A_N(net1521));
 sg13g2_a21oi_1 _4608_ (.A1(_0519_),
    .A2(_0640_),
    .Y(_0641_),
    .B1(net1516));
 sg13g2_a21oi_1 _4609_ (.A1(net1516),
    .A2(_0639_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_a221oi_1 _4610_ (.B2(net1676),
    .C1(_0635_),
    .B1(_0642_),
    .A1(net1685),
    .Y(_0643_),
    .A2(_0618_));
 sg13g2_nand2_1 _4611_ (.Y(_0644_),
    .A(net1506),
    .B(net727));
 sg13g2_mux2_1 _4612_ (.A0(\s0.data_out[24][7] ),
    .A1(\s0.data_out[23][7] ),
    .S(net1508),
    .X(_0645_));
 sg13g2_nor2b_1 _4613_ (.A(net1499),
    .B_N(net1321),
    .Y(_0646_));
 sg13g2_a21o_1 _4614_ (.A2(_0645_),
    .A1(net1500),
    .B1(_0646_),
    .X(_0647_));
 sg13g2_nand2b_1 _4615_ (.Y(_0648_),
    .B(\s0.data_out[23][7] ),
    .A_N(net1520));
 sg13g2_a21oi_1 _4616_ (.A1(_0530_),
    .A2(_0648_),
    .Y(_0649_),
    .B1(net1513));
 sg13g2_a21oi_1 _4617_ (.A1(net1513),
    .A2(_0647_),
    .Y(_0650_),
    .B1(_0649_));
 sg13g2_nand2_1 _4618_ (.Y(_0651_),
    .A(net1506),
    .B(net570));
 sg13g2_mux2_1 _4619_ (.A0(\s0.data_out[24][6] ),
    .A1(\s0.data_out[23][6] ),
    .S(net1508),
    .X(_0652_));
 sg13g2_nor2b_1 _4620_ (.A(net1499),
    .B_N(net1326),
    .Y(_0653_));
 sg13g2_a21o_1 _4621_ (.A2(_0652_),
    .A1(net1500),
    .B1(_0653_),
    .X(_0654_));
 sg13g2_nand2b_1 _4622_ (.Y(_0655_),
    .B(\s0.data_out[23][6] ),
    .A_N(net1520));
 sg13g2_a21oi_1 _4623_ (.A1(_0537_),
    .A2(_0655_),
    .Y(_0656_),
    .B1(net1513));
 sg13g2_a21oi_1 _4624_ (.A1(net1513),
    .A2(_0654_),
    .Y(_0657_),
    .B1(_0656_));
 sg13g2_a22oi_1 _4625_ (.Y(_0658_),
    .B1(_0657_),
    .B2(net1648),
    .A2(_0650_),
    .A1(net1638));
 sg13g2_or2_1 _4626_ (.X(_0659_),
    .B(_0657_),
    .A(net1648));
 sg13g2_or2_1 _4627_ (.X(_0660_),
    .B(_0650_),
    .A(net1638));
 sg13g2_nand3_1 _4628_ (.B(_0659_),
    .C(_0660_),
    .A(_0658_),
    .Y(_0661_));
 sg13g2_mux2_1 _4629_ (.A0(\s0.data_out[24][4] ),
    .A1(\s0.data_out[23][4] ),
    .S(net1508),
    .X(_0662_));
 sg13g2_nor2b_1 _4630_ (.A(net1499),
    .B_N(net1336),
    .Y(_0663_));
 sg13g2_a21o_1 _4631_ (.A2(_0662_),
    .A1(net1499),
    .B1(_0663_),
    .X(_0664_));
 sg13g2_nand2b_1 _4632_ (.Y(_0665_),
    .B(\s0.data_out[23][4] ),
    .A_N(net1520));
 sg13g2_a21oi_1 _4633_ (.A1(_0558_),
    .A2(_0665_),
    .Y(_0666_),
    .B1(net1514));
 sg13g2_a21oi_1 _4634_ (.A1(net1514),
    .A2(_0664_),
    .Y(_0667_),
    .B1(_0666_));
 sg13g2_mux2_1 _4635_ (.A0(\s0.data_out[24][5] ),
    .A1(\s0.data_out[23][5] ),
    .S(net1508),
    .X(_0668_));
 sg13g2_nor2b_1 _4636_ (.A(net1499),
    .B_N(net1331),
    .Y(_0669_));
 sg13g2_a21o_1 _4637_ (.A2(_0668_),
    .A1(net1499),
    .B1(_0669_),
    .X(_0670_));
 sg13g2_nand2b_1 _4638_ (.Y(_0671_),
    .B(\s0.data_out[23][5] ),
    .A_N(net1520));
 sg13g2_a21oi_1 _4639_ (.A1(_0549_),
    .A2(_0671_),
    .Y(_0672_),
    .B1(net1514));
 sg13g2_a21oi_1 _4640_ (.A1(net1514),
    .A2(_0670_),
    .Y(_0673_),
    .B1(_0672_));
 sg13g2_a22oi_1 _4641_ (.Y(_0674_),
    .B1(_0673_),
    .B2(net1658),
    .A2(_0667_),
    .A1(net1667));
 sg13g2_nor2_1 _4642_ (.A(net1676),
    .B(_0642_),
    .Y(_0675_));
 sg13g2_nor2_1 _4643_ (.A(net1658),
    .B(_0673_),
    .Y(_0676_));
 sg13g2_nor2_1 _4644_ (.A(net1667),
    .B(_0667_),
    .Y(_0677_));
 sg13g2_nor3_1 _4645_ (.A(_0675_),
    .B(_0676_),
    .C(_0677_),
    .Y(_0678_));
 sg13g2_nand2_1 _4646_ (.Y(_0679_),
    .A(_0674_),
    .B(_0678_));
 sg13g2_or3_1 _4647_ (.A(_0643_),
    .B(_0661_),
    .C(_0679_),
    .X(_0680_));
 sg13g2_nor3_1 _4648_ (.A(_0661_),
    .B(_0674_),
    .C(_0676_),
    .Y(_0681_));
 sg13g2_nor2b_1 _4649_ (.A(_0658_),
    .B_N(_0660_),
    .Y(_0682_));
 sg13g2_nor3_1 _4650_ (.A(_0606_),
    .B(_0681_),
    .C(_0682_),
    .Y(_0683_));
 sg13g2_or2_1 _4651_ (.X(_0684_),
    .B(net1556),
    .A(net382));
 sg13g2_a21oi_1 _4652_ (.A1(_0680_),
    .A2(_0683_),
    .Y(_0148_),
    .B1(_0684_));
 sg13g2_and2_1 _4653_ (.A(net1501),
    .B(\s0.data_out[23][0] ),
    .X(_0685_));
 sg13g2_o21ai_1 _4654_ (.B1(net1515),
    .Y(_0686_),
    .A1(_0628_),
    .A2(_0685_));
 sg13g2_nand3_1 _4655_ (.B(_0632_),
    .C(_0686_),
    .A(net1714),
    .Y(_0687_));
 sg13g2_o21ai_1 _4656_ (.B1(_0687_),
    .Y(_0688_),
    .A1(net1715),
    .A2(net677));
 sg13g2_inv_1 _4657_ (.Y(_0149_),
    .A(_0688_));
 sg13g2_nor2_1 _4658_ (.A(net1175),
    .B(_3436_),
    .Y(_0689_));
 sg13g2_o21ai_1 _4659_ (.B1(net1516),
    .Y(_0690_),
    .A1(_0622_),
    .A2(_0689_));
 sg13g2_nor2_1 _4660_ (.A(net1579),
    .B(_0625_),
    .Y(_0691_));
 sg13g2_a22oi_1 _4661_ (.Y(_0150_),
    .B1(_0690_),
    .B2(_0691_),
    .A2(_3431_),
    .A1(net1579));
 sg13g2_nor2_1 _4662_ (.A(net1175),
    .B(_3435_),
    .Y(_0692_));
 sg13g2_o21ai_1 _4663_ (.B1(net1515),
    .Y(_0693_),
    .A1(_0614_),
    .A2(_0692_));
 sg13g2_nor2_1 _4664_ (.A(net1578),
    .B(_0617_),
    .Y(_0694_));
 sg13g2_a22oi_1 _4665_ (.Y(_0151_),
    .B1(_0693_),
    .B2(_0694_),
    .A2(_3430_),
    .A1(net1578));
 sg13g2_nor2_1 _4666_ (.A(net1175),
    .B(_3434_),
    .Y(_0695_));
 sg13g2_o21ai_1 _4667_ (.B1(net1515),
    .Y(_0696_),
    .A1(_0638_),
    .A2(_0695_));
 sg13g2_nor2_1 _4668_ (.A(net1579),
    .B(_0641_),
    .Y(_0697_));
 sg13g2_a22oi_1 _4669_ (.Y(_0152_),
    .B1(_0696_),
    .B2(_0697_),
    .A2(_3429_),
    .A1(net1580));
 sg13g2_and2_1 _4670_ (.A(net1499),
    .B(\s0.data_out[23][4] ),
    .X(_0698_));
 sg13g2_o21ai_1 _4671_ (.B1(net1514),
    .Y(_0699_),
    .A1(_0663_),
    .A2(_0698_));
 sg13g2_nor2_1 _4672_ (.A(net1578),
    .B(_0666_),
    .Y(_0700_));
 sg13g2_a22oi_1 _4673_ (.Y(_0153_),
    .B1(_0699_),
    .B2(_0700_),
    .A2(_3428_),
    .A1(net1578));
 sg13g2_and2_1 _4674_ (.A(net1499),
    .B(net614),
    .X(_0701_));
 sg13g2_o21ai_1 _4675_ (.B1(net1514),
    .Y(_0702_),
    .A1(_0669_),
    .A2(_0701_));
 sg13g2_nor2_1 _4676_ (.A(net1578),
    .B(net430),
    .Y(_0703_));
 sg13g2_a22oi_1 _4677_ (.Y(_0154_),
    .B1(net615),
    .B2(_0703_),
    .A2(_3427_),
    .A1(net1579));
 sg13g2_nor2_1 _4678_ (.A(net1174),
    .B(_3433_),
    .Y(_0704_));
 sg13g2_o21ai_1 _4679_ (.B1(net1513),
    .Y(_0705_),
    .A1(_0653_),
    .A2(_0704_));
 sg13g2_nor2_1 _4680_ (.A(net1580),
    .B(_0656_),
    .Y(_0706_));
 sg13g2_a22oi_1 _4681_ (.Y(_0155_),
    .B1(_0705_),
    .B2(_0706_),
    .A2(_3426_),
    .A1(net1580));
 sg13g2_nor2_1 _4682_ (.A(net1174),
    .B(_3432_),
    .Y(_0707_));
 sg13g2_o21ai_1 _4683_ (.B1(net1513),
    .Y(_0708_),
    .A1(_0646_),
    .A2(_0707_));
 sg13g2_nor2_1 _4684_ (.A(net1580),
    .B(_0649_),
    .Y(_0709_));
 sg13g2_a22oi_1 _4685_ (.Y(_0156_),
    .B1(_0708_),
    .B2(_0709_),
    .A2(_3425_),
    .A1(net1580));
 sg13g2_o21ai_1 _4686_ (.B1(net1503),
    .Y(_0710_),
    .A1(net1629),
    .A2(net1486));
 sg13g2_a21oi_1 _4687_ (.A1(net1622),
    .A2(net1495),
    .Y(_0711_),
    .B1(_0710_));
 sg13g2_a21oi_1 _4688_ (.A1(net1174),
    .A2(_0604_),
    .Y(_0712_),
    .B1(_0711_));
 sg13g2_o21ai_1 _4689_ (.B1(_0711_),
    .Y(_0713_),
    .A1(net411),
    .A2(net1495));
 sg13g2_nor2_1 _4690_ (.A(net1486),
    .B(_0710_),
    .Y(_0714_));
 sg13g2_o21ai_1 _4691_ (.B1(net1174),
    .Y(_0715_),
    .A1(net411),
    .A2(net1506));
 sg13g2_nand2_1 _4692_ (.Y(_0716_),
    .A(_0713_),
    .B(_0715_));
 sg13g2_o21ai_1 _4693_ (.B1(net1716),
    .Y(_0717_),
    .A1(_0714_),
    .A2(_0716_));
 sg13g2_a21oi_1 _4694_ (.A1(_3370_),
    .A2(_0712_),
    .Y(_0157_),
    .B1(_0717_));
 sg13g2_and2_1 _4695_ (.A(net1716),
    .B(_0712_),
    .X(_0158_));
 sg13g2_and2_1 _4696_ (.A(net1722),
    .B(net374),
    .X(_0159_));
 sg13g2_nand2_1 _4697_ (.Y(_0718_),
    .A(net1495),
    .B(net658));
 sg13g2_o21ai_1 _4698_ (.B1(_0718_),
    .Y(_0719_),
    .A1(net1496),
    .A2(_3436_));
 sg13g2_nor2b_1 _4699_ (.A(net1488),
    .B_N(net1347),
    .Y(_0720_));
 sg13g2_a21o_1 _4700_ (.A2(_0719_),
    .A1(net1488),
    .B1(_0720_),
    .X(_0721_));
 sg13g2_nand2b_1 _4701_ (.Y(_0722_),
    .B(net658),
    .A_N(net1507));
 sg13g2_a21oi_1 _4702_ (.A1(_0620_),
    .A2(_0722_),
    .Y(_0723_),
    .B1(net1504));
 sg13g2_a21oi_1 _4703_ (.A1(net1504),
    .A2(_0721_),
    .Y(_0724_),
    .B1(_0723_));
 sg13g2_mux2_1 _4704_ (.A0(\s0.data_out[22][0] ),
    .A1(\s0.data_out[23][0] ),
    .S(net1507),
    .X(_0725_));
 sg13g2_nand2_1 _4705_ (.Y(_0726_),
    .A(net1175),
    .B(_0725_));
 sg13g2_nor2b_1 _4706_ (.A(net1488),
    .B_N(net1351),
    .Y(_0727_));
 sg13g2_mux2_1 _4707_ (.A0(\s0.data_out[23][0] ),
    .A1(\s0.data_out[22][0] ),
    .S(net1496),
    .X(_0728_));
 sg13g2_a21oi_1 _4708_ (.A1(net1488),
    .A2(_0728_),
    .Y(_0729_),
    .B1(_0727_));
 sg13g2_nand2b_1 _4709_ (.Y(_0730_),
    .B(net1504),
    .A_N(_0729_));
 sg13g2_a221oi_1 _4710_ (.B2(_0730_),
    .C1(net1701),
    .B1(_0726_),
    .A1(net1694),
    .Y(_0731_),
    .A2(_0724_));
 sg13g2_nand2_1 _4711_ (.Y(_0732_),
    .A(net1495),
    .B(\s0.data_out[22][2] ));
 sg13g2_o21ai_1 _4712_ (.B1(_0732_),
    .Y(_0733_),
    .A1(net1496),
    .A2(_3435_));
 sg13g2_nor2b_1 _4713_ (.A(net1489),
    .B_N(net1341),
    .Y(_0734_));
 sg13g2_a21oi_1 _4714_ (.A1(net1489),
    .A2(_0733_),
    .Y(_0735_),
    .B1(_0734_));
 sg13g2_mux2_1 _4715_ (.A0(\s0.data_out[22][2] ),
    .A1(\s0.data_out[23][2] ),
    .S(net1507),
    .X(_0736_));
 sg13g2_nand2_1 _4716_ (.Y(_0737_),
    .A(net1176),
    .B(_0736_));
 sg13g2_o21ai_1 _4717_ (.B1(_0737_),
    .Y(_0738_),
    .A1(net1175),
    .A2(_0735_));
 sg13g2_or2_1 _4718_ (.X(_0739_),
    .B(_0738_),
    .A(net1561));
 sg13g2_xnor2_1 _4719_ (.Y(_0740_),
    .A(net1561),
    .B(_0738_));
 sg13g2_nor2_1 _4720_ (.A(net1694),
    .B(_0724_),
    .Y(_0741_));
 sg13g2_nand2_1 _4721_ (.Y(_0742_),
    .A(net1496),
    .B(\s0.data_out[22][3] ));
 sg13g2_o21ai_1 _4722_ (.B1(_0742_),
    .Y(_0743_),
    .A1(net1496),
    .A2(_3434_));
 sg13g2_nor2_1 _4723_ (.A(net1488),
    .B(net1162),
    .Y(_0744_));
 sg13g2_a21o_1 _4724_ (.A2(_0743_),
    .A1(net1488),
    .B1(_0744_),
    .X(_0745_));
 sg13g2_nand2b_1 _4725_ (.Y(_0746_),
    .B(net611),
    .A_N(net1507));
 sg13g2_a21oi_1 _4726_ (.A1(_0636_),
    .A2(_0746_),
    .Y(_0747_),
    .B1(net1505));
 sg13g2_a21oi_1 _4727_ (.A1(net1504),
    .A2(_0745_),
    .Y(_0748_),
    .B1(_0747_));
 sg13g2_nor2_1 _4728_ (.A(net1678),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_nor4_1 _4729_ (.A(_0731_),
    .B(_0740_),
    .C(_0741_),
    .D(_0749_),
    .Y(_0750_));
 sg13g2_nand2_1 _4730_ (.Y(_0751_),
    .A(net1678),
    .B(_0748_));
 sg13g2_o21ai_1 _4731_ (.B1(_0751_),
    .Y(_0752_),
    .A1(_0739_),
    .A2(_0749_));
 sg13g2_nand2_1 _4732_ (.Y(_0753_),
    .A(net1497),
    .B(net526));
 sg13g2_mux2_1 _4733_ (.A0(\s0.data_out[23][7] ),
    .A1(\s0.data_out[22][7] ),
    .S(net1495),
    .X(_0754_));
 sg13g2_nor2b_1 _4734_ (.A(net1486),
    .B_N(net1321),
    .Y(_0755_));
 sg13g2_a21o_1 _4735_ (.A2(_0754_),
    .A1(net1486),
    .B1(_0755_),
    .X(_0756_));
 sg13g2_nand2b_1 _4736_ (.Y(_0757_),
    .B(net526),
    .A_N(net1506));
 sg13g2_a21oi_1 _4737_ (.A1(_0644_),
    .A2(_0757_),
    .Y(_0758_),
    .B1(net1503));
 sg13g2_a21oi_1 _4738_ (.A1(net1503),
    .A2(_0756_),
    .Y(_0759_),
    .B1(_0758_));
 sg13g2_nand2_1 _4739_ (.Y(_0760_),
    .A(net1497),
    .B(net488));
 sg13g2_mux2_1 _4740_ (.A0(\s0.data_out[23][6] ),
    .A1(\s0.data_out[22][6] ),
    .S(net1495),
    .X(_0761_));
 sg13g2_nor2b_1 _4741_ (.A(net1486),
    .B_N(net1326),
    .Y(_0762_));
 sg13g2_a21o_1 _4742_ (.A2(_0761_),
    .A1(net1486),
    .B1(_0762_),
    .X(_0763_));
 sg13g2_nand2b_1 _4743_ (.Y(_0764_),
    .B(net488),
    .A_N(net1506));
 sg13g2_a21oi_1 _4744_ (.A1(_0651_),
    .A2(_0764_),
    .Y(_0765_),
    .B1(net1503));
 sg13g2_a21oi_1 _4745_ (.A1(net1503),
    .A2(_0763_),
    .Y(_0766_),
    .B1(_0765_));
 sg13g2_a22oi_1 _4746_ (.Y(_0767_),
    .B1(_0766_),
    .B2(net1648),
    .A2(_0759_),
    .A1(net1638));
 sg13g2_or2_1 _4747_ (.X(_0768_),
    .B(_0766_),
    .A(net1648));
 sg13g2_nor2_1 _4748_ (.A(net1638),
    .B(_0759_),
    .Y(_0769_));
 sg13g2_nand3b_1 _4749_ (.B(_0767_),
    .C(_0768_),
    .Y(_0770_),
    .A_N(_0769_));
 sg13g2_nand2_1 _4750_ (.Y(_0771_),
    .A(net1497),
    .B(\s0.data_out[22][5] ));
 sg13g2_mux2_1 _4751_ (.A0(\s0.data_out[23][5] ),
    .A1(\s0.data_out[22][5] ),
    .S(net1495),
    .X(_0772_));
 sg13g2_nor2b_1 _4752_ (.A(net1487),
    .B_N(net1331),
    .Y(_0773_));
 sg13g2_a21oi_1 _4753_ (.A1(net1487),
    .A2(_0772_),
    .Y(_0774_),
    .B1(_0773_));
 sg13g2_nand2b_1 _4754_ (.Y(_0775_),
    .B(net1503),
    .A_N(_0774_));
 sg13g2_mux2_1 _4755_ (.A0(\s0.data_out[22][5] ),
    .A1(\s0.data_out[23][5] ),
    .S(net1506),
    .X(_0776_));
 sg13g2_nand2_1 _4756_ (.Y(_0777_),
    .A(net1174),
    .B(_0776_));
 sg13g2_nand3_1 _4757_ (.B(_0775_),
    .C(_0777_),
    .A(net1658),
    .Y(_0778_));
 sg13g2_nor2b_1 _4758_ (.A(net1487),
    .B_N(net1336),
    .Y(_0779_));
 sg13g2_mux2_1 _4759_ (.A0(\s0.data_out[23][4] ),
    .A1(\s0.data_out[22][4] ),
    .S(net1495),
    .X(_0780_));
 sg13g2_a21oi_1 _4760_ (.A1(net1487),
    .A2(_0780_),
    .Y(_0781_),
    .B1(_0779_));
 sg13g2_nand2b_1 _4761_ (.Y(_0782_),
    .B(net1504),
    .A_N(_0781_));
 sg13g2_mux2_1 _4762_ (.A0(\s0.data_out[22][4] ),
    .A1(\s0.data_out[23][4] ),
    .S(net1507),
    .X(_0783_));
 sg13g2_nand2_1 _4763_ (.Y(_0784_),
    .A(net1174),
    .B(_0783_));
 sg13g2_nand3_1 _4764_ (.B(_0782_),
    .C(_0784_),
    .A(net1667),
    .Y(_0785_));
 sg13g2_nand2_1 _4765_ (.Y(_0786_),
    .A(_0778_),
    .B(_0785_));
 sg13g2_a21oi_1 _4766_ (.A1(_0782_),
    .A2(_0784_),
    .Y(_0787_),
    .B1(net1667));
 sg13g2_a21oi_1 _4767_ (.A1(_0775_),
    .A2(_0777_),
    .Y(_0788_),
    .B1(net1658));
 sg13g2_a21o_1 _4768_ (.A2(_0777_),
    .A1(_0775_),
    .B1(net1658),
    .X(_0789_));
 sg13g2_nor4_1 _4769_ (.A(_0770_),
    .B(_0786_),
    .C(_0787_),
    .D(_0788_),
    .Y(_0790_));
 sg13g2_o21ai_1 _4770_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_0750_),
    .A2(_0752_));
 sg13g2_a21oi_1 _4771_ (.A1(_0778_),
    .A2(_0785_),
    .Y(_0792_),
    .B1(_0770_));
 sg13g2_o21ai_1 _4772_ (.B1(_0712_),
    .Y(_0793_),
    .A1(_0767_),
    .A2(_0769_));
 sg13g2_a21oi_1 _4773_ (.A1(_0789_),
    .A2(_0792_),
    .Y(_0794_),
    .B1(_0793_));
 sg13g2_or2_1 _4774_ (.X(_0795_),
    .B(net1556),
    .A(net378));
 sg13g2_a21oi_1 _4775_ (.A1(_0791_),
    .A2(_0794_),
    .Y(_0160_),
    .B1(_0795_));
 sg13g2_a21oi_1 _4776_ (.A1(net1488),
    .A2(\s0.data_out[22][0] ),
    .Y(_0796_),
    .B1(_0727_));
 sg13g2_a21oi_1 _4777_ (.A1(net1175),
    .A2(_0725_),
    .Y(_0797_),
    .B1(net1582));
 sg13g2_o21ai_1 _4778_ (.B1(_0797_),
    .Y(_0798_),
    .A1(net1175),
    .A2(_0796_));
 sg13g2_o21ai_1 _4779_ (.B1(_0798_),
    .Y(_0799_),
    .A1(net1716),
    .A2(net738));
 sg13g2_inv_1 _4780_ (.Y(_0161_),
    .A(net739));
 sg13g2_and2_1 _4781_ (.A(net1489),
    .B(net658),
    .X(_0800_));
 sg13g2_o21ai_1 _4782_ (.B1(net1504),
    .Y(_0801_),
    .A1(_0720_),
    .A2(_0800_));
 sg13g2_nor2_1 _4783_ (.A(net1582),
    .B(_0723_),
    .Y(_0802_));
 sg13g2_a22oi_1 _4784_ (.Y(_0162_),
    .B1(_0801_),
    .B2(_0802_),
    .A2(_3436_),
    .A1(net1582));
 sg13g2_a21oi_1 _4785_ (.A1(net1489),
    .A2(\s0.data_out[22][2] ),
    .Y(_0803_),
    .B1(_0734_));
 sg13g2_a21oi_1 _4786_ (.A1(net1176),
    .A2(_0736_),
    .Y(_0804_),
    .B1(net1580));
 sg13g2_o21ai_1 _4787_ (.B1(_0804_),
    .Y(_0805_),
    .A1(net1175),
    .A2(_0803_));
 sg13g2_o21ai_1 _4788_ (.B1(_0805_),
    .Y(_0806_),
    .A1(net1716),
    .A2(net678));
 sg13g2_inv_1 _4789_ (.Y(_0163_),
    .A(net679));
 sg13g2_and2_1 _4790_ (.A(net1488),
    .B(net611),
    .X(_0807_));
 sg13g2_o21ai_1 _4791_ (.B1(net1505),
    .Y(_0808_),
    .A1(_0744_),
    .A2(_0807_));
 sg13g2_nor2_1 _4792_ (.A(net1582),
    .B(_0747_),
    .Y(_0809_));
 sg13g2_a22oi_1 _4793_ (.Y(_0164_),
    .B1(_0808_),
    .B2(_0809_),
    .A2(_3434_),
    .A1(net1582));
 sg13g2_a21oi_1 _4794_ (.A1(net1487),
    .A2(net415),
    .Y(_0810_),
    .B1(_0779_));
 sg13g2_a21oi_1 _4795_ (.A1(net1174),
    .A2(_0783_),
    .Y(_0811_),
    .B1(net1581));
 sg13g2_o21ai_1 _4796_ (.B1(_0811_),
    .Y(_0812_),
    .A1(net1174),
    .A2(_0810_));
 sg13g2_o21ai_1 _4797_ (.B1(_0812_),
    .Y(_0813_),
    .A1(net1716),
    .A2(net743));
 sg13g2_inv_1 _4798_ (.Y(_0165_),
    .A(_0813_));
 sg13g2_a21oi_1 _4799_ (.A1(net1487),
    .A2(net720),
    .Y(_0814_),
    .B1(_0773_));
 sg13g2_a21oi_1 _4800_ (.A1(net1176),
    .A2(_0776_),
    .Y(_0815_),
    .B1(net1581));
 sg13g2_o21ai_1 _4801_ (.B1(_0815_),
    .Y(_0816_),
    .A1(net1176),
    .A2(_0814_));
 sg13g2_o21ai_1 _4802_ (.B1(_0816_),
    .Y(_0817_),
    .A1(net1716),
    .A2(net614));
 sg13g2_inv_1 _4803_ (.Y(_0166_),
    .A(_0817_));
 sg13g2_and2_1 _4804_ (.A(net1486),
    .B(net488),
    .X(_0818_));
 sg13g2_o21ai_1 _4805_ (.B1(net1503),
    .Y(_0819_),
    .A1(_0762_),
    .A2(_0818_));
 sg13g2_nor2_1 _4806_ (.A(net1581),
    .B(_0765_),
    .Y(_0820_));
 sg13g2_a22oi_1 _4807_ (.Y(_0167_),
    .B1(_0819_),
    .B2(_0820_),
    .A2(_3433_),
    .A1(net1580));
 sg13g2_and2_1 _4808_ (.A(net1486),
    .B(net526),
    .X(_0821_));
 sg13g2_o21ai_1 _4809_ (.B1(net1503),
    .Y(_0822_),
    .A1(_0755_),
    .A2(_0821_));
 sg13g2_nor2_1 _4810_ (.A(net1581),
    .B(_0758_),
    .Y(_0823_));
 sg13g2_a22oi_1 _4811_ (.Y(_0168_),
    .B1(_0822_),
    .B2(_0823_),
    .A2(_3432_),
    .A1(net1580));
 sg13g2_o21ai_1 _4812_ (.B1(net1490),
    .Y(_0824_),
    .A1(net1630),
    .A2(net1474));
 sg13g2_nor2b_1 _4813_ (.A(net1630),
    .B_N(net1483),
    .Y(_0825_));
 sg13g2_nor2_1 _4814_ (.A(_0824_),
    .B(_0825_),
    .Y(_0826_));
 sg13g2_a21oi_1 _4815_ (.A1(net1623),
    .A2(net1497),
    .Y(_0827_),
    .B1(net1490));
 sg13g2_nor2_1 _4816_ (.A(_0826_),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_o21ai_1 _4817_ (.B1(_0826_),
    .Y(_0829_),
    .A1(net400),
    .A2(net1483));
 sg13g2_nor2_1 _4818_ (.A(net1474),
    .B(_0824_),
    .Y(_0830_));
 sg13g2_nor2_1 _4819_ (.A(net400),
    .B(net1497),
    .Y(_0831_));
 sg13g2_o21ai_1 _4820_ (.B1(_0829_),
    .Y(_0832_),
    .A1(net1490),
    .A2(_0831_));
 sg13g2_o21ai_1 _4821_ (.B1(net1722),
    .Y(_0833_),
    .A1(_0830_),
    .A2(_0832_));
 sg13g2_a21oi_1 _4822_ (.A1(_3369_),
    .A2(_0828_),
    .Y(_0169_),
    .B1(_0833_));
 sg13g2_nor3_1 _4823_ (.A(net1592),
    .B(_0826_),
    .C(_0827_),
    .Y(_0170_));
 sg13g2_and2_1 _4824_ (.A(net1724),
    .B(net387),
    .X(_0171_));
 sg13g2_nand2_1 _4825_ (.Y(_0834_),
    .A(net1484),
    .B(\s0.data_out[21][2] ));
 sg13g2_mux2_1 _4826_ (.A0(\s0.data_out[22][2] ),
    .A1(\s0.data_out[21][2] ),
    .S(net1484),
    .X(_0835_));
 sg13g2_nor2b_1 _4827_ (.A(net1478),
    .B_N(net1343),
    .Y(_0836_));
 sg13g2_a21oi_1 _4828_ (.A1(net1478),
    .A2(_0835_),
    .Y(_0837_),
    .B1(_0836_));
 sg13g2_nand2b_1 _4829_ (.Y(_0838_),
    .B(net1492),
    .A_N(_0837_));
 sg13g2_o21ai_1 _4830_ (.B1(_0732_),
    .Y(_0839_),
    .A1(net1498),
    .A2(_3444_));
 sg13g2_nand2b_1 _4831_ (.Y(_0840_),
    .B(_0839_),
    .A_N(net1492));
 sg13g2_and2_1 _4832_ (.A(_0838_),
    .B(_0840_),
    .X(_0841_));
 sg13g2_a21o_1 _4833_ (.A2(_0840_),
    .A1(_0838_),
    .B1(net1688),
    .X(_0842_));
 sg13g2_nand2_1 _4834_ (.Y(_0843_),
    .A(net1484),
    .B(\s0.data_out[21][1] ));
 sg13g2_o21ai_1 _4835_ (.B1(_0843_),
    .Y(_0844_),
    .A1(net1484),
    .A2(_3440_));
 sg13g2_nor2b_1 _4836_ (.A(net1478),
    .B_N(net1347),
    .Y(_0845_));
 sg13g2_a21o_1 _4837_ (.A2(_0844_),
    .A1(net1479),
    .B1(_0845_),
    .X(_0846_));
 sg13g2_nand2b_1 _4838_ (.Y(_0847_),
    .B(net551),
    .A_N(net1498));
 sg13g2_a21oi_1 _4839_ (.A1(_0718_),
    .A2(_0847_),
    .Y(_0848_),
    .B1(net1492));
 sg13g2_a21oi_1 _4840_ (.A1(net1492),
    .A2(_0846_),
    .Y(_0849_),
    .B1(_0848_));
 sg13g2_mux2_1 _4841_ (.A0(\s0.data_out[22][0] ),
    .A1(\s0.data_out[21][0] ),
    .S(net1484),
    .X(_0850_));
 sg13g2_nor2b_1 _4842_ (.A(net1478),
    .B_N(net1351),
    .Y(_0851_));
 sg13g2_a21oi_1 _4843_ (.A1(net1478),
    .A2(_0850_),
    .Y(_0852_),
    .B1(_0851_));
 sg13g2_nand2b_1 _4844_ (.Y(_0853_),
    .B(net1492),
    .A_N(_0852_));
 sg13g2_mux2_1 _4845_ (.A0(\s0.data_out[21][0] ),
    .A1(\s0.data_out[22][0] ),
    .S(net1498),
    .X(_0854_));
 sg13g2_nand2b_1 _4846_ (.Y(_0855_),
    .B(_0854_),
    .A_N(net1493));
 sg13g2_a221oi_1 _4847_ (.B2(_0855_),
    .C1(net1701),
    .B1(_0853_),
    .A1(net1694),
    .Y(_0856_),
    .A2(_0849_));
 sg13g2_o21ai_1 _4848_ (.B1(_0842_),
    .Y(_0857_),
    .A1(net1694),
    .A2(_0849_));
 sg13g2_nor2_1 _4849_ (.A(net1478),
    .B(net1161),
    .Y(_0858_));
 sg13g2_nand2_1 _4850_ (.Y(_0859_),
    .A(net1484),
    .B(net499));
 sg13g2_o21ai_1 _4851_ (.B1(_0859_),
    .Y(_0860_),
    .A1(net1484),
    .A2(_3439_));
 sg13g2_a21o_1 _4852_ (.A2(_0860_),
    .A1(net1478),
    .B1(_0858_),
    .X(_0861_));
 sg13g2_nand2b_1 _4853_ (.Y(_0862_),
    .B(\s0.data_out[21][3] ),
    .A_N(net1498));
 sg13g2_a21oi_1 _4854_ (.A1(_0742_),
    .A2(_0862_),
    .Y(_0863_),
    .B1(net1494));
 sg13g2_a21oi_1 _4855_ (.A1(net1492),
    .A2(_0861_),
    .Y(_0864_),
    .B1(_0863_));
 sg13g2_a22oi_1 _4856_ (.Y(_0865_),
    .B1(_0864_),
    .B2(net1678),
    .A2(_0841_),
    .A1(net1688));
 sg13g2_o21ai_1 _4857_ (.B1(_0865_),
    .Y(_0866_),
    .A1(_0856_),
    .A2(_0857_));
 sg13g2_nand2_1 _4858_ (.Y(_0867_),
    .A(net1482),
    .B(net544));
 sg13g2_mux2_1 _4859_ (.A0(\s0.data_out[22][7] ),
    .A1(\s0.data_out[21][7] ),
    .S(net1483),
    .X(_0868_));
 sg13g2_nor2b_1 _4860_ (.A(net1474),
    .B_N(net1322),
    .Y(_0869_));
 sg13g2_a21o_1 _4861_ (.A2(_0868_),
    .A1(net1474),
    .B1(_0869_),
    .X(_0870_));
 sg13g2_nand2b_1 _4862_ (.Y(_0871_),
    .B(\s0.data_out[21][7] ),
    .A_N(net1497));
 sg13g2_a21oi_1 _4863_ (.A1(_0753_),
    .A2(_0871_),
    .Y(_0872_),
    .B1(net1490));
 sg13g2_a21oi_1 _4864_ (.A1(net1490),
    .A2(_0870_),
    .Y(_0873_),
    .B1(_0872_));
 sg13g2_nand2_1 _4865_ (.Y(_0874_),
    .A(net1482),
    .B(net715));
 sg13g2_mux2_1 _4866_ (.A0(\s0.data_out[22][6] ),
    .A1(\s0.data_out[21][6] ),
    .S(net1483),
    .X(_0875_));
 sg13g2_nor2b_1 _4867_ (.A(net1474),
    .B_N(net1327),
    .Y(_0876_));
 sg13g2_a21o_1 _4868_ (.A2(_0875_),
    .A1(net1474),
    .B1(_0876_),
    .X(_0877_));
 sg13g2_nand2b_1 _4869_ (.Y(_0878_),
    .B(\s0.data_out[21][6] ),
    .A_N(net1497));
 sg13g2_a21oi_1 _4870_ (.A1(_0760_),
    .A2(_0878_),
    .Y(_0879_),
    .B1(net1491));
 sg13g2_a21oi_1 _4871_ (.A1(net1491),
    .A2(_0877_),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_a22oi_1 _4872_ (.Y(_0881_),
    .B1(_0880_),
    .B2(net1651),
    .A2(_0873_),
    .A1(net1641));
 sg13g2_inv_1 _4873_ (.Y(_0882_),
    .A(_0881_));
 sg13g2_nor2_1 _4874_ (.A(net1651),
    .B(_0880_),
    .Y(_0883_));
 sg13g2_nor2_1 _4875_ (.A(net1641),
    .B(_0873_),
    .Y(_0884_));
 sg13g2_nor3_1 _4876_ (.A(_0882_),
    .B(_0883_),
    .C(_0884_),
    .Y(_0885_));
 sg13g2_nand2_1 _4877_ (.Y(_0886_),
    .A(net1482),
    .B(net449));
 sg13g2_mux2_1 _4878_ (.A0(\s0.data_out[22][5] ),
    .A1(\s0.data_out[21][5] ),
    .S(net1483),
    .X(_0887_));
 sg13g2_nor2b_1 _4879_ (.A(net1474),
    .B_N(net1332),
    .Y(_0888_));
 sg13g2_a21oi_1 _4880_ (.A1(net1477),
    .A2(_0887_),
    .Y(_0889_),
    .B1(_0888_));
 sg13g2_nand2b_1 _4881_ (.Y(_0890_),
    .B(net1490),
    .A_N(_0889_));
 sg13g2_o21ai_1 _4882_ (.B1(_0771_),
    .Y(_0891_),
    .A1(net1498),
    .A2(_3442_));
 sg13g2_nand2b_1 _4883_ (.Y(_0892_),
    .B(_0891_),
    .A_N(net1491));
 sg13g2_nand3_1 _4884_ (.B(_0890_),
    .C(_0892_),
    .A(net1660),
    .Y(_0893_));
 sg13g2_nor2b_1 _4885_ (.A(net1480),
    .B_N(net1338),
    .Y(_0894_));
 sg13g2_nand2_1 _4886_ (.Y(_0895_),
    .A(net1483),
    .B(\s0.data_out[21][4] ));
 sg13g2_mux2_1 _4887_ (.A0(\s0.data_out[22][4] ),
    .A1(\s0.data_out[21][4] ),
    .S(net1483),
    .X(_0896_));
 sg13g2_a21oi_1 _4888_ (.A1(net1480),
    .A2(_0896_),
    .Y(_0897_),
    .B1(_0894_));
 sg13g2_nand2b_1 _4889_ (.Y(_0898_),
    .B(net1490),
    .A_N(_0897_));
 sg13g2_mux2_1 _4890_ (.A0(\s0.data_out[21][4] ),
    .A1(\s0.data_out[22][4] ),
    .S(net1497),
    .X(_0899_));
 sg13g2_nand2b_1 _4891_ (.Y(_0900_),
    .B(_0899_),
    .A_N(net1491));
 sg13g2_nand3_1 _4892_ (.B(_0898_),
    .C(_0900_),
    .A(net1670),
    .Y(_0901_));
 sg13g2_nand2_1 _4893_ (.Y(_0902_),
    .A(_0893_),
    .B(_0901_));
 sg13g2_a21oi_1 _4894_ (.A1(_0898_),
    .A2(_0900_),
    .Y(_0903_),
    .B1(net1670));
 sg13g2_a21oi_1 _4895_ (.A1(_0890_),
    .A2(_0892_),
    .Y(_0904_),
    .B1(net1660));
 sg13g2_nor2_1 _4896_ (.A(net1678),
    .B(_0864_),
    .Y(_0905_));
 sg13g2_nor4_1 _4897_ (.A(_0902_),
    .B(_0903_),
    .C(_0904_),
    .D(_0905_),
    .Y(_0906_));
 sg13g2_nand3_1 _4898_ (.B(_0885_),
    .C(_0906_),
    .A(_0866_),
    .Y(_0907_));
 sg13g2_o21ai_1 _4899_ (.B1(_0893_),
    .Y(_0908_),
    .A1(_0901_),
    .A2(_0904_));
 sg13g2_o21ai_1 _4900_ (.B1(_0828_),
    .Y(_0909_),
    .A1(_0881_),
    .A2(_0884_));
 sg13g2_a21oi_1 _4901_ (.A1(_0885_),
    .A2(_0908_),
    .Y(_0910_),
    .B1(_0909_));
 sg13g2_or2_1 _4902_ (.X(_0911_),
    .B(net1558),
    .A(net374));
 sg13g2_a21oi_1 _4903_ (.A1(_0907_),
    .A2(_0910_),
    .Y(_0172_),
    .B1(_0911_));
 sg13g2_and2_1 _4904_ (.A(net1478),
    .B(\s0.data_out[21][0] ),
    .X(_0912_));
 sg13g2_o21ai_1 _4905_ (.B1(net1493),
    .Y(_0913_),
    .A1(_0851_),
    .A2(_0912_));
 sg13g2_nand3_1 _4906_ (.B(_0855_),
    .C(_0913_),
    .A(net1723),
    .Y(_0914_));
 sg13g2_o21ai_1 _4907_ (.B1(_0914_),
    .Y(_0915_),
    .A1(net1723),
    .A2(net754));
 sg13g2_inv_1 _4908_ (.Y(_0173_),
    .A(_0915_));
 sg13g2_and2_1 _4909_ (.A(net1479),
    .B(net551),
    .X(_0916_));
 sg13g2_o21ai_1 _4910_ (.B1(net1492),
    .Y(_0917_),
    .A1(_0845_),
    .A2(_0916_));
 sg13g2_nor2_1 _4911_ (.A(net1593),
    .B(_0848_),
    .Y(_0918_));
 sg13g2_a22oi_1 _4912_ (.Y(_0174_),
    .B1(_0917_),
    .B2(_0918_),
    .A2(_3440_),
    .A1(net1593));
 sg13g2_nor2_1 _4913_ (.A(net1172),
    .B(_3444_),
    .Y(_0919_));
 sg13g2_o21ai_1 _4914_ (.B1(net1493),
    .Y(_0920_),
    .A1(_0836_),
    .A2(_0919_));
 sg13g2_nand3_1 _4915_ (.B(_0840_),
    .C(_0920_),
    .A(net1723),
    .Y(_0921_));
 sg13g2_o21ai_1 _4916_ (.B1(_0921_),
    .Y(_0922_),
    .A1(net1723),
    .A2(net690));
 sg13g2_inv_1 _4917_ (.Y(_0175_),
    .A(_0922_));
 sg13g2_nor2_1 _4918_ (.A(net1172),
    .B(_3443_),
    .Y(_0923_));
 sg13g2_o21ai_1 _4919_ (.B1(net1492),
    .Y(_0924_),
    .A1(_0858_),
    .A2(_0923_));
 sg13g2_nor2_1 _4920_ (.A(net1593),
    .B(net414),
    .Y(_0925_));
 sg13g2_a22oi_1 _4921_ (.Y(_0176_),
    .B1(_0924_),
    .B2(_0925_),
    .A2(_3439_),
    .A1(net1593));
 sg13g2_and2_1 _4922_ (.A(net1477),
    .B(\s0.data_out[21][4] ),
    .X(_0926_));
 sg13g2_o21ai_1 _4923_ (.B1(net1493),
    .Y(_0927_),
    .A1(_0894_),
    .A2(_0926_));
 sg13g2_nand3_1 _4924_ (.B(_0900_),
    .C(_0927_),
    .A(net1722),
    .Y(_0928_));
 sg13g2_o21ai_1 _4925_ (.B1(_0928_),
    .Y(_0929_),
    .A1(net1722),
    .A2(net415));
 sg13g2_inv_1 _4926_ (.Y(_0177_),
    .A(_0929_));
 sg13g2_nor2_1 _4927_ (.A(net1173),
    .B(_3442_),
    .Y(_0930_));
 sg13g2_o21ai_1 _4928_ (.B1(net1491),
    .Y(_0931_),
    .A1(_0888_),
    .A2(_0930_));
 sg13g2_nand3_1 _4929_ (.B(_0892_),
    .C(_0931_),
    .A(net1722),
    .Y(_0932_));
 sg13g2_o21ai_1 _4930_ (.B1(_0932_),
    .Y(_0933_),
    .A1(net1722),
    .A2(net720));
 sg13g2_inv_1 _4931_ (.Y(_0178_),
    .A(_0933_));
 sg13g2_and2_1 _4932_ (.A(net1474),
    .B(\s0.data_out[21][6] ),
    .X(_0934_));
 sg13g2_o21ai_1 _4933_ (.B1(net1491),
    .Y(_0935_),
    .A1(_0876_),
    .A2(_0934_));
 sg13g2_nor2_1 _4934_ (.A(net1592),
    .B(_0879_),
    .Y(_0936_));
 sg13g2_a22oi_1 _4935_ (.Y(_0179_),
    .B1(_0935_),
    .B2(_0936_),
    .A2(_3438_),
    .A1(net1592));
 sg13g2_nor2_1 _4936_ (.A(net1173),
    .B(_3441_),
    .Y(_0937_));
 sg13g2_o21ai_1 _4937_ (.B1(net1490),
    .Y(_0938_),
    .A1(_0869_),
    .A2(_0937_));
 sg13g2_nor2_1 _4938_ (.A(net1592),
    .B(_0872_),
    .Y(_0939_));
 sg13g2_a22oi_1 _4939_ (.Y(_0180_),
    .B1(_0938_),
    .B2(_0939_),
    .A2(_3437_),
    .A1(net1593));
 sg13g2_o21ai_1 _4940_ (.B1(net1475),
    .Y(_0940_),
    .A1(net1630),
    .A2(net1461));
 sg13g2_nor2_1 _4941_ (.A(net1630),
    .B(_3392_),
    .Y(_0941_));
 sg13g2_nor2_2 _4942_ (.A(_0940_),
    .B(_0941_),
    .Y(_0942_));
 sg13g2_nor2_1 _4943_ (.A(net1475),
    .B(_0825_),
    .Y(_0943_));
 sg13g2_nor2_1 _4944_ (.A(_0942_),
    .B(_0943_),
    .Y(_0944_));
 sg13g2_o21ai_1 _4945_ (.B1(_0942_),
    .Y(_0945_),
    .A1(\s0.was_valid_out[20] [0]),
    .A2(net1470));
 sg13g2_nor2_1 _4946_ (.A(net1461),
    .B(_0940_),
    .Y(_0946_));
 sg13g2_o21ai_1 _4947_ (.B1(net1173),
    .Y(_0947_),
    .A1(\s0.was_valid_out[20] [0]),
    .A2(net1482));
 sg13g2_nand2_1 _4948_ (.Y(_0948_),
    .A(_0945_),
    .B(_0947_));
 sg13g2_o21ai_1 _4949_ (.B1(net1724),
    .Y(_0949_),
    .A1(_0946_),
    .A2(_0948_));
 sg13g2_a21oi_1 _4950_ (.A1(_3368_),
    .A2(_0944_),
    .Y(_0181_),
    .B1(_0949_));
 sg13g2_nor3_1 _4951_ (.A(net1594),
    .B(_0942_),
    .C(_0943_),
    .Y(_0182_));
 sg13g2_nand2_1 _4952_ (.Y(_0950_),
    .A(net1470),
    .B(net691));
 sg13g2_o21ai_1 _4953_ (.B1(_0950_),
    .Y(_0951_),
    .A1(net1470),
    .A2(_3444_));
 sg13g2_nor2b_1 _4954_ (.A(net1463),
    .B_N(net1343),
    .Y(_0952_));
 sg13g2_a21oi_1 _4955_ (.A1(net1463),
    .A2(_0951_),
    .Y(_0953_),
    .B1(_0952_));
 sg13g2_o21ai_1 _4956_ (.B1(_0834_),
    .Y(_0954_),
    .A1(net1484),
    .A2(_3449_));
 sg13g2_nand2_1 _4957_ (.Y(_0955_),
    .A(net1171),
    .B(_0954_));
 sg13g2_o21ai_1 _4958_ (.B1(_0955_),
    .Y(_0956_),
    .A1(net1171),
    .A2(_0953_));
 sg13g2_nor2b_1 _4959_ (.A(net1463),
    .B_N(net1346),
    .Y(_0957_));
 sg13g2_nand2_1 _4960_ (.Y(_0958_),
    .A(net1472),
    .B(net560));
 sg13g2_mux2_1 _4961_ (.A0(\s0.data_out[21][1] ),
    .A1(\s0.data_out[20][1] ),
    .S(net1471),
    .X(_0959_));
 sg13g2_a21oi_1 _4962_ (.A1(net1463),
    .A2(_0959_),
    .Y(_0960_),
    .B1(_0957_));
 sg13g2_nand2b_1 _4963_ (.Y(_0961_),
    .B(net1481),
    .A_N(_0960_));
 sg13g2_o21ai_1 _4964_ (.B1(_0843_),
    .Y(_0962_),
    .A1(net1485),
    .A2(_3450_));
 sg13g2_nand2_1 _4965_ (.Y(_0963_),
    .A(net1171),
    .B(_0962_));
 sg13g2_nand3_1 _4966_ (.B(_0961_),
    .C(_0963_),
    .A(net1695),
    .Y(_0964_));
 sg13g2_a21oi_1 _4967_ (.A1(_0961_),
    .A2(_0963_),
    .Y(_0965_),
    .B1(net1695));
 sg13g2_mux2_1 _4968_ (.A0(\s0.data_out[21][0] ),
    .A1(\s0.data_out[20][0] ),
    .S(net1471),
    .X(_0966_));
 sg13g2_nor2b_1 _4969_ (.A(net1464),
    .B_N(net1350),
    .Y(_0967_));
 sg13g2_a21oi_1 _4970_ (.A1(net1463),
    .A2(_0966_),
    .Y(_0968_),
    .B1(_0967_));
 sg13g2_mux2_1 _4971_ (.A0(\s0.data_out[20][0] ),
    .A1(\s0.data_out[21][0] ),
    .S(net1485),
    .X(_0969_));
 sg13g2_nand2_1 _4972_ (.Y(_0970_),
    .A(net1172),
    .B(_0969_));
 sg13g2_o21ai_1 _4973_ (.B1(_0970_),
    .Y(_0971_),
    .A1(net1172),
    .A2(_0968_));
 sg13g2_and2_1 _4974_ (.A(net1559),
    .B(_0971_),
    .X(_0972_));
 sg13g2_a221oi_1 _4975_ (.B2(_0972_),
    .C1(_0965_),
    .B1(_0964_),
    .A1(net1562),
    .Y(_0973_),
    .A2(_0956_));
 sg13g2_nand2_1 _4976_ (.Y(_0974_),
    .A(net1473),
    .B(net644));
 sg13g2_mux2_1 _4977_ (.A0(\s0.data_out[21][3] ),
    .A1(\s0.data_out[20][3] ),
    .S(net1471),
    .X(_0975_));
 sg13g2_nor2b_1 _4978_ (.A(net1464),
    .B_N(net1339),
    .Y(_0976_));
 sg13g2_a21o_1 _4979_ (.A2(_0975_),
    .A1(net1464),
    .B1(_0976_),
    .X(_0977_));
 sg13g2_nand2b_1 _4980_ (.Y(_0978_),
    .B(\s0.data_out[20][3] ),
    .A_N(net1485));
 sg13g2_a21oi_1 _4981_ (.A1(_0859_),
    .A2(_0978_),
    .Y(_0979_),
    .B1(net1479));
 sg13g2_a21oi_1 _4982_ (.A1(net1481),
    .A2(_0977_),
    .Y(_0980_),
    .B1(_0979_));
 sg13g2_nand2_1 _4983_ (.Y(_0981_),
    .A(net1678),
    .B(_0980_));
 sg13g2_o21ai_1 _4984_ (.B1(_0981_),
    .Y(_0982_),
    .A1(net1562),
    .A2(_0956_));
 sg13g2_nor2_1 _4985_ (.A(_0973_),
    .B(_0982_),
    .Y(_0983_));
 sg13g2_nand2_1 _4986_ (.Y(_0984_),
    .A(net1472),
    .B(net694));
 sg13g2_mux2_1 _4987_ (.A0(\s0.data_out[21][7] ),
    .A1(\s0.data_out[20][7] ),
    .S(net1470),
    .X(_0985_));
 sg13g2_nor2b_1 _4988_ (.A(net1462),
    .B_N(net1322),
    .Y(_0986_));
 sg13g2_a21o_1 _4989_ (.A2(_0985_),
    .A1(net1462),
    .B1(_0986_),
    .X(_0987_));
 sg13g2_nand2b_1 _4990_ (.Y(_0988_),
    .B(\s0.data_out[20][7] ),
    .A_N(net1482));
 sg13g2_a21oi_1 _4991_ (.A1(_0867_),
    .A2(_0988_),
    .Y(_0989_),
    .B1(net1475));
 sg13g2_a21oi_1 _4992_ (.A1(net1475),
    .A2(_0987_),
    .Y(_0990_),
    .B1(_0989_));
 sg13g2_nand2_1 _4993_ (.Y(_0991_),
    .A(net1472),
    .B(net781));
 sg13g2_mux2_1 _4994_ (.A0(\s0.data_out[21][6] ),
    .A1(\s0.data_out[20][6] ),
    .S(net1470),
    .X(_0992_));
 sg13g2_nor2b_1 _4995_ (.A(net1461),
    .B_N(net1327),
    .Y(_0993_));
 sg13g2_a21o_1 _4996_ (.A2(_0992_),
    .A1(net1461),
    .B1(_0993_),
    .X(_0994_));
 sg13g2_nand2b_1 _4997_ (.Y(_0995_),
    .B(net835),
    .A_N(net1482));
 sg13g2_a21oi_1 _4998_ (.A1(_0874_),
    .A2(_0995_),
    .Y(_0996_),
    .B1(net1475));
 sg13g2_a21oi_1 _4999_ (.A1(net1475),
    .A2(_0994_),
    .Y(_0997_),
    .B1(_0996_));
 sg13g2_a22oi_1 _5000_ (.Y(_0998_),
    .B1(_0997_),
    .B2(net1651),
    .A2(_0990_),
    .A1(net1641));
 sg13g2_nor2_1 _5001_ (.A(net1651),
    .B(_0997_),
    .Y(_0999_));
 sg13g2_or2_1 _5002_ (.X(_1000_),
    .B(_0990_),
    .A(net1641));
 sg13g2_nand3b_1 _5003_ (.B(_1000_),
    .C(_0998_),
    .Y(_1001_),
    .A_N(_0999_));
 sg13g2_nand2_1 _5004_ (.Y(_1002_),
    .A(net1470),
    .B(net492));
 sg13g2_mux2_1 _5005_ (.A0(\s0.data_out[21][5] ),
    .A1(\s0.data_out[20][5] ),
    .S(net1470),
    .X(_1003_));
 sg13g2_nor2b_1 _5006_ (.A(net1462),
    .B_N(net1332),
    .Y(_1004_));
 sg13g2_a21o_1 _5007_ (.A2(_1003_),
    .A1(net1462),
    .B1(_1004_),
    .X(_1005_));
 sg13g2_nand2b_1 _5008_ (.Y(_1006_),
    .B(\s0.data_out[20][5] ),
    .A_N(net1482));
 sg13g2_a21oi_1 _5009_ (.A1(_0886_),
    .A2(_1006_),
    .Y(_1007_),
    .B1(net1476));
 sg13g2_a21oi_1 _5010_ (.A1(net1476),
    .A2(_1005_),
    .Y(_1008_),
    .B1(_1007_));
 sg13g2_nand2_1 _5011_ (.Y(_1009_),
    .A(net1660),
    .B(_1008_));
 sg13g2_nand2_1 _5012_ (.Y(_1010_),
    .A(net1472),
    .B(net516));
 sg13g2_mux2_1 _5013_ (.A0(\s0.data_out[21][4] ),
    .A1(\s0.data_out[20][4] ),
    .S(net1470),
    .X(_1011_));
 sg13g2_nor2b_1 _5014_ (.A(net1462),
    .B_N(net1338),
    .Y(_1012_));
 sg13g2_a21oi_1 _5015_ (.A1(net1469),
    .A2(_1011_),
    .Y(_1013_),
    .B1(_1012_));
 sg13g2_nand2b_1 _5016_ (.Y(_1014_),
    .B(net1476),
    .A_N(_1013_));
 sg13g2_o21ai_1 _5017_ (.B1(_0895_),
    .Y(_1015_),
    .A1(net1482),
    .A2(_3447_));
 sg13g2_nand2_1 _5018_ (.Y(_1016_),
    .A(net1173),
    .B(_1015_));
 sg13g2_nand3_1 _5019_ (.B(_1014_),
    .C(_1016_),
    .A(net1670),
    .Y(_1017_));
 sg13g2_a21oi_1 _5020_ (.A1(_1014_),
    .A2(_1016_),
    .Y(_1018_),
    .B1(net1670));
 sg13g2_nor2_1 _5021_ (.A(net1660),
    .B(_1008_),
    .Y(_1019_));
 sg13g2_nor2_1 _5022_ (.A(net1678),
    .B(_0980_),
    .Y(_1020_));
 sg13g2_nor3_1 _5023_ (.A(_1018_),
    .B(_1019_),
    .C(_1020_),
    .Y(_1021_));
 sg13g2_nand3_1 _5024_ (.B(_1017_),
    .C(_1021_),
    .A(_1009_),
    .Y(_1022_));
 sg13g2_or3_1 _5025_ (.A(_0983_),
    .B(_1001_),
    .C(_1022_),
    .X(_1023_));
 sg13g2_o21ai_1 _5026_ (.B1(_1009_),
    .Y(_1024_),
    .A1(_1017_),
    .A2(_1019_));
 sg13g2_nor2b_1 _5027_ (.A(_1001_),
    .B_N(_1024_),
    .Y(_1025_));
 sg13g2_nor2b_1 _5028_ (.A(_0998_),
    .B_N(_1000_),
    .Y(_1026_));
 sg13g2_nor4_1 _5029_ (.A(_0942_),
    .B(_0943_),
    .C(_1025_),
    .D(_1026_),
    .Y(_1027_));
 sg13g2_or2_1 _5030_ (.X(_1028_),
    .B(net1558),
    .A(net387));
 sg13g2_a21oi_1 _5031_ (.A1(_1023_),
    .A2(_1027_),
    .Y(_0183_),
    .B1(_1028_));
 sg13g2_a21oi_1 _5032_ (.A1(net1463),
    .A2(\s0.data_out[20][0] ),
    .Y(_1029_),
    .B1(_0967_));
 sg13g2_a21oi_1 _5033_ (.A1(net1171),
    .A2(_0969_),
    .Y(_1030_),
    .B1(net1595));
 sg13g2_o21ai_1 _5034_ (.B1(_1030_),
    .Y(_1031_),
    .A1(net1172),
    .A2(_1029_));
 sg13g2_o21ai_1 _5035_ (.B1(_1031_),
    .Y(_1032_),
    .A1(net1723),
    .A2(net713));
 sg13g2_inv_1 _5036_ (.Y(_0184_),
    .A(net714));
 sg13g2_a21oi_1 _5037_ (.A1(net1463),
    .A2(\s0.data_out[20][1] ),
    .Y(_1033_),
    .B1(_0957_));
 sg13g2_a21oi_1 _5038_ (.A1(net1171),
    .A2(_0962_),
    .Y(_1034_),
    .B1(net1595));
 sg13g2_o21ai_1 _5039_ (.B1(_1034_),
    .Y(_1035_),
    .A1(net1171),
    .A2(_1033_));
 sg13g2_o21ai_1 _5040_ (.B1(_1035_),
    .Y(_1036_),
    .A1(net1722),
    .A2(net551));
 sg13g2_inv_1 _5041_ (.Y(_0185_),
    .A(net552));
 sg13g2_a21oi_1 _5042_ (.A1(net1463),
    .A2(\s0.data_out[20][2] ),
    .Y(_1037_),
    .B1(_0952_));
 sg13g2_a21oi_1 _5043_ (.A1(net1171),
    .A2(_0954_),
    .Y(_1038_),
    .B1(net1595));
 sg13g2_o21ai_1 _5044_ (.B1(_1038_),
    .Y(_1039_),
    .A1(net1171),
    .A2(_1037_));
 sg13g2_o21ai_1 _5045_ (.B1(_1039_),
    .Y(_1040_),
    .A1(net1722),
    .A2(net520));
 sg13g2_inv_1 _5046_ (.Y(_0186_),
    .A(net521));
 sg13g2_and2_1 _5047_ (.A(net1465),
    .B(\s0.data_out[20][3] ),
    .X(_1041_));
 sg13g2_o21ai_1 _5048_ (.B1(net1481),
    .Y(_1042_),
    .A1(_0976_),
    .A2(_1041_));
 sg13g2_nor2_1 _5049_ (.A(net1593),
    .B(_0979_),
    .Y(_1043_));
 sg13g2_a22oi_1 _5050_ (.Y(_0187_),
    .B1(_1042_),
    .B2(_1043_),
    .A2(_3443_),
    .A1(net1593));
 sg13g2_a21oi_1 _5051_ (.A1(net1461),
    .A2(net516),
    .Y(_1044_),
    .B1(_1012_));
 sg13g2_a21oi_1 _5052_ (.A1(net1173),
    .A2(_1015_),
    .Y(_1045_),
    .B1(net1594));
 sg13g2_o21ai_1 _5053_ (.B1(_1045_),
    .Y(_1046_),
    .A1(net1173),
    .A2(_1044_));
 sg13g2_o21ai_1 _5054_ (.B1(_1046_),
    .Y(_1047_),
    .A1(net1724),
    .A2(net702));
 sg13g2_inv_1 _5055_ (.Y(_0188_),
    .A(_1047_));
 sg13g2_and2_1 _5056_ (.A(net1462),
    .B(net492),
    .X(_1048_));
 sg13g2_o21ai_1 _5057_ (.B1(net1476),
    .Y(_1049_),
    .A1(_1004_),
    .A2(_1048_));
 sg13g2_nor2_1 _5058_ (.A(net1592),
    .B(net450),
    .Y(_1050_));
 sg13g2_a22oi_1 _5059_ (.Y(_0189_),
    .B1(_1049_),
    .B2(_1050_),
    .A2(_3442_),
    .A1(net1592));
 sg13g2_and2_1 _5060_ (.A(net1461),
    .B(\s0.data_out[20][6] ),
    .X(_1051_));
 sg13g2_o21ai_1 _5061_ (.B1(net1475),
    .Y(_1052_),
    .A1(_0993_),
    .A2(_1051_));
 sg13g2_nand3b_1 _5062_ (.B(_1052_),
    .C(net1724),
    .Y(_1053_),
    .A_N(_0996_));
 sg13g2_o21ai_1 _5063_ (.B1(net836),
    .Y(_1054_),
    .A1(net1724),
    .A2(net715));
 sg13g2_inv_1 _5064_ (.Y(_0190_),
    .A(_1054_));
 sg13g2_and2_1 _5065_ (.A(net1462),
    .B(\s0.data_out[20][7] ),
    .X(_1055_));
 sg13g2_o21ai_1 _5066_ (.B1(net1475),
    .Y(_1056_),
    .A1(_0986_),
    .A2(_1055_));
 sg13g2_nor2_1 _5067_ (.A(net1592),
    .B(_0989_),
    .Y(_1057_));
 sg13g2_a22oi_1 _5068_ (.Y(_0191_),
    .B1(_1056_),
    .B2(_1057_),
    .A2(_3441_),
    .A1(net1592));
 sg13g2_and2_1 _5069_ (.A(net1724),
    .B(net376),
    .X(_0192_));
 sg13g2_o21ai_1 _5070_ (.B1(net1467),
    .Y(_1058_),
    .A1(net1632),
    .A2(net1453));
 sg13g2_nand2_1 _5071_ (.Y(_1059_),
    .A(net1623),
    .B(net1457));
 sg13g2_nand2b_1 _5072_ (.Y(_1060_),
    .B(_1059_),
    .A_N(_1058_));
 sg13g2_o21ai_1 _5073_ (.B1(_1060_),
    .Y(_1061_),
    .A1(net1466),
    .A2(_0941_));
 sg13g2_nor2_1 _5074_ (.A(net409),
    .B(net1457),
    .Y(_1062_));
 sg13g2_or2_1 _5075_ (.X(_1063_),
    .B(_1062_),
    .A(_1060_));
 sg13g2_nor2_1 _5076_ (.A(net1453),
    .B(_1058_),
    .Y(_1064_));
 sg13g2_a21oi_1 _5077_ (.A1(_3367_),
    .A2(_3392_),
    .Y(_1065_),
    .B1(net1466));
 sg13g2_nor2_1 _5078_ (.A(_1064_),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_o21ai_1 _5079_ (.B1(net1724),
    .Y(_1067_),
    .A1(net618),
    .A2(_1061_));
 sg13g2_a21oi_1 _5080_ (.A1(_1063_),
    .A2(_1066_),
    .Y(_0193_),
    .B1(_1067_));
 sg13g2_nor2_1 _5081_ (.A(net1594),
    .B(_1061_),
    .Y(_0194_));
 sg13g2_and2_1 _5082_ (.A(net1713),
    .B(net395),
    .X(_0195_));
 sg13g2_nand2_1 _5083_ (.Y(_1068_),
    .A(net1460),
    .B(net662));
 sg13g2_mux2_1 _5084_ (.A0(\s0.data_out[20][2] ),
    .A1(\s0.data_out[19][2] ),
    .S(net1457),
    .X(_1069_));
 sg13g2_nor2b_1 _5085_ (.A(net1451),
    .B_N(net1342),
    .Y(_1070_));
 sg13g2_a21o_1 _5086_ (.A2(_1069_),
    .A1(net1451),
    .B1(_1070_),
    .X(_1071_));
 sg13g2_nand2b_1 _5087_ (.Y(_1072_),
    .B(net662),
    .A_N(net1471));
 sg13g2_a21oi_1 _5088_ (.A1(_0950_),
    .A2(_1072_),
    .Y(_1073_),
    .B1(net1465));
 sg13g2_a21oi_1 _5089_ (.A1(net1465),
    .A2(_1071_),
    .Y(_1074_),
    .B1(_1073_));
 sg13g2_or2_1 _5090_ (.X(_1075_),
    .B(_1074_),
    .A(net1686));
 sg13g2_nand2_1 _5091_ (.Y(_1076_),
    .A(net1458),
    .B(net725));
 sg13g2_o21ai_1 _5092_ (.B1(_1076_),
    .Y(_1077_),
    .A1(net1457),
    .A2(_3450_));
 sg13g2_nor2b_1 _5093_ (.A(net1451),
    .B_N(net1346),
    .Y(_1078_));
 sg13g2_a21o_1 _5094_ (.A2(_1077_),
    .A1(net1451),
    .B1(_1078_),
    .X(_1079_));
 sg13g2_nand2_1 _5095_ (.Y(_1080_),
    .A(_3392_),
    .B(\s0.data_out[19][1] ));
 sg13g2_a21oi_1 _5096_ (.A1(_0958_),
    .A2(_1080_),
    .Y(_1081_),
    .B1(net1468));
 sg13g2_a21oi_1 _5097_ (.A1(net1468),
    .A2(_1079_),
    .Y(_1082_),
    .B1(_1081_));
 sg13g2_mux2_1 _5098_ (.A0(\s0.data_out[20][0] ),
    .A1(\s0.data_out[19][0] ),
    .S(net1457),
    .X(_1083_));
 sg13g2_nor2b_1 _5099_ (.A(net1451),
    .B_N(net1350),
    .Y(_1084_));
 sg13g2_a21oi_1 _5100_ (.A1(net1451),
    .A2(_1083_),
    .Y(_1085_),
    .B1(_1084_));
 sg13g2_nand2b_1 _5101_ (.Y(_1086_),
    .B(net1465),
    .A_N(_1085_));
 sg13g2_mux2_1 _5102_ (.A0(\s0.data_out[19][0] ),
    .A1(\s0.data_out[20][0] ),
    .S(net1471),
    .X(_1087_));
 sg13g2_nand2b_1 _5103_ (.Y(_1088_),
    .B(_1087_),
    .A_N(net1465));
 sg13g2_a221oi_1 _5104_ (.B2(_1088_),
    .C1(net1702),
    .B1(_1086_),
    .A1(net1695),
    .Y(_1089_),
    .A2(_1082_));
 sg13g2_o21ai_1 _5105_ (.B1(_1075_),
    .Y(_1090_),
    .A1(net1695),
    .A2(_1082_));
 sg13g2_nand2_1 _5106_ (.Y(_1091_),
    .A(net1458),
    .B(net656));
 sg13g2_o21ai_1 _5107_ (.B1(_1091_),
    .Y(_1092_),
    .A1(net1457),
    .A2(_3448_));
 sg13g2_nor2_1 _5108_ (.A(net1452),
    .B(net1161),
    .Y(_1093_));
 sg13g2_a21o_1 _5109_ (.A2(_1092_),
    .A1(net1452),
    .B1(_1093_),
    .X(_1094_));
 sg13g2_nand2_1 _5110_ (.Y(_1095_),
    .A(_3392_),
    .B(\s0.data_out[19][3] ));
 sg13g2_a21oi_1 _5111_ (.A1(_0974_),
    .A2(_1095_),
    .Y(_1096_),
    .B1(net1468));
 sg13g2_a21oi_1 _5112_ (.A1(net1469),
    .A2(_1094_),
    .Y(_1097_),
    .B1(_1096_));
 sg13g2_a22oi_1 _5113_ (.Y(_1098_),
    .B1(_1097_),
    .B2(net1680),
    .A2(_1074_),
    .A1(net1686));
 sg13g2_o21ai_1 _5114_ (.B1(_1098_),
    .Y(_1099_),
    .A1(_1089_),
    .A2(_1090_));
 sg13g2_nand2_1 _5115_ (.Y(_1100_),
    .A(net1459),
    .B(net764));
 sg13g2_mux2_1 _5116_ (.A0(\s0.data_out[20][6] ),
    .A1(\s0.data_out[19][6] ),
    .S(net1459),
    .X(_1101_));
 sg13g2_nor2b_1 _5117_ (.A(net1454),
    .B_N(net1328),
    .Y(_1102_));
 sg13g2_a21o_1 _5118_ (.A2(_1101_),
    .A1(net1454),
    .B1(_1102_),
    .X(_1103_));
 sg13g2_nand2b_1 _5119_ (.Y(_1104_),
    .B(net764),
    .A_N(net1472));
 sg13g2_a21oi_1 _5120_ (.A1(_0991_),
    .A2(_1104_),
    .Y(_1105_),
    .B1(net1466));
 sg13g2_a21oi_1 _5121_ (.A1(net1467),
    .A2(_1103_),
    .Y(_1106_),
    .B1(_1105_));
 sg13g2_nand2_1 _5122_ (.Y(_1107_),
    .A(net1459),
    .B(net755));
 sg13g2_mux2_1 _5123_ (.A0(\s0.data_out[20][7] ),
    .A1(\s0.data_out[19][7] ),
    .S(net1459),
    .X(_1108_));
 sg13g2_nor2b_1 _5124_ (.A(net1454),
    .B_N(net1323),
    .Y(_1109_));
 sg13g2_a21o_1 _5125_ (.A2(_1108_),
    .A1(net1454),
    .B1(_1109_),
    .X(_1110_));
 sg13g2_nand2b_1 _5126_ (.Y(_1111_),
    .B(\s0.data_out[19][7] ),
    .A_N(net1472));
 sg13g2_a21oi_1 _5127_ (.A1(_0984_),
    .A2(_1111_),
    .Y(_1112_),
    .B1(net1467));
 sg13g2_a21oi_1 _5128_ (.A1(net1467),
    .A2(_1110_),
    .Y(_1113_),
    .B1(_1112_));
 sg13g2_a22oi_1 _5129_ (.Y(_1114_),
    .B1(_1113_),
    .B2(net1643),
    .A2(_1106_),
    .A1(net1653));
 sg13g2_nor2_1 _5130_ (.A(net1653),
    .B(_1106_),
    .Y(_1115_));
 sg13g2_or2_1 _5131_ (.X(_1116_),
    .B(_1113_),
    .A(net1643));
 sg13g2_nand3b_1 _5132_ (.B(_1116_),
    .C(_1114_),
    .Y(_1117_),
    .A_N(_1115_));
 sg13g2_nand2_1 _5133_ (.Y(_1118_),
    .A(net1459),
    .B(net790));
 sg13g2_o21ai_1 _5134_ (.B1(_1118_),
    .Y(_1119_),
    .A1(net1457),
    .A2(_3447_));
 sg13g2_nor2b_1 _5135_ (.A(net1453),
    .B_N(net1337),
    .Y(_1120_));
 sg13g2_a21o_1 _5136_ (.A2(_1119_),
    .A1(net1453),
    .B1(_1120_),
    .X(_1121_));
 sg13g2_nand2_1 _5137_ (.Y(_1122_),
    .A(_3392_),
    .B(\s0.data_out[19][4] ));
 sg13g2_a21oi_1 _5138_ (.A1(_1010_),
    .A2(_1122_),
    .Y(_1123_),
    .B1(net1466));
 sg13g2_a21oi_1 _5139_ (.A1(net1466),
    .A2(_1121_),
    .Y(_1124_),
    .B1(_1123_));
 sg13g2_nand2_1 _5140_ (.Y(_1125_),
    .A(net1460),
    .B(\s0.data_out[19][5] ));
 sg13g2_mux2_1 _5141_ (.A0(\s0.data_out[20][5] ),
    .A1(\s0.data_out[19][5] ),
    .S(net1457),
    .X(_1126_));
 sg13g2_nor2b_1 _5142_ (.A(net1453),
    .B_N(net1332),
    .Y(_1127_));
 sg13g2_a21o_1 _5143_ (.A2(_1126_),
    .A1(net1453),
    .B1(_1127_),
    .X(_1128_));
 sg13g2_nand2b_1 _5144_ (.Y(_1129_),
    .B(\s0.data_out[19][5] ),
    .A_N(net1472));
 sg13g2_a21oi_1 _5145_ (.A1(_1002_),
    .A2(_1129_),
    .Y(_1130_),
    .B1(net1461));
 sg13g2_a21oi_1 _5146_ (.A1(net1466),
    .A2(_1128_),
    .Y(_1131_),
    .B1(_1130_));
 sg13g2_nor2_1 _5147_ (.A(net1661),
    .B(_1131_),
    .Y(_1132_));
 sg13g2_nand2_1 _5148_ (.Y(_1133_),
    .A(net1661),
    .B(_1131_));
 sg13g2_o21ai_1 _5149_ (.B1(_1133_),
    .Y(_1134_),
    .A1(net1680),
    .A2(_1097_));
 sg13g2_xnor2_1 _5150_ (.Y(_1135_),
    .A(net1671),
    .B(_1124_));
 sg13g2_nor4_1 _5151_ (.A(_1117_),
    .B(_1132_),
    .C(_1134_),
    .D(_1135_),
    .Y(_1136_));
 sg13g2_nand2_1 _5152_ (.Y(_1137_),
    .A(_1099_),
    .B(_1136_));
 sg13g2_nand3b_1 _5153_ (.B(_1124_),
    .C(net1671),
    .Y(_1138_),
    .A_N(_1132_));
 sg13g2_a21oi_1 _5154_ (.A1(_1133_),
    .A2(_1138_),
    .Y(_1139_),
    .B1(_1117_));
 sg13g2_nor2b_1 _5155_ (.A(_1114_),
    .B_N(_1116_),
    .Y(_1140_));
 sg13g2_nor3_1 _5156_ (.A(_1061_),
    .B(_1139_),
    .C(_1140_),
    .Y(_1141_));
 sg13g2_or2_1 _5157_ (.X(_1142_),
    .B(net1557),
    .A(net376));
 sg13g2_a21oi_1 _5158_ (.A1(_1137_),
    .A2(_1141_),
    .Y(_0196_),
    .B1(_1142_));
 sg13g2_and2_1 _5159_ (.A(net1451),
    .B(\s0.data_out[19][0] ),
    .X(_1143_));
 sg13g2_o21ai_1 _5160_ (.B1(net1465),
    .Y(_1144_),
    .A1(_1084_),
    .A2(_1143_));
 sg13g2_nand3_1 _5161_ (.B(_1088_),
    .C(_1144_),
    .A(net1725),
    .Y(_1145_));
 sg13g2_o21ai_1 _5162_ (.B1(_1145_),
    .Y(_1146_),
    .A1(net1725),
    .A2(net733));
 sg13g2_inv_1 _5163_ (.Y(_0197_),
    .A(_1146_));
 sg13g2_nor2_1 _5164_ (.A(net1191),
    .B(_3456_),
    .Y(_1147_));
 sg13g2_o21ai_1 _5165_ (.B1(net1468),
    .Y(_1148_),
    .A1(_1078_),
    .A2(_1147_));
 sg13g2_nor2_1 _5166_ (.A(net1594),
    .B(_1081_),
    .Y(_1149_));
 sg13g2_a22oi_1 _5167_ (.Y(_0198_),
    .B1(_1148_),
    .B2(_1149_),
    .A2(_3450_),
    .A1(net1595));
 sg13g2_nor2_1 _5168_ (.A(net1191),
    .B(_3455_),
    .Y(_1150_));
 sg13g2_o21ai_1 _5169_ (.B1(net1468),
    .Y(_1151_),
    .A1(_1070_),
    .A2(_1150_));
 sg13g2_nor2_1 _5170_ (.A(net1595),
    .B(_1073_),
    .Y(_1152_));
 sg13g2_a22oi_1 _5171_ (.Y(_0199_),
    .B1(_1151_),
    .B2(_1152_),
    .A2(_3449_),
    .A1(net1595));
 sg13g2_nor2_1 _5172_ (.A(net1191),
    .B(_3454_),
    .Y(_1153_));
 sg13g2_o21ai_1 _5173_ (.B1(net1468),
    .Y(_1154_),
    .A1(_1093_),
    .A2(_1153_));
 sg13g2_nor2_1 _5174_ (.A(net1605),
    .B(_1096_),
    .Y(_1155_));
 sg13g2_a22oi_1 _5175_ (.Y(_0200_),
    .B1(_1154_),
    .B2(_1155_),
    .A2(_3448_),
    .A1(net1605));
 sg13g2_nor2_1 _5176_ (.A(net1191),
    .B(_3453_),
    .Y(_1156_));
 sg13g2_o21ai_1 _5177_ (.B1(net1466),
    .Y(_1157_),
    .A1(_1120_),
    .A2(_1156_));
 sg13g2_nor2_1 _5178_ (.A(net1594),
    .B(_1123_),
    .Y(_1158_));
 sg13g2_a22oi_1 _5179_ (.Y(_0201_),
    .B1(_1157_),
    .B2(_1158_),
    .A2(_3447_),
    .A1(net1594));
 sg13g2_and2_1 _5180_ (.A(net1453),
    .B(\s0.data_out[19][5] ),
    .X(_1159_));
 sg13g2_o21ai_1 _5181_ (.B1(net1461),
    .Y(_1160_),
    .A1(_1127_),
    .A2(_1159_));
 sg13g2_nor2_1 _5182_ (.A(net1594),
    .B(_1130_),
    .Y(_1161_));
 sg13g2_a22oi_1 _5183_ (.Y(_0202_),
    .B1(_1160_),
    .B2(_1161_),
    .A2(_3446_),
    .A1(net1594));
 sg13g2_nor2_1 _5184_ (.A(net1191),
    .B(_3452_),
    .Y(_1162_));
 sg13g2_o21ai_1 _5185_ (.B1(net1466),
    .Y(_1163_),
    .A1(_1102_),
    .A2(_1162_));
 sg13g2_nand3b_1 _5186_ (.B(_1163_),
    .C(net1731),
    .Y(_1164_),
    .A_N(_1105_));
 sg13g2_o21ai_1 _5187_ (.B1(_1164_),
    .Y(_1165_),
    .A1(net1731),
    .A2(net781));
 sg13g2_inv_1 _5188_ (.Y(_0203_),
    .A(_1165_));
 sg13g2_nor2_1 _5189_ (.A(net1192),
    .B(_3451_),
    .Y(_1166_));
 sg13g2_o21ai_1 _5190_ (.B1(net1467),
    .Y(_1167_),
    .A1(_1109_),
    .A2(_1166_));
 sg13g2_nor2_1 _5191_ (.A(net1605),
    .B(_1112_),
    .Y(_1168_));
 sg13g2_a22oi_1 _5192_ (.Y(_0204_),
    .B1(_1167_),
    .B2(_1168_),
    .A2(_3445_),
    .A1(net1605));
 sg13g2_o21ai_1 _5193_ (.B1(net1455),
    .Y(_1169_),
    .A1(net1632),
    .A2(net1441));
 sg13g2_a21oi_1 _5194_ (.A1(net1623),
    .A2(net1447),
    .Y(_1170_),
    .B1(_1169_));
 sg13g2_o21ai_1 _5195_ (.B1(_1170_),
    .Y(_1171_),
    .A1(\s0.was_valid_out[18] [0]),
    .A2(net1447));
 sg13g2_nor2_1 _5196_ (.A(net1441),
    .B(_1169_),
    .Y(_1172_));
 sg13g2_o21ai_1 _5197_ (.B1(net1192),
    .Y(_1173_),
    .A1(\s0.was_valid_out[18] [0]),
    .A2(net1459));
 sg13g2_nand2_1 _5198_ (.Y(_1174_),
    .A(_1171_),
    .B(_1173_));
 sg13g2_a21oi_2 _5199_ (.B1(_1170_),
    .Y(_1175_),
    .A2(_1059_),
    .A1(net1191));
 sg13g2_o21ai_1 _5200_ (.B1(net1731),
    .Y(_1176_),
    .A1(_1172_),
    .A2(_1174_));
 sg13g2_a21oi_1 _5201_ (.A1(_3367_),
    .A2(_1175_),
    .Y(_0205_),
    .B1(_1176_));
 sg13g2_and2_1 _5202_ (.A(net1731),
    .B(_1175_),
    .X(_0206_));
 sg13g2_and2_1 _5203_ (.A(net1733),
    .B(net381),
    .X(_0207_));
 sg13g2_nand2_1 _5204_ (.Y(_1177_),
    .A(net1448),
    .B(net627));
 sg13g2_mux2_1 _5205_ (.A0(\s0.data_out[19][2] ),
    .A1(\s0.data_out[18][2] ),
    .S(net1447),
    .X(_1178_));
 sg13g2_nor2b_1 _5206_ (.A(net1440),
    .B_N(net1342),
    .Y(_1179_));
 sg13g2_a21o_1 _5207_ (.A2(_1178_),
    .A1(net1441),
    .B1(_1179_),
    .X(_1180_));
 sg13g2_nand2b_1 _5208_ (.Y(_1181_),
    .B(net627),
    .A_N(net1460));
 sg13g2_a21oi_1 _5209_ (.A1(_1068_),
    .A2(_1181_),
    .Y(_1182_),
    .B1(net1456));
 sg13g2_a21oi_1 _5210_ (.A1(net1456),
    .A2(_1180_),
    .Y(_1183_),
    .B1(_1182_));
 sg13g2_or2_1 _5211_ (.X(_1184_),
    .B(_1183_),
    .A(net1686));
 sg13g2_nand2_1 _5212_ (.Y(_1185_),
    .A(net1447),
    .B(\s0.data_out[18][1] ));
 sg13g2_o21ai_1 _5213_ (.B1(_1185_),
    .Y(_1186_),
    .A1(net1447),
    .A2(_3456_));
 sg13g2_nor2b_1 _5214_ (.A(net1440),
    .B_N(net1346),
    .Y(_1187_));
 sg13g2_a21o_1 _5215_ (.A2(_1186_),
    .A1(net1440),
    .B1(_1187_),
    .X(_1188_));
 sg13g2_nand2b_1 _5216_ (.Y(_1189_),
    .B(\s0.data_out[18][1] ),
    .A_N(net1458));
 sg13g2_a21oi_1 _5217_ (.A1(_1076_),
    .A2(_1189_),
    .Y(_1190_),
    .B1(net1452));
 sg13g2_a21oi_1 _5218_ (.A1(net1452),
    .A2(_1188_),
    .Y(_1191_),
    .B1(_1190_));
 sg13g2_mux2_1 _5219_ (.A0(\s0.data_out[19][0] ),
    .A1(\s0.data_out[18][0] ),
    .S(net1447),
    .X(_1192_));
 sg13g2_nor2b_1 _5220_ (.A(net1440),
    .B_N(net1350),
    .Y(_1193_));
 sg13g2_a21oi_1 _5221_ (.A1(net1440),
    .A2(_1192_),
    .Y(_1194_),
    .B1(_1193_));
 sg13g2_nand2b_1 _5222_ (.Y(_1195_),
    .B(net1452),
    .A_N(_1194_));
 sg13g2_mux2_1 _5223_ (.A0(\s0.data_out[18][0] ),
    .A1(\s0.data_out[19][0] ),
    .S(net1458),
    .X(_1196_));
 sg13g2_nand2_1 _5224_ (.Y(_1197_),
    .A(net1191),
    .B(_1196_));
 sg13g2_a221oi_1 _5225_ (.B2(_1197_),
    .C1(net1702),
    .B1(_1195_),
    .A1(net1696),
    .Y(_1198_),
    .A2(_1191_));
 sg13g2_o21ai_1 _5226_ (.B1(_1184_),
    .Y(_1199_),
    .A1(net1696),
    .A2(_1191_));
 sg13g2_nand2_1 _5227_ (.Y(_1200_),
    .A(net1448),
    .B(net482));
 sg13g2_o21ai_1 _5228_ (.B1(_1200_),
    .Y(_1201_),
    .A1(net1448),
    .A2(_3454_));
 sg13g2_nor2_1 _5229_ (.A(net1443),
    .B(net1161),
    .Y(_1202_));
 sg13g2_a21o_1 _5230_ (.A2(_1201_),
    .A1(net1443),
    .B1(_1202_),
    .X(_1203_));
 sg13g2_nand2b_1 _5231_ (.Y(_1204_),
    .B(net482),
    .A_N(net1460));
 sg13g2_a21oi_1 _5232_ (.A1(_1091_),
    .A2(_1204_),
    .Y(_1205_),
    .B1(net1456));
 sg13g2_a21oi_1 _5233_ (.A1(net1456),
    .A2(_1203_),
    .Y(_1206_),
    .B1(_1205_));
 sg13g2_a22oi_1 _5234_ (.Y(_1207_),
    .B1(_1206_),
    .B2(net1680),
    .A2(_1183_),
    .A1(net1686));
 sg13g2_o21ai_1 _5235_ (.B1(_1207_),
    .Y(_1208_),
    .A1(_1198_),
    .A2(_1199_));
 sg13g2_nand2_1 _5236_ (.Y(_1209_),
    .A(net1449),
    .B(\s0.data_out[18][6] ));
 sg13g2_mux2_1 _5237_ (.A0(\s0.data_out[19][6] ),
    .A1(\s0.data_out[18][6] ),
    .S(net1448),
    .X(_1210_));
 sg13g2_nor2b_1 _5238_ (.A(net1441),
    .B_N(net1328),
    .Y(_1211_));
 sg13g2_a21o_1 _5239_ (.A2(_1210_),
    .A1(net1442),
    .B1(_1211_),
    .X(_1212_));
 sg13g2_nand2b_1 _5240_ (.Y(_1213_),
    .B(\s0.data_out[18][6] ),
    .A_N(net1459));
 sg13g2_a21oi_1 _5241_ (.A1(_1100_),
    .A2(_1213_),
    .Y(_1214_),
    .B1(net1454));
 sg13g2_a21oi_1 _5242_ (.A1(net1454),
    .A2(_1212_),
    .Y(_1215_),
    .B1(_1214_));
 sg13g2_nand2_1 _5243_ (.Y(_1216_),
    .A(net1449),
    .B(net805));
 sg13g2_mux2_1 _5244_ (.A0(\s0.data_out[19][7] ),
    .A1(\s0.data_out[18][7] ),
    .S(net1448),
    .X(_1217_));
 sg13g2_nor2b_1 _5245_ (.A(net1442),
    .B_N(net1323),
    .Y(_1218_));
 sg13g2_a21o_1 _5246_ (.A2(_1217_),
    .A1(net1442),
    .B1(_1218_),
    .X(_1219_));
 sg13g2_nand2b_1 _5247_ (.Y(_1220_),
    .B(\s0.data_out[18][7] ),
    .A_N(net1460));
 sg13g2_a21oi_1 _5248_ (.A1(_1107_),
    .A2(_1220_),
    .Y(_1221_),
    .B1(net1455));
 sg13g2_a21oi_1 _5249_ (.A1(net1455),
    .A2(_1219_),
    .Y(_1222_),
    .B1(_1221_));
 sg13g2_a22oi_1 _5250_ (.Y(_1223_),
    .B1(_1222_),
    .B2(net1643),
    .A2(_1215_),
    .A1(net1653));
 sg13g2_or2_1 _5251_ (.X(_1224_),
    .B(_1215_),
    .A(net1653));
 sg13g2_nor2_1 _5252_ (.A(net1643),
    .B(_1222_),
    .Y(_1225_));
 sg13g2_nand3b_1 _5253_ (.B(_1223_),
    .C(_1224_),
    .Y(_1226_),
    .A_N(_1225_));
 sg13g2_nand2_1 _5254_ (.Y(_1227_),
    .A(net1449),
    .B(net574));
 sg13g2_mux2_1 _5255_ (.A0(\s0.data_out[19][5] ),
    .A1(\s0.data_out[18][5] ),
    .S(net1449),
    .X(_1228_));
 sg13g2_nor2b_1 _5256_ (.A(net1444),
    .B_N(net1333),
    .Y(_1229_));
 sg13g2_a21oi_1 _5257_ (.A1(net1444),
    .A2(_1228_),
    .Y(_1230_),
    .B1(_1229_));
 sg13g2_nand2b_1 _5258_ (.Y(_1231_),
    .B(net1456),
    .A_N(_1230_));
 sg13g2_o21ai_1 _5259_ (.B1(_1125_),
    .Y(_1232_),
    .A1(net1460),
    .A2(_3458_));
 sg13g2_nand2_1 _5260_ (.Y(_1233_),
    .A(net1192),
    .B(_1232_));
 sg13g2_nand3_1 _5261_ (.B(_1231_),
    .C(_1233_),
    .A(net1661),
    .Y(_1234_));
 sg13g2_nor2b_1 _5262_ (.A(net1442),
    .B_N(net1337),
    .Y(_1235_));
 sg13g2_nand2_1 _5263_ (.Y(_1236_),
    .A(net1449),
    .B(net598));
 sg13g2_mux2_1 _5264_ (.A0(\s0.data_out[19][4] ),
    .A1(\s0.data_out[18][4] ),
    .S(net1448),
    .X(_1237_));
 sg13g2_a21o_1 _5265_ (.A2(_1237_),
    .A1(net1442),
    .B1(_1235_),
    .X(_1238_));
 sg13g2_nand2b_1 _5266_ (.Y(_1239_),
    .B(net598),
    .A_N(net1459));
 sg13g2_a21oi_1 _5267_ (.A1(_1118_),
    .A2(_1239_),
    .Y(_1240_),
    .B1(net1454));
 sg13g2_a21oi_1 _5268_ (.A1(net1455),
    .A2(_1238_),
    .Y(_1241_),
    .B1(_1240_));
 sg13g2_nand2_1 _5269_ (.Y(_1242_),
    .A(net1671),
    .B(_1241_));
 sg13g2_nand2_1 _5270_ (.Y(_1243_),
    .A(_1234_),
    .B(_1242_));
 sg13g2_nor2_1 _5271_ (.A(net1671),
    .B(_1241_),
    .Y(_1244_));
 sg13g2_a21o_1 _5272_ (.A2(_1233_),
    .A1(_1231_),
    .B1(net1661),
    .X(_1245_));
 sg13g2_o21ai_1 _5273_ (.B1(_1245_),
    .Y(_1246_),
    .A1(net1682),
    .A2(_1206_));
 sg13g2_nor4_1 _5274_ (.A(_1226_),
    .B(_1243_),
    .C(_1244_),
    .D(_1246_),
    .Y(_1247_));
 sg13g2_nor2b_1 _5275_ (.A(_1226_),
    .B_N(_1243_),
    .Y(_1248_));
 sg13g2_o21ai_1 _5276_ (.B1(_1175_),
    .Y(_1249_),
    .A1(_1223_),
    .A2(_1225_));
 sg13g2_a221oi_1 _5277_ (.B2(_1245_),
    .C1(_1249_),
    .B1(_1248_),
    .A1(_1208_),
    .Y(_1250_),
    .A2(_1247_));
 sg13g2_nor3_1 _5278_ (.A(net370),
    .B(net1557),
    .C(_1250_),
    .Y(_0208_));
 sg13g2_a21oi_1 _5279_ (.A1(net1440),
    .A2(\s0.data_out[18][0] ),
    .Y(_1251_),
    .B1(_1193_));
 sg13g2_a21oi_1 _5280_ (.A1(net1191),
    .A2(_1196_),
    .Y(_1252_),
    .B1(net1608));
 sg13g2_o21ai_1 _5281_ (.B1(_1252_),
    .Y(_1253_),
    .A1(net1192),
    .A2(_1251_));
 sg13g2_o21ai_1 _5282_ (.B1(_1253_),
    .Y(_1254_),
    .A1(net1724),
    .A2(net683));
 sg13g2_inv_1 _5283_ (.Y(_0209_),
    .A(net684));
 sg13g2_and2_1 _5284_ (.A(net1440),
    .B(\s0.data_out[18][1] ),
    .X(_1255_));
 sg13g2_o21ai_1 _5285_ (.B1(net1451),
    .Y(_1256_),
    .A1(_1187_),
    .A2(_1255_));
 sg13g2_nor2_1 _5286_ (.A(net1608),
    .B(_1190_),
    .Y(_1257_));
 sg13g2_a22oi_1 _5287_ (.Y(_0210_),
    .B1(_1256_),
    .B2(_1257_),
    .A2(_3456_),
    .A1(net1608));
 sg13g2_nor2_1 _5288_ (.A(net1196),
    .B(_3461_),
    .Y(_1258_));
 sg13g2_o21ai_1 _5289_ (.B1(net1456),
    .Y(_1259_),
    .A1(_1179_),
    .A2(_1258_));
 sg13g2_nor2_1 _5290_ (.A(net1605),
    .B(_1182_),
    .Y(_1260_));
 sg13g2_a22oi_1 _5291_ (.Y(_0211_),
    .B1(_1259_),
    .B2(_1260_),
    .A2(_3455_),
    .A1(net1605));
 sg13g2_nor2_1 _5292_ (.A(net1197),
    .B(_3460_),
    .Y(_1261_));
 sg13g2_o21ai_1 _5293_ (.B1(net1456),
    .Y(_1262_),
    .A1(_1202_),
    .A2(_1261_));
 sg13g2_nor2_1 _5294_ (.A(net1606),
    .B(_1205_),
    .Y(_1263_));
 sg13g2_a22oi_1 _5295_ (.Y(_0212_),
    .B1(_1262_),
    .B2(_1263_),
    .A2(_3454_),
    .A1(net1606));
 sg13g2_nor2_1 _5296_ (.A(net1197),
    .B(_3459_),
    .Y(_1264_));
 sg13g2_o21ai_1 _5297_ (.B1(net1455),
    .Y(_1265_),
    .A1(_1235_),
    .A2(_1264_));
 sg13g2_nor2_1 _5298_ (.A(net1606),
    .B(_1240_),
    .Y(_1266_));
 sg13g2_a22oi_1 _5299_ (.Y(_0213_),
    .B1(_1265_),
    .B2(_1266_),
    .A2(_3453_),
    .A1(net1605));
 sg13g2_a21oi_1 _5300_ (.A1(net1444),
    .A2(net574),
    .Y(_1267_),
    .B1(_1229_));
 sg13g2_a21oi_1 _5301_ (.A1(net1192),
    .A2(_1232_),
    .Y(_1268_),
    .B1(net1609));
 sg13g2_o21ai_1 _5302_ (.B1(_1268_),
    .Y(_1269_),
    .A1(net1192),
    .A2(_1267_));
 sg13g2_o21ai_1 _5303_ (.B1(_1269_),
    .Y(_1270_),
    .A1(net1733),
    .A2(net804));
 sg13g2_inv_1 _5304_ (.Y(_0214_),
    .A(_1270_));
 sg13g2_and2_1 _5305_ (.A(net1441),
    .B(\s0.data_out[18][6] ),
    .X(_1271_));
 sg13g2_o21ai_1 _5306_ (.B1(net1454),
    .Y(_1272_),
    .A1(_1211_),
    .A2(_1271_));
 sg13g2_nor2_1 _5307_ (.A(net1605),
    .B(_1214_),
    .Y(_1273_));
 sg13g2_a22oi_1 _5308_ (.Y(_0215_),
    .B1(_1272_),
    .B2(_1273_),
    .A2(_3452_),
    .A1(net1606));
 sg13g2_nor2_1 _5309_ (.A(net1197),
    .B(_3457_),
    .Y(_1274_));
 sg13g2_o21ai_1 _5310_ (.B1(net1455),
    .Y(_1275_),
    .A1(_1218_),
    .A2(_1274_));
 sg13g2_nor2_1 _5311_ (.A(net1606),
    .B(_1221_),
    .Y(_1276_));
 sg13g2_a22oi_1 _5312_ (.Y(_0216_),
    .B1(_1275_),
    .B2(_1276_),
    .A2(_3451_),
    .A1(net1606));
 sg13g2_o21ai_1 _5313_ (.B1(net1446),
    .Y(_1277_),
    .A1(net1632),
    .A2(net1432));
 sg13g2_a21oi_1 _5314_ (.A1(net1623),
    .A2(net1436),
    .Y(_1278_),
    .B1(_1277_));
 sg13g2_a21oi_1 _5315_ (.A1(net1624),
    .A2(net1450),
    .Y(_1279_),
    .B1(net1446));
 sg13g2_nor3_1 _5316_ (.A(net826),
    .B(_1278_),
    .C(net404),
    .Y(_1280_));
 sg13g2_or2_1 _5317_ (.X(_1281_),
    .B(net1436),
    .A(net420));
 sg13g2_nor2_1 _5318_ (.A(net1431),
    .B(_1277_),
    .Y(_1282_));
 sg13g2_or2_1 _5319_ (.X(_1283_),
    .B(net1450),
    .A(net420));
 sg13g2_a221oi_1 _5320_ (.B2(net1197),
    .C1(_1282_),
    .B1(_1283_),
    .A1(_1278_),
    .Y(_1284_),
    .A2(_1281_));
 sg13g2_nor3_1 _5321_ (.A(net1609),
    .B(_1280_),
    .C(_1284_),
    .Y(_0217_));
 sg13g2_nor3_1 _5322_ (.A(net1611),
    .B(_1278_),
    .C(net404),
    .Y(_0218_));
 sg13g2_and2_1 _5323_ (.A(net1733),
    .B(net390),
    .X(_0219_));
 sg13g2_nand2_1 _5324_ (.Y(_1285_),
    .A(net1435),
    .B(\s0.data_out[17][2] ));
 sg13g2_o21ai_1 _5325_ (.B1(_1285_),
    .Y(_1286_),
    .A1(net1435),
    .A2(_3461_));
 sg13g2_nor2b_1 _5326_ (.A(net1430),
    .B_N(net1342),
    .Y(_1287_));
 sg13g2_a21oi_1 _5327_ (.A1(net1429),
    .A2(_1286_),
    .Y(_1288_),
    .B1(_1287_));
 sg13g2_o21ai_1 _5328_ (.B1(_1177_),
    .Y(_1289_),
    .A1(net1448),
    .A2(_3464_));
 sg13g2_nand2_1 _5329_ (.Y(_1290_),
    .A(net1197),
    .B(_1289_));
 sg13g2_o21ai_1 _5330_ (.B1(_1290_),
    .Y(_1291_),
    .A1(net1197),
    .A2(_1288_));
 sg13g2_nand2_1 _5331_ (.Y(_1292_),
    .A(net1435),
    .B(net823));
 sg13g2_mux2_1 _5332_ (.A0(\s0.data_out[18][1] ),
    .A1(\s0.data_out[17][1] ),
    .S(net1435),
    .X(_1293_));
 sg13g2_nor2b_1 _5333_ (.A(net1428),
    .B_N(net1346),
    .Y(_1294_));
 sg13g2_a21oi_1 _5334_ (.A1(net1428),
    .A2(_1293_),
    .Y(_1295_),
    .B1(_1294_));
 sg13g2_nand2b_1 _5335_ (.Y(_1296_),
    .B(net1440),
    .A_N(_1295_));
 sg13g2_o21ai_1 _5336_ (.B1(_1185_),
    .Y(_1297_),
    .A1(net1447),
    .A2(_3465_));
 sg13g2_nand2_1 _5337_ (.Y(_1298_),
    .A(net1196),
    .B(_1297_));
 sg13g2_nand3_1 _5338_ (.B(_1296_),
    .C(_1298_),
    .A(net1696),
    .Y(_1299_));
 sg13g2_mux2_1 _5339_ (.A0(\s0.data_out[18][0] ),
    .A1(\s0.data_out[17][0] ),
    .S(net1435),
    .X(_1300_));
 sg13g2_nor2b_1 _5340_ (.A(net1428),
    .B_N(net1350),
    .Y(_1301_));
 sg13g2_a21oi_1 _5341_ (.A1(net1428),
    .A2(_1300_),
    .Y(_1302_),
    .B1(_1301_));
 sg13g2_mux2_1 _5342_ (.A0(\s0.data_out[17][0] ),
    .A1(\s0.data_out[18][0] ),
    .S(net1447),
    .X(_1303_));
 sg13g2_nand2_1 _5343_ (.Y(_1304_),
    .A(net1196),
    .B(_1303_));
 sg13g2_o21ai_1 _5344_ (.B1(_1304_),
    .Y(_1305_),
    .A1(net1196),
    .A2(_1302_));
 sg13g2_and2_1 _5345_ (.A(net1559),
    .B(_1305_),
    .X(_1306_));
 sg13g2_a21oi_1 _5346_ (.A1(_1296_),
    .A2(_1298_),
    .Y(_1307_),
    .B1(net1696));
 sg13g2_a221oi_1 _5347_ (.B2(_1306_),
    .C1(_1307_),
    .B1(_1299_),
    .A1(net1562),
    .Y(_1308_),
    .A2(_1291_));
 sg13g2_nand2_1 _5348_ (.Y(_1309_),
    .A(net1435),
    .B(net819));
 sg13g2_mux2_1 _5349_ (.A0(\s0.data_out[18][3] ),
    .A1(\s0.data_out[17][3] ),
    .S(net1439),
    .X(_1310_));
 sg13g2_nor2b_1 _5350_ (.A(net1430),
    .B_N(net1339),
    .Y(_1311_));
 sg13g2_a21o_1 _5351_ (.A2(_1310_),
    .A1(net1430),
    .B1(_1311_),
    .X(_1312_));
 sg13g2_nand2b_1 _5352_ (.Y(_1313_),
    .B(\s0.data_out[17][3] ),
    .A_N(net1448));
 sg13g2_a21oi_1 _5353_ (.A1(_1200_),
    .A2(_1313_),
    .Y(_1314_),
    .B1(net1443));
 sg13g2_a21oi_1 _5354_ (.A1(net1442),
    .A2(_1312_),
    .Y(_1315_),
    .B1(_1314_));
 sg13g2_nand2_1 _5355_ (.Y(_1316_),
    .A(net1680),
    .B(_1315_));
 sg13g2_o21ai_1 _5356_ (.B1(_1316_),
    .Y(_1317_),
    .A1(net1562),
    .A2(_1291_));
 sg13g2_nand2_1 _5357_ (.Y(_1318_),
    .A(net1436),
    .B(net638));
 sg13g2_mux2_1 _5358_ (.A0(\s0.data_out[18][6] ),
    .A1(\s0.data_out[17][6] ),
    .S(net1436),
    .X(_1319_));
 sg13g2_nor2b_1 _5359_ (.A(net1432),
    .B_N(net1328),
    .Y(_1320_));
 sg13g2_a21o_1 _5360_ (.A2(_1319_),
    .A1(net1432),
    .B1(_1320_),
    .X(_1321_));
 sg13g2_nand2b_1 _5361_ (.Y(_1322_),
    .B(\s0.data_out[17][6] ),
    .A_N(net1449));
 sg13g2_a21oi_1 _5362_ (.A1(_1209_),
    .A2(_1322_),
    .Y(_1323_),
    .B1(net1445));
 sg13g2_a21oi_1 _5363_ (.A1(net1445),
    .A2(_1321_),
    .Y(_1324_),
    .B1(_1323_));
 sg13g2_nand2_1 _5364_ (.Y(_1325_),
    .A(net1436),
    .B(net582));
 sg13g2_mux2_1 _5365_ (.A0(\s0.data_out[18][7] ),
    .A1(\s0.data_out[17][7] ),
    .S(net1436),
    .X(_1326_));
 sg13g2_nor2b_1 _5366_ (.A(net1432),
    .B_N(net1323),
    .Y(_1327_));
 sg13g2_a21o_1 _5367_ (.A2(_1326_),
    .A1(net1432),
    .B1(_1327_),
    .X(_1328_));
 sg13g2_nand2b_1 _5368_ (.Y(_1329_),
    .B(net582),
    .A_N(net1450));
 sg13g2_a21oi_1 _5369_ (.A1(_1216_),
    .A2(_1329_),
    .Y(_1330_),
    .B1(net1445));
 sg13g2_a21oi_1 _5370_ (.A1(net1446),
    .A2(_1328_),
    .Y(_1331_),
    .B1(_1330_));
 sg13g2_a22oi_1 _5371_ (.Y(_1332_),
    .B1(_1331_),
    .B2(net1643),
    .A2(_1324_),
    .A1(net1653));
 sg13g2_nor2_1 _5372_ (.A(net1653),
    .B(_1324_),
    .Y(_1333_));
 sg13g2_or2_1 _5373_ (.X(_1334_),
    .B(_1331_),
    .A(net1643));
 sg13g2_nand3b_1 _5374_ (.B(_1334_),
    .C(_1332_),
    .Y(_1335_),
    .A_N(_1333_));
 sg13g2_nand2_1 _5375_ (.Y(_1336_),
    .A(net1438),
    .B(\s0.data_out[17][4] ));
 sg13g2_o21ai_1 _5376_ (.B1(_1336_),
    .Y(_1337_),
    .A1(net1438),
    .A2(_3459_));
 sg13g2_nor2b_1 _5377_ (.A(net1431),
    .B_N(net1337),
    .Y(_1338_));
 sg13g2_a21o_1 _5378_ (.A2(_1337_),
    .A1(net1431),
    .B1(_1338_),
    .X(_1339_));
 sg13g2_nand2b_1 _5379_ (.Y(_1340_),
    .B(\s0.data_out[17][4] ),
    .A_N(net1449));
 sg13g2_a21oi_1 _5380_ (.A1(_1236_),
    .A2(_1340_),
    .Y(_1341_),
    .B1(net1444));
 sg13g2_a21oi_1 _5381_ (.A1(net1445),
    .A2(_1339_),
    .Y(_1342_),
    .B1(_1341_));
 sg13g2_nand2_1 _5382_ (.Y(_1343_),
    .A(net1436),
    .B(\s0.data_out[17][5] ));
 sg13g2_mux2_1 _5383_ (.A0(\s0.data_out[18][5] ),
    .A1(\s0.data_out[17][5] ),
    .S(net1438),
    .X(_1344_));
 sg13g2_nor2b_1 _5384_ (.A(net1431),
    .B_N(net1333),
    .Y(_1345_));
 sg13g2_a21o_1 _5385_ (.A2(_1344_),
    .A1(net1431),
    .B1(_1345_),
    .X(_1346_));
 sg13g2_nand2b_1 _5386_ (.Y(_1347_),
    .B(\s0.data_out[17][5] ),
    .A_N(net1449));
 sg13g2_a21oi_1 _5387_ (.A1(_1227_),
    .A2(_1347_),
    .Y(_1348_),
    .B1(net1444));
 sg13g2_a21oi_1 _5388_ (.A1(net1444),
    .A2(_1346_),
    .Y(_1349_),
    .B1(_1348_));
 sg13g2_a22oi_1 _5389_ (.Y(_1350_),
    .B1(_1349_),
    .B2(net1661),
    .A2(_1342_),
    .A1(net1672));
 sg13g2_nor2_1 _5390_ (.A(net1663),
    .B(_1349_),
    .Y(_1351_));
 sg13g2_nor2_1 _5391_ (.A(net1680),
    .B(_1315_),
    .Y(_1352_));
 sg13g2_nor2_1 _5392_ (.A(_1351_),
    .B(_1352_),
    .Y(_1353_));
 sg13g2_o21ai_1 _5393_ (.B1(_1350_),
    .Y(_1354_),
    .A1(net1672),
    .A2(_1342_));
 sg13g2_o21ai_1 _5394_ (.B1(_1353_),
    .Y(_1355_),
    .A1(_1308_),
    .A2(_1317_));
 sg13g2_or3_1 _5395_ (.A(_1335_),
    .B(_1354_),
    .C(_1355_),
    .X(_1356_));
 sg13g2_nor3_1 _5396_ (.A(_1335_),
    .B(_1350_),
    .C(_1351_),
    .Y(_1357_));
 sg13g2_nor2b_1 _5397_ (.A(_1332_),
    .B_N(_1334_),
    .Y(_1358_));
 sg13g2_nor4_1 _5398_ (.A(_1278_),
    .B(_1279_),
    .C(_1357_),
    .D(_1358_),
    .Y(_1359_));
 sg13g2_or2_1 _5399_ (.X(_1360_),
    .B(net1557),
    .A(net381));
 sg13g2_a21oi_1 _5400_ (.A1(_1356_),
    .A2(net405),
    .Y(_0220_),
    .B1(_1360_));
 sg13g2_a21oi_1 _5401_ (.A1(net1428),
    .A2(net780),
    .Y(_1361_),
    .B1(_1301_));
 sg13g2_a21oi_1 _5402_ (.A1(net1196),
    .A2(_1303_),
    .Y(_1362_),
    .B1(net1608));
 sg13g2_o21ai_1 _5403_ (.B1(_1362_),
    .Y(_1363_),
    .A1(net1196),
    .A2(_1361_));
 sg13g2_o21ai_1 _5404_ (.B1(_1363_),
    .Y(_1364_),
    .A1(net1732),
    .A2(net787));
 sg13g2_inv_1 _5405_ (.Y(_0221_),
    .A(_1364_));
 sg13g2_a21oi_1 _5406_ (.A1(net1428),
    .A2(\s0.data_out[17][1] ),
    .Y(_1365_),
    .B1(_1294_));
 sg13g2_a21oi_1 _5407_ (.A1(net1196),
    .A2(_1297_),
    .Y(_1366_),
    .B1(net1607));
 sg13g2_o21ai_1 _5408_ (.B1(_1366_),
    .Y(_1367_),
    .A1(net1196),
    .A2(_1365_));
 sg13g2_o21ai_1 _5409_ (.B1(_1367_),
    .Y(_1368_),
    .A1(net1732),
    .A2(net798));
 sg13g2_inv_1 _5410_ (.Y(_0222_),
    .A(net799));
 sg13g2_nor2_1 _5411_ (.A(net1198),
    .B(_3464_),
    .Y(_1369_));
 sg13g2_o21ai_1 _5412_ (.B1(net1442),
    .Y(_1370_),
    .A1(_1287_),
    .A2(_1369_));
 sg13g2_nand3_1 _5413_ (.B(_1290_),
    .C(_1370_),
    .A(net1732),
    .Y(_1371_));
 sg13g2_o21ai_1 _5414_ (.B1(_1371_),
    .Y(_1372_),
    .A1(net1732),
    .A2(net627));
 sg13g2_inv_1 _5415_ (.Y(_0223_),
    .A(net628));
 sg13g2_nor2_1 _5416_ (.A(net1198),
    .B(_3463_),
    .Y(_1373_));
 sg13g2_o21ai_1 _5417_ (.B1(net1442),
    .Y(_1374_),
    .A1(_1311_),
    .A2(_1373_));
 sg13g2_nor2_1 _5418_ (.A(net1609),
    .B(_1314_),
    .Y(_1375_));
 sg13g2_a22oi_1 _5419_ (.Y(_0224_),
    .B1(_1374_),
    .B2(_1375_),
    .A2(_3460_),
    .A1(net1609));
 sg13g2_and2_1 _5420_ (.A(net1431),
    .B(\s0.data_out[17][4] ),
    .X(_1376_));
 sg13g2_o21ai_1 _5421_ (.B1(net1444),
    .Y(_1377_),
    .A1(_1338_),
    .A2(_1376_));
 sg13g2_nor2_1 _5422_ (.A(net1609),
    .B(_1341_),
    .Y(_1378_));
 sg13g2_a22oi_1 _5423_ (.Y(_0225_),
    .B1(_1377_),
    .B2(_1378_),
    .A2(_3459_),
    .A1(net1609));
 sg13g2_and2_1 _5424_ (.A(net1431),
    .B(\s0.data_out[17][5] ),
    .X(_1379_));
 sg13g2_o21ai_1 _5425_ (.B1(net1444),
    .Y(_1380_),
    .A1(_1345_),
    .A2(_1379_));
 sg13g2_nor2_1 _5426_ (.A(net1609),
    .B(_1348_),
    .Y(_1381_));
 sg13g2_a22oi_1 _5427_ (.Y(_0226_),
    .B1(_1380_),
    .B2(_1381_),
    .A2(_3458_),
    .A1(net1609));
 sg13g2_and2_1 _5428_ (.A(net1432),
    .B(\s0.data_out[17][6] ),
    .X(_1382_));
 sg13g2_o21ai_1 _5429_ (.B1(net1445),
    .Y(_1383_),
    .A1(_1320_),
    .A2(_1382_));
 sg13g2_nand3b_1 _5430_ (.B(_1383_),
    .C(net1733),
    .Y(_1384_),
    .A_N(_1323_));
 sg13g2_o21ai_1 _5431_ (.B1(_1384_),
    .Y(_1385_),
    .A1(net1733),
    .A2(net808));
 sg13g2_inv_1 _5432_ (.Y(_0227_),
    .A(net809));
 sg13g2_nor2_1 _5433_ (.A(net1199),
    .B(_3462_),
    .Y(_1386_));
 sg13g2_o21ai_1 _5434_ (.B1(net1445),
    .Y(_1387_),
    .A1(_1327_),
    .A2(_1386_));
 sg13g2_nor2_1 _5435_ (.A(net1611),
    .B(_1330_),
    .Y(_1388_));
 sg13g2_a22oi_1 _5436_ (.Y(_0228_),
    .B1(_1387_),
    .B2(_1388_),
    .A2(_3457_),
    .A1(net1611));
 sg13g2_o21ai_1 _5437_ (.B1(net1433),
    .Y(_1389_),
    .A1(net1632),
    .A2(net1420));
 sg13g2_nor2_1 _5438_ (.A(net1632),
    .B(_3376_),
    .Y(_1390_));
 sg13g2_nor2_1 _5439_ (.A(_1389_),
    .B(_1390_),
    .Y(_1391_));
 sg13g2_a21oi_1 _5440_ (.A1(net1623),
    .A2(net1437),
    .Y(_1392_),
    .B1(net1433));
 sg13g2_nor2_1 _5441_ (.A(_1391_),
    .B(_1392_),
    .Y(_1393_));
 sg13g2_o21ai_1 _5442_ (.B1(_1391_),
    .Y(_1394_),
    .A1(\s0.was_valid_out[16] [0]),
    .A2(net1425));
 sg13g2_nor2_1 _5443_ (.A(net1420),
    .B(_1389_),
    .Y(_1395_));
 sg13g2_o21ai_1 _5444_ (.B1(net1199),
    .Y(_1396_),
    .A1(\s0.was_valid_out[16] [0]),
    .A2(net1436));
 sg13g2_nand2_1 _5445_ (.Y(_1397_),
    .A(_1394_),
    .B(_1396_));
 sg13g2_o21ai_1 _5446_ (.B1(net1734),
    .Y(_1398_),
    .A1(_1395_),
    .A2(_1397_));
 sg13g2_a21oi_1 _5447_ (.A1(_3366_),
    .A2(_1393_),
    .Y(_0229_),
    .B1(_1398_));
 sg13g2_nor3_1 _5448_ (.A(net1610),
    .B(_1391_),
    .C(_1392_),
    .Y(_0230_));
 sg13g2_and2_1 _5449_ (.A(net1736),
    .B(net389),
    .X(_0231_));
 sg13g2_nand2_1 _5450_ (.Y(_1399_),
    .A(net1424),
    .B(net484));
 sg13g2_o21ai_1 _5451_ (.B1(_1399_),
    .Y(_1400_),
    .A1(net1424),
    .A2(_3465_));
 sg13g2_nor2b_1 _5452_ (.A(net1415),
    .B_N(net1346),
    .Y(_1401_));
 sg13g2_a21o_1 _5453_ (.A2(_1400_),
    .A1(net1415),
    .B1(_1401_),
    .X(_1402_));
 sg13g2_nand2b_1 _5454_ (.Y(_1403_),
    .B(net484),
    .A_N(net1435));
 sg13g2_a21oi_1 _5455_ (.A1(_1292_),
    .A2(_1403_),
    .Y(_1404_),
    .B1(net1428));
 sg13g2_a21oi_1 _5456_ (.A1(net1429),
    .A2(_1402_),
    .Y(_1405_),
    .B1(_1404_));
 sg13g2_mux2_1 _5457_ (.A0(\s0.data_out[16][0] ),
    .A1(\s0.data_out[17][0] ),
    .S(net1435),
    .X(_1406_));
 sg13g2_nand2_1 _5458_ (.Y(_1407_),
    .A(net1198),
    .B(_1406_));
 sg13g2_nor2b_1 _5459_ (.A(net1415),
    .B_N(net1350),
    .Y(_1408_));
 sg13g2_mux2_1 _5460_ (.A0(\s0.data_out[17][0] ),
    .A1(\s0.data_out[16][0] ),
    .S(net1424),
    .X(_1409_));
 sg13g2_a21oi_1 _5461_ (.A1(net1415),
    .A2(_1409_),
    .Y(_1410_),
    .B1(_1408_));
 sg13g2_nand2b_1 _5462_ (.Y(_1411_),
    .B(net1429),
    .A_N(_1410_));
 sg13g2_a221oi_1 _5463_ (.B2(_1411_),
    .C1(net1701),
    .B1(_1407_),
    .A1(net1695),
    .Y(_1412_),
    .A2(_1405_));
 sg13g2_nand2_1 _5464_ (.Y(_1413_),
    .A(net1427),
    .B(net564));
 sg13g2_o21ai_1 _5465_ (.B1(_1413_),
    .Y(_1414_),
    .A1(net1427),
    .A2(_3464_));
 sg13g2_nor2b_1 _5466_ (.A(net1415),
    .B_N(net1342),
    .Y(_1415_));
 sg13g2_a21oi_1 _5467_ (.A1(net1416),
    .A2(_1414_),
    .Y(_1416_),
    .B1(_1415_));
 sg13g2_o21ai_1 _5468_ (.B1(_1285_),
    .Y(_1417_),
    .A1(net1439),
    .A2(_3470_));
 sg13g2_nand2_1 _5469_ (.Y(_1418_),
    .A(net1198),
    .B(_1417_));
 sg13g2_o21ai_1 _5470_ (.B1(_1418_),
    .Y(_1419_),
    .A1(net1198),
    .A2(_1416_));
 sg13g2_or2_1 _5471_ (.X(_1420_),
    .B(_1419_),
    .A(net1562));
 sg13g2_xnor2_1 _5472_ (.Y(_1421_),
    .A(net1562),
    .B(_1419_));
 sg13g2_nor2_1 _5473_ (.A(net1695),
    .B(_1405_),
    .Y(_1422_));
 sg13g2_nand2_1 _5474_ (.Y(_1423_),
    .A(net1424),
    .B(net471));
 sg13g2_o21ai_1 _5475_ (.B1(_1423_),
    .Y(_1424_),
    .A1(net1424),
    .A2(_3463_));
 sg13g2_nor2_1 _5476_ (.A(net1416),
    .B(net1161),
    .Y(_1425_));
 sg13g2_a21o_1 _5477_ (.A2(_1424_),
    .A1(net1416),
    .B1(_1425_),
    .X(_1426_));
 sg13g2_nand2b_1 _5478_ (.Y(_1427_),
    .B(net471),
    .A_N(net1439));
 sg13g2_a21oi_1 _5479_ (.A1(_1309_),
    .A2(_1427_),
    .Y(_1428_),
    .B1(net1430));
 sg13g2_a21oi_1 _5480_ (.A1(net1430),
    .A2(_1426_),
    .Y(_1429_),
    .B1(_1428_));
 sg13g2_nor2_1 _5481_ (.A(net1680),
    .B(_1429_),
    .Y(_1430_));
 sg13g2_nor4_1 _5482_ (.A(_1412_),
    .B(_1421_),
    .C(_1422_),
    .D(_1430_),
    .Y(_1431_));
 sg13g2_nand2_1 _5483_ (.Y(_1432_),
    .A(net1680),
    .B(_1429_));
 sg13g2_o21ai_1 _5484_ (.B1(_1432_),
    .Y(_1433_),
    .A1(_1420_),
    .A2(_1430_));
 sg13g2_nand2_1 _5485_ (.Y(_1434_),
    .A(net1426),
    .B(net538));
 sg13g2_mux2_1 _5486_ (.A0(\s0.data_out[17][7] ),
    .A1(\s0.data_out[16][7] ),
    .S(net1425),
    .X(_1435_));
 sg13g2_nor2b_1 _5487_ (.A(net1420),
    .B_N(net1322),
    .Y(_1436_));
 sg13g2_a21o_1 _5488_ (.A2(_1435_),
    .A1(net1419),
    .B1(_1436_),
    .X(_1437_));
 sg13g2_nand2b_1 _5489_ (.Y(_1438_),
    .B(net538),
    .A_N(net1437));
 sg13g2_a21oi_1 _5490_ (.A1(_1325_),
    .A2(_1438_),
    .Y(_1439_),
    .B1(net1432));
 sg13g2_a21oi_1 _5491_ (.A1(net1432),
    .A2(_1437_),
    .Y(_1440_),
    .B1(_1439_));
 sg13g2_nand2_1 _5492_ (.Y(_1441_),
    .A(net1425),
    .B(net752));
 sg13g2_mux2_1 _5493_ (.A0(\s0.data_out[17][6] ),
    .A1(\s0.data_out[16][6] ),
    .S(net1425),
    .X(_1442_));
 sg13g2_nor2b_1 _5494_ (.A(net1420),
    .B_N(net1327),
    .Y(_1443_));
 sg13g2_a21o_1 _5495_ (.A2(_1442_),
    .A1(net1419),
    .B1(_1443_),
    .X(_1444_));
 sg13g2_nand2b_1 _5496_ (.Y(_1445_),
    .B(\s0.data_out[16][6] ),
    .A_N(net1437));
 sg13g2_a21oi_1 _5497_ (.A1(_1318_),
    .A2(_1445_),
    .Y(_1446_),
    .B1(net1433));
 sg13g2_a21oi_1 _5498_ (.A1(net1433),
    .A2(_1444_),
    .Y(_1447_),
    .B1(_1446_));
 sg13g2_a22oi_1 _5499_ (.Y(_1448_),
    .B1(_1447_),
    .B2(net1653),
    .A2(_1440_),
    .A1(net1643));
 sg13g2_nor2_1 _5500_ (.A(net1653),
    .B(_1447_),
    .Y(_1449_));
 sg13g2_or2_1 _5501_ (.X(_1450_),
    .B(_1440_),
    .A(net1643));
 sg13g2_inv_1 _5502_ (.Y(_1451_),
    .A(_1450_));
 sg13g2_nand3b_1 _5503_ (.B(_1450_),
    .C(_1448_),
    .Y(_1452_),
    .A_N(_1449_));
 sg13g2_nand2_1 _5504_ (.Y(_1453_),
    .A(net1426),
    .B(net465));
 sg13g2_mux2_1 _5505_ (.A0(\s0.data_out[17][5] ),
    .A1(\s0.data_out[16][5] ),
    .S(net1426),
    .X(_1454_));
 sg13g2_nor2b_1 _5506_ (.A(net1419),
    .B_N(net1332),
    .Y(_1455_));
 sg13g2_a21oi_1 _5507_ (.A1(net1419),
    .A2(_1454_),
    .Y(_1456_),
    .B1(_1455_));
 sg13g2_nand2b_1 _5508_ (.Y(_1457_),
    .B(net1431),
    .A_N(_1456_));
 sg13g2_o21ai_1 _5509_ (.B1(_1343_),
    .Y(_1458_),
    .A1(net1437),
    .A2(_3467_));
 sg13g2_nand2_1 _5510_ (.Y(_1459_),
    .A(_3375_),
    .B(_1458_));
 sg13g2_nand3_1 _5511_ (.B(_1457_),
    .C(_1459_),
    .A(net1661),
    .Y(_1460_));
 sg13g2_nor2b_1 _5512_ (.A(net1419),
    .B_N(net1337),
    .Y(_1461_));
 sg13g2_nand2_1 _5513_ (.Y(_1462_),
    .A(net1426),
    .B(net716));
 sg13g2_mux2_1 _5514_ (.A0(\s0.data_out[17][4] ),
    .A1(\s0.data_out[16][4] ),
    .S(net1426),
    .X(_1463_));
 sg13g2_a21oi_1 _5515_ (.A1(net1419),
    .A2(_1463_),
    .Y(_1464_),
    .B1(_1461_));
 sg13g2_nand2b_1 _5516_ (.Y(_1465_),
    .B(net1434),
    .A_N(_1464_));
 sg13g2_o21ai_1 _5517_ (.B1(_1336_),
    .Y(_1466_),
    .A1(net1438),
    .A2(_3468_));
 sg13g2_nand2_1 _5518_ (.Y(_1467_),
    .A(net1199),
    .B(_1466_));
 sg13g2_nand3_1 _5519_ (.B(_1465_),
    .C(_1467_),
    .A(net1671),
    .Y(_1468_));
 sg13g2_nand2_1 _5520_ (.Y(_1469_),
    .A(_1460_),
    .B(_1468_));
 sg13g2_a21oi_1 _5521_ (.A1(_1457_),
    .A2(_1459_),
    .Y(_1470_),
    .B1(net1661));
 sg13g2_inv_1 _5522_ (.Y(_1471_),
    .A(_1470_));
 sg13g2_a21oi_1 _5523_ (.A1(_1465_),
    .A2(_1467_),
    .Y(_1472_),
    .B1(net1671));
 sg13g2_nor4_1 _5524_ (.A(_1452_),
    .B(_1469_),
    .C(_1470_),
    .D(_1472_),
    .Y(_1473_));
 sg13g2_o21ai_1 _5525_ (.B1(_1473_),
    .Y(_1474_),
    .A1(_1431_),
    .A2(_1433_));
 sg13g2_a21oi_1 _5526_ (.A1(_1460_),
    .A2(_1468_),
    .Y(_1475_),
    .B1(_1452_));
 sg13g2_o21ai_1 _5527_ (.B1(_1393_),
    .Y(_1476_),
    .A1(_1448_),
    .A2(_1451_));
 sg13g2_a21oi_1 _5528_ (.A1(_1471_),
    .A2(_1475_),
    .Y(_1477_),
    .B1(_1476_));
 sg13g2_or2_1 _5529_ (.X(_1478_),
    .B(net1557),
    .A(net390));
 sg13g2_a21oi_1 _5530_ (.A1(_1474_),
    .A2(_1477_),
    .Y(_0232_),
    .B1(_1478_));
 sg13g2_a21oi_1 _5531_ (.A1(net1415),
    .A2(net653),
    .Y(_1479_),
    .B1(_1408_));
 sg13g2_a21oi_1 _5532_ (.A1(net1198),
    .A2(_1406_),
    .Y(_1480_),
    .B1(net1608));
 sg13g2_o21ai_1 _5533_ (.B1(_1480_),
    .Y(_1481_),
    .A1(net1198),
    .A2(_1479_));
 sg13g2_o21ai_1 _5534_ (.B1(_1481_),
    .Y(_1482_),
    .A1(net1732),
    .A2(net780));
 sg13g2_inv_1 _5535_ (.Y(_0233_),
    .A(_1482_));
 sg13g2_and2_1 _5536_ (.A(net1415),
    .B(net484),
    .X(_1483_));
 sg13g2_o21ai_1 _5537_ (.B1(net1428),
    .Y(_1484_),
    .A1(_1401_),
    .A2(_1483_));
 sg13g2_nor2_1 _5538_ (.A(net1607),
    .B(_1404_),
    .Y(_1485_));
 sg13g2_a22oi_1 _5539_ (.Y(_0234_),
    .B1(_1484_),
    .B2(_1485_),
    .A2(_3465_),
    .A1(net1607));
 sg13g2_a21oi_1 _5540_ (.A1(net1415),
    .A2(\s0.data_out[16][2] ),
    .Y(_1486_),
    .B1(_1415_));
 sg13g2_a21oi_1 _5541_ (.A1(net1198),
    .A2(_1417_),
    .Y(_1487_),
    .B1(net1607));
 sg13g2_o21ai_1 _5542_ (.B1(_1487_),
    .Y(_1488_),
    .A1(net1199),
    .A2(_1486_));
 sg13g2_o21ai_1 _5543_ (.B1(_1488_),
    .Y(_1489_),
    .A1(net1731),
    .A2(net530));
 sg13g2_inv_1 _5544_ (.Y(_0235_),
    .A(net531));
 sg13g2_and2_1 _5545_ (.A(net1416),
    .B(net471),
    .X(_1490_));
 sg13g2_o21ai_1 _5546_ (.B1(net1430),
    .Y(_1491_),
    .A1(_1425_),
    .A2(_1490_));
 sg13g2_nor2_1 _5547_ (.A(net1610),
    .B(_1428_),
    .Y(_1492_));
 sg13g2_a22oi_1 _5548_ (.Y(_0236_),
    .B1(_1491_),
    .B2(_1492_),
    .A2(_3463_),
    .A1(net1610));
 sg13g2_a21oi_1 _5549_ (.A1(net1419),
    .A2(\s0.data_out[16][4] ),
    .Y(_1493_),
    .B1(_1461_));
 sg13g2_a21oi_1 _5550_ (.A1(_3375_),
    .A2(_1466_),
    .Y(_1494_),
    .B1(net1610));
 sg13g2_o21ai_1 _5551_ (.B1(_1494_),
    .Y(_1495_),
    .A1(net1199),
    .A2(_1493_));
 sg13g2_o21ai_1 _5552_ (.B1(_1495_),
    .Y(_1496_),
    .A1(net1734),
    .A2(net681));
 sg13g2_inv_1 _5553_ (.Y(_0237_),
    .A(net682));
 sg13g2_a21oi_1 _5554_ (.A1(net1419),
    .A2(net465),
    .Y(_1497_),
    .B1(_1455_));
 sg13g2_a21oi_1 _5555_ (.A1(net1199),
    .A2(_1458_),
    .Y(_1498_),
    .B1(net1611));
 sg13g2_o21ai_1 _5556_ (.B1(_1498_),
    .Y(_1499_),
    .A1(net1199),
    .A2(_1497_));
 sg13g2_o21ai_1 _5557_ (.B1(_1499_),
    .Y(_1500_),
    .A1(net1734),
    .A2(net708));
 sg13g2_inv_1 _5558_ (.Y(_0238_),
    .A(_1500_));
 sg13g2_and2_1 _5559_ (.A(net1420),
    .B(\s0.data_out[16][6] ),
    .X(_1501_));
 sg13g2_o21ai_1 _5560_ (.B1(net1433),
    .Y(_1502_),
    .A1(_1443_),
    .A2(_1501_));
 sg13g2_nand3b_1 _5561_ (.B(_1502_),
    .C(net1734),
    .Y(_1503_),
    .A_N(_1446_));
 sg13g2_o21ai_1 _5562_ (.B1(_1503_),
    .Y(_1504_),
    .A1(net1734),
    .A2(net638));
 sg13g2_inv_1 _5563_ (.Y(_0239_),
    .A(net639));
 sg13g2_and2_1 _5564_ (.A(net1420),
    .B(net538),
    .X(_1505_));
 sg13g2_o21ai_1 _5565_ (.B1(net1433),
    .Y(_1506_),
    .A1(_1436_),
    .A2(_1505_));
 sg13g2_nor2_1 _5566_ (.A(net1610),
    .B(_1439_),
    .Y(_1507_));
 sg13g2_a22oi_1 _5567_ (.Y(_0240_),
    .B1(_1506_),
    .B2(_1507_),
    .A2(_3462_),
    .A1(net1610));
 sg13g2_o21ai_1 _5568_ (.B1(net1421),
    .Y(_1508_),
    .A1(net1632),
    .A2(net1408));
 sg13g2_nand2_1 _5569_ (.Y(_1509_),
    .A(net1623),
    .B(net1414));
 sg13g2_nand2b_1 _5570_ (.Y(_1510_),
    .B(_1509_),
    .A_N(_1508_));
 sg13g2_o21ai_1 _5571_ (.B1(_1510_),
    .Y(_1511_),
    .A1(net1421),
    .A2(_1390_));
 sg13g2_nor2_1 _5572_ (.A(net398),
    .B(net1414),
    .Y(_1512_));
 sg13g2_or2_1 _5573_ (.X(_1513_),
    .B(_1512_),
    .A(_1510_));
 sg13g2_nor2_1 _5574_ (.A(net1407),
    .B(_1508_),
    .Y(_1514_));
 sg13g2_a21oi_1 _5575_ (.A1(_3365_),
    .A2(_3376_),
    .Y(_1515_),
    .B1(net1422));
 sg13g2_nor2_1 _5576_ (.A(_1514_),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_o21ai_1 _5577_ (.B1(net1733),
    .Y(_1517_),
    .A1(net616),
    .A2(_1511_));
 sg13g2_a21oi_1 _5578_ (.A1(_1513_),
    .A2(_1516_),
    .Y(_0241_),
    .B1(_1517_));
 sg13g2_nor2_1 _5579_ (.A(net1617),
    .B(_1511_),
    .Y(_0242_));
 sg13g2_and2_1 _5580_ (.A(net1737),
    .B(net394),
    .X(_0243_));
 sg13g2_nand2_1 _5581_ (.Y(_1518_),
    .A(net1411),
    .B(net585));
 sg13g2_mux2_1 _5582_ (.A0(\s0.data_out[16][2] ),
    .A1(\s0.data_out[15][2] ),
    .S(net1411),
    .X(_1519_));
 sg13g2_nor2b_1 _5583_ (.A(net1404),
    .B_N(net1342),
    .Y(_1520_));
 sg13g2_a21o_1 _5584_ (.A2(_1519_),
    .A1(net1405),
    .B1(_1520_),
    .X(_1521_));
 sg13g2_nand2b_1 _5585_ (.Y(_1522_),
    .B(\s0.data_out[15][2] ),
    .A_N(net1427));
 sg13g2_a21oi_1 _5586_ (.A1(_1413_),
    .A2(_1522_),
    .Y(_1523_),
    .B1(net1416));
 sg13g2_a21oi_1 _5587_ (.A1(net1417),
    .A2(_1521_),
    .Y(_1524_),
    .B1(_1523_));
 sg13g2_nor2_1 _5588_ (.A(net1686),
    .B(_1524_),
    .Y(_1525_));
 sg13g2_nand2_1 _5589_ (.Y(_1526_),
    .A(net1411),
    .B(net814));
 sg13g2_mux2_1 _5590_ (.A0(\s0.data_out[16][1] ),
    .A1(\s0.data_out[15][1] ),
    .S(net1411),
    .X(_1527_));
 sg13g2_nor2b_1 _5591_ (.A(net1404),
    .B_N(net1346),
    .Y(_1528_));
 sg13g2_a21o_1 _5592_ (.A2(_1527_),
    .A1(net1404),
    .B1(_1528_),
    .X(_1529_));
 sg13g2_nand2b_1 _5593_ (.Y(_1530_),
    .B(\s0.data_out[15][1] ),
    .A_N(net1424));
 sg13g2_a21oi_1 _5594_ (.A1(_1399_),
    .A2(_1530_),
    .Y(_1531_),
    .B1(net1417));
 sg13g2_a21oi_1 _5595_ (.A1(net1417),
    .A2(_1529_),
    .Y(_1532_),
    .B1(_1531_));
 sg13g2_nor2_1 _5596_ (.A(net1695),
    .B(_1532_),
    .Y(_1533_));
 sg13g2_mux2_1 _5597_ (.A0(\s0.data_out[16][0] ),
    .A1(\s0.data_out[15][0] ),
    .S(net1411),
    .X(_1534_));
 sg13g2_nor2b_1 _5598_ (.A(net1404),
    .B_N(net1350),
    .Y(_1535_));
 sg13g2_a21oi_1 _5599_ (.A1(net1404),
    .A2(_1534_),
    .Y(_1536_),
    .B1(_1535_));
 sg13g2_nand2b_1 _5600_ (.Y(_1537_),
    .B(net1417),
    .A_N(_1536_));
 sg13g2_mux2_1 _5601_ (.A0(\s0.data_out[15][0] ),
    .A1(\s0.data_out[16][0] ),
    .S(net1424),
    .X(_1538_));
 sg13g2_nand2b_1 _5602_ (.Y(_1539_),
    .B(_1538_),
    .A_N(net1417));
 sg13g2_a221oi_1 _5603_ (.B2(_1539_),
    .C1(net1701),
    .B1(_1537_),
    .A1(net1695),
    .Y(_1540_),
    .A2(_1532_));
 sg13g2_nor3_1 _5604_ (.A(_1525_),
    .B(_1533_),
    .C(_1540_),
    .Y(_1541_));
 sg13g2_nand2_1 _5605_ (.Y(_1542_),
    .A(net1411),
    .B(net786));
 sg13g2_mux2_1 _5606_ (.A0(\s0.data_out[16][3] ),
    .A1(\s0.data_out[15][3] ),
    .S(net1412),
    .X(_1543_));
 sg13g2_nor2b_1 _5607_ (.A(net1405),
    .B_N(\s0.data_new_delayed[3] ),
    .Y(_1544_));
 sg13g2_a21o_1 _5608_ (.A2(_1543_),
    .A1(net1405),
    .B1(_1544_),
    .X(_1545_));
 sg13g2_nand2b_1 _5609_ (.Y(_1546_),
    .B(\s0.data_out[15][3] ),
    .A_N(net1424));
 sg13g2_a21oi_1 _5610_ (.A1(_1423_),
    .A2(_1546_),
    .Y(_1547_),
    .B1(net1418));
 sg13g2_a21oi_1 _5611_ (.A1(net1418),
    .A2(_1545_),
    .Y(_1548_),
    .B1(_1547_));
 sg13g2_a221oi_1 _5612_ (.B2(net1682),
    .C1(_1541_),
    .B1(_1548_),
    .A1(net1686),
    .Y(_1549_),
    .A2(_1524_));
 sg13g2_nand2_1 _5613_ (.Y(_1550_),
    .A(net1413),
    .B(net578));
 sg13g2_mux2_1 _5614_ (.A0(\s0.data_out[16][7] ),
    .A1(\s0.data_out[15][7] ),
    .S(net1414),
    .X(_1551_));
 sg13g2_nor2b_1 _5615_ (.A(net1407),
    .B_N(net1322),
    .Y(_1552_));
 sg13g2_a21o_1 _5616_ (.A2(_1551_),
    .A1(net1407),
    .B1(_1552_),
    .X(_1553_));
 sg13g2_nand2b_1 _5617_ (.Y(_1554_),
    .B(\s0.data_out[15][7] ),
    .A_N(net1425));
 sg13g2_a21oi_1 _5618_ (.A1(_1434_),
    .A2(_1554_),
    .Y(_1555_),
    .B1(net1421));
 sg13g2_a21oi_1 _5619_ (.A1(net1422),
    .A2(_1553_),
    .Y(_1556_),
    .B1(_1555_));
 sg13g2_nand2_1 _5620_ (.Y(_1557_),
    .A(net1413),
    .B(net842));
 sg13g2_mux2_1 _5621_ (.A0(\s0.data_out[16][6] ),
    .A1(\s0.data_out[15][6] ),
    .S(net1414),
    .X(_1558_));
 sg13g2_nor2b_1 _5622_ (.A(net1407),
    .B_N(net1327),
    .Y(_1559_));
 sg13g2_a21o_1 _5623_ (.A2(_1558_),
    .A1(net1407),
    .B1(_1559_),
    .X(_1560_));
 sg13g2_nand2b_1 _5624_ (.Y(_1561_),
    .B(net841),
    .A_N(net1425));
 sg13g2_a21oi_1 _5625_ (.A1(_1441_),
    .A2(_1561_),
    .Y(_1562_),
    .B1(net1421));
 sg13g2_a21oi_1 _5626_ (.A1(net1421),
    .A2(_1560_),
    .Y(_1563_),
    .B1(_1562_));
 sg13g2_a22oi_1 _5627_ (.Y(_1564_),
    .B1(_1563_),
    .B2(net1652),
    .A2(_1556_),
    .A1(net1642));
 sg13g2_or2_1 _5628_ (.X(_1565_),
    .B(_1556_),
    .A(net1644));
 sg13g2_nor2_1 _5629_ (.A(net1652),
    .B(_1563_),
    .Y(_1566_));
 sg13g2_nand3b_1 _5630_ (.B(_1564_),
    .C(_1565_),
    .Y(_1567_),
    .A_N(_1566_));
 sg13g2_nand2_1 _5631_ (.Y(_1568_),
    .A(net1413),
    .B(\s0.data_out[15][4] ));
 sg13g2_mux2_1 _5632_ (.A0(\s0.data_out[16][4] ),
    .A1(\s0.data_out[15][4] ),
    .S(net1414),
    .X(_1569_));
 sg13g2_nor2b_1 _5633_ (.A(net1408),
    .B_N(net1337),
    .Y(_1570_));
 sg13g2_a21o_1 _5634_ (.A2(_1569_),
    .A1(net1408),
    .B1(_1570_),
    .X(_1571_));
 sg13g2_nand2b_1 _5635_ (.Y(_1572_),
    .B(\s0.data_out[15][4] ),
    .A_N(net1426));
 sg13g2_a21oi_1 _5636_ (.A1(_1462_),
    .A2(_1572_),
    .Y(_1573_),
    .B1(net1422));
 sg13g2_a21oi_1 _5637_ (.A1(net1422),
    .A2(_1571_),
    .Y(_1574_),
    .B1(_1573_));
 sg13g2_nand2_1 _5638_ (.Y(_1575_),
    .A(net1413),
    .B(\s0.data_out[15][5] ));
 sg13g2_mux2_1 _5639_ (.A0(\s0.data_out[16][5] ),
    .A1(\s0.data_out[15][5] ),
    .S(net1414),
    .X(_1576_));
 sg13g2_nor2b_1 _5640_ (.A(net1408),
    .B_N(net1332),
    .Y(_1577_));
 sg13g2_a21o_1 _5641_ (.A2(_1576_),
    .A1(net1407),
    .B1(_1577_),
    .X(_1578_));
 sg13g2_nand2b_1 _5642_ (.Y(_1579_),
    .B(\s0.data_out[15][5] ),
    .A_N(net1425));
 sg13g2_a21oi_1 _5643_ (.A1(_1453_),
    .A2(_1579_),
    .Y(_1580_),
    .B1(net1421));
 sg13g2_a21oi_1 _5644_ (.A1(net1422),
    .A2(_1578_),
    .Y(_1581_),
    .B1(_1580_));
 sg13g2_a22oi_1 _5645_ (.Y(_1582_),
    .B1(_1581_),
    .B2(net1662),
    .A2(_1574_),
    .A1(net1671));
 sg13g2_nor2_1 _5646_ (.A(net1680),
    .B(_1548_),
    .Y(_1583_));
 sg13g2_nor2_1 _5647_ (.A(net1671),
    .B(_1574_),
    .Y(_1584_));
 sg13g2_nor2_1 _5648_ (.A(net1661),
    .B(_1581_),
    .Y(_1585_));
 sg13g2_nor3_1 _5649_ (.A(_1583_),
    .B(_1584_),
    .C(_1585_),
    .Y(_1586_));
 sg13g2_nand2_1 _5650_ (.Y(_1587_),
    .A(_1582_),
    .B(_1586_));
 sg13g2_or3_1 _5651_ (.A(_1549_),
    .B(_1567_),
    .C(_1587_),
    .X(_1588_));
 sg13g2_nor3_1 _5652_ (.A(_1567_),
    .B(_1582_),
    .C(_1585_),
    .Y(_1589_));
 sg13g2_nor2b_1 _5653_ (.A(_1564_),
    .B_N(_1565_),
    .Y(_1590_));
 sg13g2_nor3_1 _5654_ (.A(_1511_),
    .B(_1589_),
    .C(_1590_),
    .Y(_1591_));
 sg13g2_or2_1 _5655_ (.X(_1592_),
    .B(net1557),
    .A(net389));
 sg13g2_a21oi_1 _5656_ (.A1(_1588_),
    .A2(_1591_),
    .Y(_0244_),
    .B1(_1592_));
 sg13g2_and2_1 _5657_ (.A(net1404),
    .B(\s0.data_out[15][0] ),
    .X(_1593_));
 sg13g2_o21ai_1 _5658_ (.B1(net1417),
    .Y(_1594_),
    .A1(_1535_),
    .A2(_1593_));
 sg13g2_nand3_1 _5659_ (.B(_1539_),
    .C(_1594_),
    .A(net1731),
    .Y(_1595_));
 sg13g2_o21ai_1 _5660_ (.B1(_1595_),
    .Y(_1596_),
    .A1(net1731),
    .A2(net653));
 sg13g2_inv_1 _5661_ (.Y(_0245_),
    .A(_1596_));
 sg13g2_nor2_1 _5662_ (.A(net1190),
    .B(_3475_),
    .Y(_1597_));
 sg13g2_o21ai_1 _5663_ (.B1(net1417),
    .Y(_1598_),
    .A1(_1528_),
    .A2(_1597_));
 sg13g2_nor2_1 _5664_ (.A(net1607),
    .B(_1531_),
    .Y(_1599_));
 sg13g2_a22oi_1 _5665_ (.Y(_0246_),
    .B1(_1598_),
    .B2(_1599_),
    .A2(_3471_),
    .A1(net1607));
 sg13g2_nor2_1 _5666_ (.A(net1190),
    .B(_3474_),
    .Y(_1600_));
 sg13g2_o21ai_1 _5667_ (.B1(net1417),
    .Y(_1601_),
    .A1(_1520_),
    .A2(_1600_));
 sg13g2_nor2_1 _5668_ (.A(net1607),
    .B(_1523_),
    .Y(_1602_));
 sg13g2_a22oi_1 _5669_ (.Y(_0247_),
    .B1(_1601_),
    .B2(_1602_),
    .A2(_3470_),
    .A1(net1607));
 sg13g2_nor2_1 _5670_ (.A(net1190),
    .B(_3473_),
    .Y(_1603_));
 sg13g2_o21ai_1 _5671_ (.B1(net1418),
    .Y(_1604_),
    .A1(_1544_),
    .A2(_1603_));
 sg13g2_nor2_1 _5672_ (.A(net1617),
    .B(_1547_),
    .Y(_1605_));
 sg13g2_a22oi_1 _5673_ (.Y(_0248_),
    .B1(_1604_),
    .B2(_1605_),
    .A2(_3469_),
    .A1(net1617));
 sg13g2_and2_1 _5674_ (.A(net1408),
    .B(\s0.data_out[15][4] ),
    .X(_1606_));
 sg13g2_o21ai_1 _5675_ (.B1(net1422),
    .Y(_1607_),
    .A1(_1570_),
    .A2(_1606_));
 sg13g2_nor2_1 _5676_ (.A(net1611),
    .B(_1573_),
    .Y(_1608_));
 sg13g2_a22oi_1 _5677_ (.Y(_0249_),
    .B1(_1607_),
    .B2(_1608_),
    .A2(_3468_),
    .A1(net1610));
 sg13g2_and2_1 _5678_ (.A(net1407),
    .B(net589),
    .X(_1609_));
 sg13g2_o21ai_1 _5679_ (.B1(net1421),
    .Y(_1610_),
    .A1(_1577_),
    .A2(_1609_));
 sg13g2_nor2_1 _5680_ (.A(net1611),
    .B(net466),
    .Y(_1611_));
 sg13g2_a22oi_1 _5681_ (.Y(_0250_),
    .B1(_1610_),
    .B2(_1611_),
    .A2(_3467_),
    .A1(net1610));
 sg13g2_and2_1 _5682_ (.A(net1407),
    .B(\s0.data_out[15][6] ),
    .X(_1612_));
 sg13g2_o21ai_1 _5683_ (.B1(net1421),
    .Y(_1613_),
    .A1(_1559_),
    .A2(_1612_));
 sg13g2_nand3b_1 _5684_ (.B(_1613_),
    .C(net1733),
    .Y(_1614_),
    .A_N(_1562_));
 sg13g2_o21ai_1 _5685_ (.B1(_1614_),
    .Y(_1615_),
    .A1(net1733),
    .A2(net752));
 sg13g2_inv_1 _5686_ (.Y(_0251_),
    .A(_1615_));
 sg13g2_nor2_1 _5687_ (.A(net1189),
    .B(_3472_),
    .Y(_1616_));
 sg13g2_o21ai_1 _5688_ (.B1(net1422),
    .Y(_1617_),
    .A1(_1552_),
    .A2(_1616_));
 sg13g2_nor2_1 _5689_ (.A(net1617),
    .B(_1555_),
    .Y(_1618_));
 sg13g2_a22oi_1 _5690_ (.Y(_0252_),
    .B1(_1617_),
    .B2(_1618_),
    .A2(_3466_),
    .A1(net1618));
 sg13g2_o21ai_1 _5691_ (.B1(net1410),
    .Y(_1619_),
    .A1(net1633),
    .A2(net1399));
 sg13g2_nor2b_1 _5692_ (.A(net1633),
    .B_N(net1402),
    .Y(_1620_));
 sg13g2_nor2_1 _5693_ (.A(_1619_),
    .B(_1620_),
    .Y(_1621_));
 sg13g2_a21oi_1 _5694_ (.A1(net1189),
    .A2(_1509_),
    .Y(_1622_),
    .B1(_1621_));
 sg13g2_o21ai_1 _5695_ (.B1(_1621_),
    .Y(_1623_),
    .A1(\s0.was_valid_out[14] [0]),
    .A2(net1403));
 sg13g2_nor2_1 _5696_ (.A(net1396),
    .B(_1619_),
    .Y(_1624_));
 sg13g2_o21ai_1 _5697_ (.B1(net1189),
    .Y(_1625_),
    .A1(\s0.was_valid_out[14] [0]),
    .A2(net1413));
 sg13g2_nand2_1 _5698_ (.Y(_1626_),
    .A(_1623_),
    .B(_1625_));
 sg13g2_o21ai_1 _5699_ (.B1(net1736),
    .Y(_1627_),
    .A1(_1624_),
    .A2(_1626_));
 sg13g2_a21oi_1 _5700_ (.A1(_3365_),
    .A2(_1622_),
    .Y(_0253_),
    .B1(_1627_));
 sg13g2_and2_1 _5701_ (.A(net1736),
    .B(_1622_),
    .X(_0254_));
 sg13g2_and2_1 _5702_ (.A(net1737),
    .B(net392),
    .X(_0255_));
 sg13g2_nand2_1 _5703_ (.Y(_1628_),
    .A(net1400),
    .B(net729));
 sg13g2_o21ai_1 _5704_ (.B1(_1628_),
    .Y(_1629_),
    .A1(net1400),
    .A2(_3475_));
 sg13g2_nor2b_1 _5705_ (.A(net1393),
    .B_N(\s0.data_new_delayed[1] ),
    .Y(_1630_));
 sg13g2_a21o_1 _5706_ (.A2(_1629_),
    .A1(net1393),
    .B1(_1630_),
    .X(_1631_));
 sg13g2_nand2b_1 _5707_ (.Y(_1632_),
    .B(net729),
    .A_N(net1411));
 sg13g2_a21oi_1 _5708_ (.A1(_1526_),
    .A2(_1632_),
    .Y(_1633_),
    .B1(net1404));
 sg13g2_a21oi_1 _5709_ (.A1(net1405),
    .A2(_1631_),
    .Y(_1634_),
    .B1(_1633_));
 sg13g2_mux2_1 _5710_ (.A0(\s0.data_out[14][0] ),
    .A1(\s0.data_out[15][0] ),
    .S(net1411),
    .X(_1635_));
 sg13g2_nand2_1 _5711_ (.Y(_1636_),
    .A(net1190),
    .B(_1635_));
 sg13g2_nor2b_1 _5712_ (.A(net1393),
    .B_N(net1350),
    .Y(_1637_));
 sg13g2_mux2_1 _5713_ (.A0(\s0.data_out[15][0] ),
    .A1(\s0.data_out[14][0] ),
    .S(net1400),
    .X(_1638_));
 sg13g2_a21oi_1 _5714_ (.A1(net1393),
    .A2(_1638_),
    .Y(_1639_),
    .B1(_1637_));
 sg13g2_nand2b_1 _5715_ (.Y(_1640_),
    .B(net1405),
    .A_N(_1639_));
 sg13g2_a221oi_1 _5716_ (.B2(_1640_),
    .C1(net1702),
    .B1(_1636_),
    .A1(net1697),
    .Y(_1641_),
    .A2(_1634_));
 sg13g2_nand2_1 _5717_ (.Y(_1642_),
    .A(net1400),
    .B(net648));
 sg13g2_o21ai_1 _5718_ (.B1(_1642_),
    .Y(_1643_),
    .A1(net1401),
    .A2(_3474_));
 sg13g2_nor2b_1 _5719_ (.A(net1394),
    .B_N(net1342),
    .Y(_1644_));
 sg13g2_a21oi_1 _5720_ (.A1(net1395),
    .A2(_1643_),
    .Y(_1645_),
    .B1(_1644_));
 sg13g2_o21ai_1 _5721_ (.B1(_1518_),
    .Y(_1646_),
    .A1(net1412),
    .A2(_3480_));
 sg13g2_nand2_1 _5722_ (.Y(_1647_),
    .A(net1190),
    .B(_1646_));
 sg13g2_o21ai_1 _5723_ (.B1(_1647_),
    .Y(_1648_),
    .A1(net1190),
    .A2(_1645_));
 sg13g2_or2_1 _5724_ (.X(_1649_),
    .B(_1648_),
    .A(net1562));
 sg13g2_xnor2_1 _5725_ (.Y(_1650_),
    .A(net1562),
    .B(_1648_));
 sg13g2_nor2_1 _5726_ (.A(net1697),
    .B(_1634_),
    .Y(_1651_));
 sg13g2_nand2_1 _5727_ (.Y(_1652_),
    .A(net1401),
    .B(net730));
 sg13g2_o21ai_1 _5728_ (.B1(_1652_),
    .Y(_1653_),
    .A1(net1401),
    .A2(_3473_));
 sg13g2_nor2_1 _5729_ (.A(net1395),
    .B(net1161),
    .Y(_1654_));
 sg13g2_a21o_1 _5730_ (.A2(_1653_),
    .A1(net1395),
    .B1(_1654_),
    .X(_1655_));
 sg13g2_nand2b_1 _5731_ (.Y(_1656_),
    .B(net730),
    .A_N(net1412));
 sg13g2_a21oi_1 _5732_ (.A1(_1542_),
    .A2(_1656_),
    .Y(_1657_),
    .B1(net1406));
 sg13g2_a21oi_1 _5733_ (.A1(net1406),
    .A2(_1655_),
    .Y(_1658_),
    .B1(_1657_));
 sg13g2_nor2_1 _5734_ (.A(net1681),
    .B(_1658_),
    .Y(_1659_));
 sg13g2_nor4_1 _5735_ (.A(_1641_),
    .B(_1650_),
    .C(_1651_),
    .D(_1659_),
    .Y(_1660_));
 sg13g2_nand2_1 _5736_ (.Y(_1661_),
    .A(net1681),
    .B(_1658_));
 sg13g2_o21ai_1 _5737_ (.B1(_1661_),
    .Y(_1662_),
    .A1(_1649_),
    .A2(_1659_));
 sg13g2_nand2_1 _5738_ (.Y(_1663_),
    .A(net1402),
    .B(net712));
 sg13g2_mux2_1 _5739_ (.A0(\s0.data_out[15][7] ),
    .A1(\s0.data_out[14][7] ),
    .S(net1403),
    .X(_1664_));
 sg13g2_nor2b_1 _5740_ (.A(net1396),
    .B_N(net1322),
    .Y(_1665_));
 sg13g2_a21o_1 _5741_ (.A2(_1664_),
    .A1(net1396),
    .B1(_1665_),
    .X(_1666_));
 sg13g2_nand2b_1 _5742_ (.Y(_1667_),
    .B(\s0.data_out[14][7] ),
    .A_N(net1413));
 sg13g2_a21oi_1 _5743_ (.A1(_1550_),
    .A2(_1667_),
    .Y(_1668_),
    .B1(net1409));
 sg13g2_a21oi_1 _5744_ (.A1(net1409),
    .A2(_1666_),
    .Y(_1669_),
    .B1(_1668_));
 sg13g2_nand2_1 _5745_ (.Y(_1670_),
    .A(net1403),
    .B(net721));
 sg13g2_mux2_1 _5746_ (.A0(\s0.data_out[15][6] ),
    .A1(\s0.data_out[14][6] ),
    .S(net1402),
    .X(_1671_));
 sg13g2_nor2b_1 _5747_ (.A(net1398),
    .B_N(net1327),
    .Y(_1672_));
 sg13g2_a21o_1 _5748_ (.A2(_1671_),
    .A1(net1398),
    .B1(_1672_),
    .X(_1673_));
 sg13g2_nand2b_1 _5749_ (.Y(_1674_),
    .B(\s0.data_out[14][6] ),
    .A_N(net1414));
 sg13g2_a21oi_1 _5750_ (.A1(_1557_),
    .A2(_1674_),
    .Y(_1675_),
    .B1(net1409));
 sg13g2_a21oi_1 _5751_ (.A1(net1409),
    .A2(_1673_),
    .Y(_1676_),
    .B1(_1675_));
 sg13g2_a22oi_1 _5752_ (.Y(_1677_),
    .B1(_1676_),
    .B2(net1652),
    .A2(_1669_),
    .A1(net1644));
 sg13g2_nor2_1 _5753_ (.A(net1652),
    .B(_1676_),
    .Y(_1678_));
 sg13g2_or2_1 _5754_ (.X(_1679_),
    .B(_1669_),
    .A(net1644));
 sg13g2_inv_1 _5755_ (.Y(_1680_),
    .A(_1679_));
 sg13g2_nand3b_1 _5756_ (.B(_1679_),
    .C(_1677_),
    .Y(_1681_),
    .A_N(_1678_));
 sg13g2_nand2_1 _5757_ (.Y(_1682_),
    .A(net1402),
    .B(net783));
 sg13g2_mux2_1 _5758_ (.A0(\s0.data_out[15][5] ),
    .A1(\s0.data_out[14][5] ),
    .S(net1403),
    .X(_1683_));
 sg13g2_nor2b_1 _5759_ (.A(net1396),
    .B_N(net1333),
    .Y(_1684_));
 sg13g2_a21oi_1 _5760_ (.A1(net1399),
    .A2(_1683_),
    .Y(_1685_),
    .B1(_1684_));
 sg13g2_nand2b_1 _5761_ (.Y(_1686_),
    .B(net1409),
    .A_N(_1685_));
 sg13g2_o21ai_1 _5762_ (.B1(_1575_),
    .Y(_1687_),
    .A1(net1413),
    .A2(_3477_));
 sg13g2_nand2_1 _5763_ (.Y(_1688_),
    .A(net1189),
    .B(_1687_));
 sg13g2_nand3_1 _5764_ (.B(_1686_),
    .C(_1688_),
    .A(net1662),
    .Y(_1689_));
 sg13g2_nor2b_1 _5765_ (.A(net1396),
    .B_N(net1337),
    .Y(_1690_));
 sg13g2_nand2_1 _5766_ (.Y(_1691_),
    .A(net1401),
    .B(\s0.data_out[14][4] ));
 sg13g2_mux2_1 _5767_ (.A0(\s0.data_out[15][4] ),
    .A1(\s0.data_out[14][4] ),
    .S(net1403),
    .X(_1692_));
 sg13g2_a21oi_1 _5768_ (.A1(net1396),
    .A2(_1692_),
    .Y(_1693_),
    .B1(_1690_));
 sg13g2_nand2b_1 _5769_ (.Y(_1694_),
    .B(net1409),
    .A_N(_1693_));
 sg13g2_o21ai_1 _5770_ (.B1(_1568_),
    .Y(_1695_),
    .A1(net1413),
    .A2(_3478_));
 sg13g2_nand2_1 _5771_ (.Y(_1696_),
    .A(net1189),
    .B(_1695_));
 sg13g2_nand3_1 _5772_ (.B(_1694_),
    .C(_1696_),
    .A(net1672),
    .Y(_1697_));
 sg13g2_nand2_1 _5773_ (.Y(_1698_),
    .A(_1689_),
    .B(_1697_));
 sg13g2_a21oi_1 _5774_ (.A1(_1686_),
    .A2(_1688_),
    .Y(_1699_),
    .B1(net1662));
 sg13g2_inv_1 _5775_ (.Y(_1700_),
    .A(_1699_));
 sg13g2_a21oi_1 _5776_ (.A1(_1694_),
    .A2(_1696_),
    .Y(_1701_),
    .B1(net1672));
 sg13g2_nor4_1 _5777_ (.A(_1681_),
    .B(_1698_),
    .C(_1699_),
    .D(_1701_),
    .Y(_1702_));
 sg13g2_o21ai_1 _5778_ (.B1(_1702_),
    .Y(_1703_),
    .A1(_1660_),
    .A2(_1662_));
 sg13g2_a21oi_1 _5779_ (.A1(_1689_),
    .A2(_1697_),
    .Y(_1704_),
    .B1(_1681_));
 sg13g2_o21ai_1 _5780_ (.B1(_1622_),
    .Y(_1705_),
    .A1(_1677_),
    .A2(_1680_));
 sg13g2_a21oi_1 _5781_ (.A1(_1700_),
    .A2(_1704_),
    .Y(_1706_),
    .B1(_1705_));
 sg13g2_or2_1 _5782_ (.X(_1707_),
    .B(net1557),
    .A(net394));
 sg13g2_a21oi_1 _5783_ (.A1(_1703_),
    .A2(_1706_),
    .Y(_0256_),
    .B1(_1707_));
 sg13g2_and2_1 _5784_ (.A(net1393),
    .B(\s0.data_out[14][0] ),
    .X(_1708_));
 sg13g2_o21ai_1 _5785_ (.B1(net1405),
    .Y(_1709_),
    .A1(_1637_),
    .A2(_1708_));
 sg13g2_nand3_1 _5786_ (.B(_1636_),
    .C(_1709_),
    .A(net1738),
    .Y(_1710_));
 sg13g2_o21ai_1 _5787_ (.B1(_1710_),
    .Y(_1711_),
    .A1(net1738),
    .A2(net621));
 sg13g2_inv_1 _5788_ (.Y(_0257_),
    .A(_1711_));
 sg13g2_nor2_1 _5789_ (.A(net1188),
    .B(_3481_),
    .Y(_1712_));
 sg13g2_o21ai_1 _5790_ (.B1(net1404),
    .Y(_1713_),
    .A1(_1630_),
    .A2(_1712_));
 sg13g2_nor2_1 _5791_ (.A(net1613),
    .B(_1633_),
    .Y(_1714_));
 sg13g2_a22oi_1 _5792_ (.Y(_0258_),
    .B1(_1713_),
    .B2(_1714_),
    .A2(_3475_),
    .A1(net1613));
 sg13g2_a21oi_1 _5793_ (.A1(net1395),
    .A2(\s0.data_out[14][2] ),
    .Y(_1715_),
    .B1(_1644_));
 sg13g2_a21oi_1 _5794_ (.A1(net1190),
    .A2(_1646_),
    .Y(_1716_),
    .B1(net1613));
 sg13g2_o21ai_1 _5795_ (.B1(_1716_),
    .Y(_1717_),
    .A1(net1190),
    .A2(_1715_));
 sg13g2_o21ai_1 _5796_ (.B1(_1717_),
    .Y(_1718_),
    .A1(net1738),
    .A2(net585));
 sg13g2_inv_1 _5797_ (.Y(_0259_),
    .A(net586));
 sg13g2_nor2_1 _5798_ (.A(net1188),
    .B(_3479_),
    .Y(_1719_));
 sg13g2_o21ai_1 _5799_ (.B1(net1406),
    .Y(_1720_),
    .A1(_1654_),
    .A2(_1719_));
 sg13g2_nor2_1 _5800_ (.A(net1617),
    .B(_1657_),
    .Y(_1721_));
 sg13g2_a22oi_1 _5801_ (.Y(_0260_),
    .B1(_1720_),
    .B2(_1721_),
    .A2(_3473_),
    .A1(net1617));
 sg13g2_a21oi_1 _5802_ (.A1(net1396),
    .A2(net532),
    .Y(_1722_),
    .B1(_1690_));
 sg13g2_a21oi_1 _5803_ (.A1(net1189),
    .A2(_1695_),
    .Y(_1723_),
    .B1(net1617));
 sg13g2_o21ai_1 _5804_ (.B1(_1723_),
    .Y(_1724_),
    .A1(net1189),
    .A2(_1722_));
 sg13g2_o21ai_1 _5805_ (.B1(_1724_),
    .Y(_1725_),
    .A1(net1736),
    .A2(net807));
 sg13g2_inv_1 _5806_ (.Y(_0261_),
    .A(_1725_));
 sg13g2_a21oi_1 _5807_ (.A1(net1399),
    .A2(net783),
    .Y(_1726_),
    .B1(_1684_));
 sg13g2_a21oi_1 _5808_ (.A1(_3380_),
    .A2(_1687_),
    .Y(_1727_),
    .B1(net1617));
 sg13g2_o21ai_1 _5809_ (.B1(_1727_),
    .Y(_1728_),
    .A1(net1189),
    .A2(_1726_));
 sg13g2_o21ai_1 _5810_ (.B1(_1728_),
    .Y(_1729_),
    .A1(net1736),
    .A2(net589));
 sg13g2_inv_1 _5811_ (.Y(_0262_),
    .A(_1729_));
 sg13g2_and2_1 _5812_ (.A(net1398),
    .B(\s0.data_out[14][6] ),
    .X(_1730_));
 sg13g2_o21ai_1 _5813_ (.B1(net1409),
    .Y(_1731_),
    .A1(_1672_),
    .A2(_1730_));
 sg13g2_nand3b_1 _5814_ (.B(_1731_),
    .C(net1736),
    .Y(_1732_),
    .A_N(_1675_));
 sg13g2_o21ai_1 _5815_ (.B1(_1732_),
    .Y(_1733_),
    .A1(net1736),
    .A2(net795));
 sg13g2_inv_1 _5816_ (.Y(_0263_),
    .A(_1733_));
 sg13g2_nor2_1 _5817_ (.A(net1188),
    .B(_3476_),
    .Y(_1734_));
 sg13g2_o21ai_1 _5818_ (.B1(net1409),
    .Y(_1735_),
    .A1(_1665_),
    .A2(_1734_));
 sg13g2_nor2_1 _5819_ (.A(net1618),
    .B(_1668_),
    .Y(_1736_));
 sg13g2_a22oi_1 _5820_ (.Y(_0264_),
    .B1(_1735_),
    .B2(_1736_),
    .A2(_3472_),
    .A1(net1618));
 sg13g2_o21ai_1 _5821_ (.B1(net1397),
    .Y(_1737_),
    .A1(net1633),
    .A2(net1387));
 sg13g2_a21oi_1 _5822_ (.A1(net1623),
    .A2(net1391),
    .Y(_1738_),
    .B1(_1737_));
 sg13g2_inv_1 _5823_ (.Y(_1739_),
    .A(_1738_));
 sg13g2_o21ai_1 _5824_ (.B1(_1739_),
    .Y(_1740_),
    .A1(net1398),
    .A2(_1620_));
 sg13g2_o21ai_1 _5825_ (.B1(_1738_),
    .Y(_1741_),
    .A1(net439),
    .A2(net1391));
 sg13g2_nor2_1 _5826_ (.A(net1387),
    .B(_1737_),
    .Y(_1742_));
 sg13g2_o21ai_1 _5827_ (.B1(net1188),
    .Y(_1743_),
    .A1(net439),
    .A2(net1402));
 sg13g2_nor2b_1 _5828_ (.A(_1742_),
    .B_N(_1743_),
    .Y(_1744_));
 sg13g2_o21ai_1 _5829_ (.B1(net1737),
    .Y(_1745_),
    .A1(net673),
    .A2(_1740_));
 sg13g2_a21oi_1 _5830_ (.A1(_1741_),
    .A2(_1744_),
    .Y(_0265_),
    .B1(_1745_));
 sg13g2_nor2_1 _5831_ (.A(net1618),
    .B(_1740_),
    .Y(_0266_));
 sg13g2_and2_1 _5832_ (.A(net1737),
    .B(net375),
    .X(_0267_));
 sg13g2_nand2_1 _5833_ (.Y(_1746_),
    .A(net1389),
    .B(\s0.data_out[13][2] ));
 sg13g2_mux2_1 _5834_ (.A0(\s0.data_out[14][2] ),
    .A1(\s0.data_out[13][2] ),
    .S(net1389),
    .X(_1747_));
 sg13g2_nor2b_1 _5835_ (.A(net1383),
    .B_N(net1342),
    .Y(_1748_));
 sg13g2_a21o_1 _5836_ (.A2(_1747_),
    .A1(net1383),
    .B1(_1748_),
    .X(_1749_));
 sg13g2_nand2b_1 _5837_ (.Y(_1750_),
    .B(\s0.data_out[13][2] ),
    .A_N(net1400));
 sg13g2_a21oi_1 _5838_ (.A1(_1642_),
    .A2(_1750_),
    .Y(_1751_),
    .B1(net1393));
 sg13g2_a21oi_1 _5839_ (.A1(net1394),
    .A2(_1749_),
    .Y(_1752_),
    .B1(_1751_));
 sg13g2_or2_1 _5840_ (.X(_1753_),
    .B(_1752_),
    .A(net1687));
 sg13g2_nand2_1 _5841_ (.Y(_1754_),
    .A(net1389),
    .B(\s0.data_out[13][1] ));
 sg13g2_o21ai_1 _5842_ (.B1(_1754_),
    .Y(_1755_),
    .A1(net1389),
    .A2(_3481_));
 sg13g2_nor2b_1 _5843_ (.A(net1382),
    .B_N(net1347),
    .Y(_1756_));
 sg13g2_a21o_1 _5844_ (.A2(_1755_),
    .A1(net1382),
    .B1(_1756_),
    .X(_1757_));
 sg13g2_nand2b_1 _5845_ (.Y(_1758_),
    .B(net587),
    .A_N(net1400));
 sg13g2_a21oi_1 _5846_ (.A1(_1628_),
    .A2(_1758_),
    .Y(_1759_),
    .B1(net1393));
 sg13g2_a21oi_1 _5847_ (.A1(net1394),
    .A2(_1757_),
    .Y(_1760_),
    .B1(_1759_));
 sg13g2_mux2_1 _5848_ (.A0(\s0.data_out[14][0] ),
    .A1(\s0.data_out[13][0] ),
    .S(net1390),
    .X(_1761_));
 sg13g2_nor2b_1 _5849_ (.A(net1382),
    .B_N(net1351),
    .Y(_1762_));
 sg13g2_a21oi_1 _5850_ (.A1(net1382),
    .A2(_1761_),
    .Y(_1763_),
    .B1(_1762_));
 sg13g2_nand2b_1 _5851_ (.Y(_1764_),
    .B(net1394),
    .A_N(_1763_));
 sg13g2_mux2_1 _5852_ (.A0(\s0.data_out[13][0] ),
    .A1(\s0.data_out[14][0] ),
    .S(net1400),
    .X(_1765_));
 sg13g2_nand2_1 _5853_ (.Y(_1766_),
    .A(net1188),
    .B(_1765_));
 sg13g2_a221oi_1 _5854_ (.B2(_1766_),
    .C1(net1702),
    .B1(_1764_),
    .A1(net1697),
    .Y(_1767_),
    .A2(_1760_));
 sg13g2_o21ai_1 _5855_ (.B1(_1753_),
    .Y(_1768_),
    .A1(net1697),
    .A2(_1760_));
 sg13g2_nand2_1 _5856_ (.Y(_1769_),
    .A(net1390),
    .B(net692));
 sg13g2_o21ai_1 _5857_ (.B1(_1769_),
    .Y(_1770_),
    .A1(net1391),
    .A2(_3479_));
 sg13g2_nor2_1 _5858_ (.A(net1383),
    .B(net1162),
    .Y(_1771_));
 sg13g2_a21o_1 _5859_ (.A2(_1770_),
    .A1(net1383),
    .B1(_1771_),
    .X(_1772_));
 sg13g2_nand2b_1 _5860_ (.Y(_1773_),
    .B(net692),
    .A_N(net1400));
 sg13g2_a21oi_1 _5861_ (.A1(_1652_),
    .A2(_1773_),
    .Y(_1774_),
    .B1(net1395));
 sg13g2_a21oi_1 _5862_ (.A1(net1395),
    .A2(_1772_),
    .Y(_1775_),
    .B1(_1774_));
 sg13g2_a22oi_1 _5863_ (.Y(_1776_),
    .B1(_1775_),
    .B2(net1681),
    .A2(_1752_),
    .A1(net1687));
 sg13g2_o21ai_1 _5864_ (.B1(_1776_),
    .Y(_1777_),
    .A1(_1767_),
    .A2(_1768_));
 sg13g2_nand2_1 _5865_ (.Y(_1778_),
    .A(net1392),
    .B(net608));
 sg13g2_mux2_1 _5866_ (.A0(\s0.data_out[14][7] ),
    .A1(\s0.data_out[13][7] ),
    .S(net1391),
    .X(_1779_));
 sg13g2_nor2b_1 _5867_ (.A(net1387),
    .B_N(net1323),
    .Y(_1780_));
 sg13g2_a21o_1 _5868_ (.A2(_1779_),
    .A1(net1387),
    .B1(_1780_),
    .X(_1781_));
 sg13g2_nand2b_1 _5869_ (.Y(_1782_),
    .B(net608),
    .A_N(net1402));
 sg13g2_a21oi_1 _5870_ (.A1(_1663_),
    .A2(_1782_),
    .Y(_1783_),
    .B1(net1397));
 sg13g2_a21oi_1 _5871_ (.A1(net1398),
    .A2(_1781_),
    .Y(_1784_),
    .B1(_1783_));
 sg13g2_nand2_1 _5872_ (.Y(_1785_),
    .A(net1391),
    .B(net760));
 sg13g2_mux2_1 _5873_ (.A0(\s0.data_out[14][6] ),
    .A1(\s0.data_out[13][6] ),
    .S(net1392),
    .X(_1786_));
 sg13g2_nor2b_1 _5874_ (.A(net1387),
    .B_N(net1328),
    .Y(_1787_));
 sg13g2_a21o_1 _5875_ (.A2(_1786_),
    .A1(net1387),
    .B1(_1787_),
    .X(_1788_));
 sg13g2_nand2b_1 _5876_ (.Y(_1789_),
    .B(\s0.data_out[13][6] ),
    .A_N(net1402));
 sg13g2_a21oi_1 _5877_ (.A1(_1670_),
    .A2(_1789_),
    .Y(_1790_),
    .B1(net1397));
 sg13g2_a21oi_1 _5878_ (.A1(net1398),
    .A2(_1788_),
    .Y(_1791_),
    .B1(_1790_));
 sg13g2_a22oi_1 _5879_ (.Y(_1792_),
    .B1(_1791_),
    .B2(net1654),
    .A2(_1784_),
    .A1(net1642));
 sg13g2_or2_1 _5880_ (.X(_1793_),
    .B(_1784_),
    .A(net1642));
 sg13g2_or2_1 _5881_ (.X(_1794_),
    .B(_1791_),
    .A(net1654));
 sg13g2_and3_1 _5882_ (.X(_1795_),
    .A(_1792_),
    .B(_1793_),
    .C(_1794_));
 sg13g2_nand3_1 _5883_ (.B(_1793_),
    .C(_1794_),
    .A(_1792_),
    .Y(_1796_));
 sg13g2_nand2_1 _5884_ (.Y(_1797_),
    .A(net1391),
    .B(net518));
 sg13g2_o21ai_1 _5885_ (.B1(_1797_),
    .Y(_1798_),
    .A1(net1391),
    .A2(_3478_));
 sg13g2_nor2b_1 _5886_ (.A(net1388),
    .B_N(net1337),
    .Y(_1799_));
 sg13g2_a21oi_1 _5887_ (.A1(net1388),
    .A2(_1798_),
    .Y(_1800_),
    .B1(_1799_));
 sg13g2_o21ai_1 _5888_ (.B1(_1691_),
    .Y(_1801_),
    .A1(net1401),
    .A2(_3484_));
 sg13g2_nand2_1 _5889_ (.Y(_1802_),
    .A(_3381_),
    .B(_1801_));
 sg13g2_o21ai_1 _5890_ (.B1(_1802_),
    .Y(_1803_),
    .A1(_3381_),
    .A2(_1800_));
 sg13g2_nand2_1 _5891_ (.Y(_1804_),
    .A(net1392),
    .B(net583));
 sg13g2_mux2_1 _5892_ (.A0(\s0.data_out[14][5] ),
    .A1(\s0.data_out[13][5] ),
    .S(net1391),
    .X(_1805_));
 sg13g2_nor2b_1 _5893_ (.A(net1387),
    .B_N(net1333),
    .Y(_1806_));
 sg13g2_a21o_1 _5894_ (.A2(_1805_),
    .A1(net1387),
    .B1(_1806_),
    .X(_1807_));
 sg13g2_nand2b_1 _5895_ (.Y(_1808_),
    .B(net583),
    .A_N(net1402));
 sg13g2_a21oi_1 _5896_ (.A1(_1682_),
    .A2(_1808_),
    .Y(_1809_),
    .B1(net1397));
 sg13g2_a21oi_1 _5897_ (.A1(net1397),
    .A2(_1807_),
    .Y(_1810_),
    .B1(_1809_));
 sg13g2_nand2_1 _5898_ (.Y(_1811_),
    .A(net1662),
    .B(_1810_));
 sg13g2_nor2_1 _5899_ (.A(net1663),
    .B(_1810_),
    .Y(_1812_));
 sg13g2_xnor2_1 _5900_ (.Y(_1813_),
    .A(_3406_),
    .B(_1803_));
 sg13g2_o21ai_1 _5901_ (.B1(_1811_),
    .Y(_1814_),
    .A1(net1681),
    .A2(_1775_));
 sg13g2_nor4_1 _5902_ (.A(_1796_),
    .B(_1812_),
    .C(_1813_),
    .D(_1814_),
    .Y(_1815_));
 sg13g2_or3_1 _5903_ (.A(_3406_),
    .B(_1803_),
    .C(_1812_),
    .X(_1816_));
 sg13g2_nand2_1 _5904_ (.Y(_1817_),
    .A(_1811_),
    .B(_1816_));
 sg13g2_nand2b_1 _5905_ (.Y(_1818_),
    .B(_1793_),
    .A_N(_1792_));
 sg13g2_a221oi_1 _5906_ (.B2(_1795_),
    .C1(_1740_),
    .B1(_1817_),
    .A1(_1777_),
    .Y(_1819_),
    .A2(_1815_));
 sg13g2_or2_1 _5907_ (.X(_1820_),
    .B(net1557),
    .A(net392));
 sg13g2_a21oi_1 _5908_ (.A1(_1818_),
    .A2(_1819_),
    .Y(_0268_),
    .B1(_1820_));
 sg13g2_a21oi_1 _5909_ (.A1(net1382),
    .A2(\s0.data_out[13][0] ),
    .Y(_1821_),
    .B1(_1762_));
 sg13g2_a21oi_1 _5910_ (.A1(net1188),
    .A2(_1765_),
    .Y(_1822_),
    .B1(net1613));
 sg13g2_o21ai_1 _5911_ (.B1(_1822_),
    .Y(_1823_),
    .A1(net1188),
    .A2(_1821_));
 sg13g2_o21ai_1 _5912_ (.B1(_1823_),
    .Y(_1824_),
    .A1(net1738),
    .A2(net636));
 sg13g2_inv_1 _5913_ (.Y(_0269_),
    .A(net637));
 sg13g2_and2_1 _5914_ (.A(net1382),
    .B(net587),
    .X(_1825_));
 sg13g2_o21ai_1 _5915_ (.B1(net1393),
    .Y(_1826_),
    .A1(_1756_),
    .A2(_1825_));
 sg13g2_nor2_1 _5916_ (.A(net1613),
    .B(_1759_),
    .Y(_1827_));
 sg13g2_a22oi_1 _5917_ (.Y(_0270_),
    .B1(_1826_),
    .B2(_1827_),
    .A2(_3481_),
    .A1(net1614));
 sg13g2_nor2_1 _5918_ (.A(net1186),
    .B(_3486_),
    .Y(_1828_));
 sg13g2_o21ai_1 _5919_ (.B1(net1394),
    .Y(_1829_),
    .A1(_1748_),
    .A2(_1828_));
 sg13g2_nor2_1 _5920_ (.A(net1614),
    .B(_1751_),
    .Y(_1830_));
 sg13g2_a22oi_1 _5921_ (.Y(_0271_),
    .B1(_1829_),
    .B2(_1830_),
    .A2(_3480_),
    .A1(net1613));
 sg13g2_nor2_1 _5922_ (.A(net1187),
    .B(_3485_),
    .Y(_1831_));
 sg13g2_o21ai_1 _5923_ (.B1(net1394),
    .Y(_1832_),
    .A1(_1771_),
    .A2(_1831_));
 sg13g2_nor2_1 _5924_ (.A(net1613),
    .B(_1774_),
    .Y(_1833_));
 sg13g2_a22oi_1 _5925_ (.Y(_0272_),
    .B1(_1832_),
    .B2(_1833_),
    .A2(_3479_),
    .A1(net1613));
 sg13g2_a21oi_1 _5926_ (.A1(net1388),
    .A2(net518),
    .Y(_1834_),
    .B1(_1799_));
 sg13g2_a21oi_1 _5927_ (.A1(_3381_),
    .A2(_1801_),
    .Y(_1835_),
    .B1(net1619));
 sg13g2_o21ai_1 _5928_ (.B1(_1835_),
    .Y(_1836_),
    .A1(net1188),
    .A2(_1834_));
 sg13g2_o21ai_1 _5929_ (.B1(_1836_),
    .Y(_1837_),
    .A1(net1736),
    .A2(net532));
 sg13g2_inv_1 _5930_ (.Y(_0273_),
    .A(net533));
 sg13g2_nor2_1 _5931_ (.A(net1187),
    .B(_3483_),
    .Y(_1838_));
 sg13g2_o21ai_1 _5932_ (.B1(net1397),
    .Y(_1839_),
    .A1(_1806_),
    .A2(_1838_));
 sg13g2_nor2_1 _5933_ (.A(net1618),
    .B(_1809_),
    .Y(_1840_));
 sg13g2_a22oi_1 _5934_ (.Y(_0274_),
    .B1(_1839_),
    .B2(_1840_),
    .A2(_3477_),
    .A1(net1618));
 sg13g2_and2_1 _5935_ (.A(net1388),
    .B(\s0.data_out[13][6] ),
    .X(_1841_));
 sg13g2_o21ai_1 _5936_ (.B1(net1397),
    .Y(_1842_),
    .A1(_1787_),
    .A2(_1841_));
 sg13g2_nand3b_1 _5937_ (.B(_1842_),
    .C(net1737),
    .Y(_1843_),
    .A_N(_1790_));
 sg13g2_o21ai_1 _5938_ (.B1(_1843_),
    .Y(_1844_),
    .A1(net1737),
    .A2(net721));
 sg13g2_inv_1 _5939_ (.Y(_0275_),
    .A(net722));
 sg13g2_nor2_1 _5940_ (.A(net1187),
    .B(_3482_),
    .Y(_1845_));
 sg13g2_o21ai_1 _5941_ (.B1(net1397),
    .Y(_1846_),
    .A1(_1780_),
    .A2(_1845_));
 sg13g2_nor2_1 _5942_ (.A(net1619),
    .B(_1783_),
    .Y(_1847_));
 sg13g2_a22oi_1 _5943_ (.Y(_0276_),
    .B1(_1846_),
    .B2(_1847_),
    .A2(_3476_),
    .A1(net1618));
 sg13g2_o21ai_1 _5944_ (.B1(net1386),
    .Y(_1848_),
    .A1(net1632),
    .A2(net1375));
 sg13g2_nor2b_1 _5945_ (.A(net1632),
    .B_N(net1381),
    .Y(_1849_));
 sg13g2_nor2_1 _5946_ (.A(_1848_),
    .B(_1849_),
    .Y(_1850_));
 sg13g2_a21oi_1 _5947_ (.A1(net1623),
    .A2(net1390),
    .Y(_1851_),
    .B1(net1385));
 sg13g2_nor2_1 _5948_ (.A(_1850_),
    .B(_1851_),
    .Y(_1852_));
 sg13g2_o21ai_1 _5949_ (.B1(_1850_),
    .Y(_1853_),
    .A1(\s0.was_valid_out[12] [0]),
    .A2(net1381));
 sg13g2_nor2_1 _5950_ (.A(net1375),
    .B(_1848_),
    .Y(_1854_));
 sg13g2_o21ai_1 _5951_ (.B1(net1187),
    .Y(_1855_),
    .A1(\s0.was_valid_out[12] [0]),
    .A2(net1390));
 sg13g2_nand2_1 _5952_ (.Y(_1856_),
    .A(_1853_),
    .B(_1855_));
 sg13g2_o21ai_1 _5953_ (.B1(net1738),
    .Y(_1857_),
    .A1(_1854_),
    .A2(_1856_));
 sg13g2_a21oi_1 _5954_ (.A1(_3364_),
    .A2(_1852_),
    .Y(_0277_),
    .B1(_1857_));
 sg13g2_nor3_1 _5955_ (.A(net1616),
    .B(_1850_),
    .C(_1851_),
    .Y(_0278_));
 sg13g2_and2_1 _5956_ (.A(net1738),
    .B(net386),
    .X(_0279_));
 sg13g2_nand2_1 _5957_ (.Y(_1858_),
    .A(net1378),
    .B(net749));
 sg13g2_o21ai_1 _5958_ (.B1(_1858_),
    .Y(_1859_),
    .A1(net1378),
    .A2(_3486_));
 sg13g2_nor2b_1 _5959_ (.A(net1369),
    .B_N(net1343),
    .Y(_1860_));
 sg13g2_a21oi_1 _5960_ (.A1(net1369),
    .A2(_1859_),
    .Y(_1861_),
    .B1(_1860_));
 sg13g2_o21ai_1 _5961_ (.B1(_1746_),
    .Y(_1862_),
    .A1(net1389),
    .A2(_3490_));
 sg13g2_nand2_1 _5962_ (.Y(_1863_),
    .A(net1185),
    .B(_1862_));
 sg13g2_o21ai_1 _5963_ (.B1(_1863_),
    .Y(_1864_),
    .A1(net1185),
    .A2(_1861_));
 sg13g2_nand2_1 _5964_ (.Y(_1865_),
    .A(net1378),
    .B(net820));
 sg13g2_mux2_1 _5965_ (.A0(\s0.data_out[13][1] ),
    .A1(\s0.data_out[12][1] ),
    .S(net1378),
    .X(_1866_));
 sg13g2_nor2b_1 _5966_ (.A(net1369),
    .B_N(net1347),
    .Y(_1867_));
 sg13g2_a21oi_1 _5967_ (.A1(net1369),
    .A2(_1866_),
    .Y(_1868_),
    .B1(_1867_));
 sg13g2_nand2b_1 _5968_ (.Y(_1869_),
    .B(net1382),
    .A_N(_1868_));
 sg13g2_o21ai_1 _5969_ (.B1(_1754_),
    .Y(_1870_),
    .A1(net1389),
    .A2(_3491_));
 sg13g2_nand2_1 _5970_ (.Y(_1871_),
    .A(net1186),
    .B(_1870_));
 sg13g2_nand3_1 _5971_ (.B(_1869_),
    .C(_1871_),
    .A(net1698),
    .Y(_1872_));
 sg13g2_mux2_1 _5972_ (.A0(\s0.data_out[13][0] ),
    .A1(\s0.data_out[12][0] ),
    .S(net1378),
    .X(_1873_));
 sg13g2_nor2b_1 _5973_ (.A(net1369),
    .B_N(net1351),
    .Y(_1874_));
 sg13g2_a21oi_1 _5974_ (.A1(net1369),
    .A2(_1873_),
    .Y(_1875_),
    .B1(_1874_));
 sg13g2_mux2_1 _5975_ (.A0(\s0.data_out[12][0] ),
    .A1(\s0.data_out[13][0] ),
    .S(net1389),
    .X(_1876_));
 sg13g2_nand2_1 _5976_ (.Y(_1877_),
    .A(net1185),
    .B(_1876_));
 sg13g2_o21ai_1 _5977_ (.B1(_1877_),
    .Y(_1878_),
    .A1(net1185),
    .A2(_1875_));
 sg13g2_and2_1 _5978_ (.A(_3418_),
    .B(_1878_),
    .X(_1879_));
 sg13g2_a21oi_1 _5979_ (.A1(_1869_),
    .A2(_1871_),
    .Y(_1880_),
    .B1(net1698));
 sg13g2_a221oi_1 _5980_ (.B2(_1879_),
    .C1(_1880_),
    .B1(_1872_),
    .A1(net1563),
    .Y(_1881_),
    .A2(_1864_));
 sg13g2_nand2_1 _5981_ (.Y(_1882_),
    .A(net1379),
    .B(net580));
 sg13g2_o21ai_1 _5982_ (.B1(_1882_),
    .Y(_1883_),
    .A1(net1379),
    .A2(_3485_));
 sg13g2_nor2_1 _5983_ (.A(net1372),
    .B(net1162),
    .Y(_1884_));
 sg13g2_a21o_1 _5984_ (.A2(_1883_),
    .A1(net1372),
    .B1(_1884_),
    .X(_1885_));
 sg13g2_nand2b_1 _5985_ (.Y(_1886_),
    .B(net580),
    .A_N(net1389));
 sg13g2_a21oi_1 _5986_ (.A1(_1769_),
    .A2(_1886_),
    .Y(_1887_),
    .B1(net1382));
 sg13g2_a21oi_1 _5987_ (.A1(net1383),
    .A2(_1885_),
    .Y(_1888_),
    .B1(_1887_));
 sg13g2_nand2_1 _5988_ (.Y(_1889_),
    .A(net1681),
    .B(_1888_));
 sg13g2_or2_1 _5989_ (.X(_1890_),
    .B(_1864_),
    .A(net1563));
 sg13g2_nand3b_1 _5990_ (.B(_1889_),
    .C(_1890_),
    .Y(_1891_),
    .A_N(_1881_));
 sg13g2_nand2_1 _5991_ (.Y(_1892_),
    .A(net1381),
    .B(\s0.data_out[12][4] ));
 sg13g2_o21ai_1 _5992_ (.B1(_1892_),
    .Y(_1893_),
    .A1(net1381),
    .A2(_3484_));
 sg13g2_nor2b_1 _5993_ (.A(net1376),
    .B_N(net1338),
    .Y(_1894_));
 sg13g2_a21o_1 _5994_ (.A2(_1893_),
    .A1(net1376),
    .B1(_1894_),
    .X(_1895_));
 sg13g2_nand2b_1 _5995_ (.Y(_1896_),
    .B(net453),
    .A_N(net1390));
 sg13g2_a21oi_1 _5996_ (.A1(_1797_),
    .A2(_1896_),
    .Y(_1897_),
    .B1(net1383));
 sg13g2_a21oi_1 _5997_ (.A1(net1384),
    .A2(_1895_),
    .Y(_1898_),
    .B1(_1897_));
 sg13g2_nand2_1 _5998_ (.Y(_1899_),
    .A(net1672),
    .B(_1898_));
 sg13g2_nand2_1 _5999_ (.Y(_1900_),
    .A(net1380),
    .B(net660));
 sg13g2_mux2_1 _6000_ (.A0(\s0.data_out[13][5] ),
    .A1(\s0.data_out[12][5] ),
    .S(net1381),
    .X(_1901_));
 sg13g2_nor2b_1 _6001_ (.A(net1376),
    .B_N(net1333),
    .Y(_1902_));
 sg13g2_a21o_1 _6002_ (.A2(_1901_),
    .A1(net1376),
    .B1(_1902_),
    .X(_1903_));
 sg13g2_nand2b_1 _6003_ (.Y(_1904_),
    .B(\s0.data_out[12][5] ),
    .A_N(net1392));
 sg13g2_a21oi_1 _6004_ (.A1(_1804_),
    .A2(_1904_),
    .Y(_1905_),
    .B1(net1384));
 sg13g2_a21oi_1 _6005_ (.A1(net1384),
    .A2(_1903_),
    .Y(_1906_),
    .B1(_1905_));
 sg13g2_nor2_1 _6006_ (.A(net1662),
    .B(_1906_),
    .Y(_1907_));
 sg13g2_nand2_1 _6007_ (.Y(_1908_),
    .A(net1662),
    .B(_1906_));
 sg13g2_o21ai_1 _6008_ (.B1(_1908_),
    .Y(_1909_),
    .A1(net1682),
    .A2(_1888_));
 sg13g2_xnor2_1 _6009_ (.Y(_1910_),
    .A(net1672),
    .B(_1898_));
 sg13g2_nand2_1 _6010_ (.Y(_1911_),
    .A(net1380),
    .B(\s0.data_out[12][6] ));
 sg13g2_mux2_1 _6011_ (.A0(\s0.data_out[13][6] ),
    .A1(\s0.data_out[12][6] ),
    .S(net1381),
    .X(_1912_));
 sg13g2_nor2b_1 _6012_ (.A(net1375),
    .B_N(net1328),
    .Y(_1913_));
 sg13g2_a21o_1 _6013_ (.A2(_1912_),
    .A1(net1375),
    .B1(_1913_),
    .X(_1914_));
 sg13g2_nand2b_1 _6014_ (.Y(_1915_),
    .B(\s0.data_out[12][6] ),
    .A_N(net1390));
 sg13g2_a21oi_1 _6015_ (.A1(_1785_),
    .A2(_1915_),
    .Y(_1916_),
    .B1(net1384));
 sg13g2_a21oi_1 _6016_ (.A1(net1384),
    .A2(_1914_),
    .Y(_1917_),
    .B1(_1916_));
 sg13g2_nand2_1 _6017_ (.Y(_1918_),
    .A(net1380),
    .B(net522));
 sg13g2_mux2_1 _6018_ (.A0(\s0.data_out[13][7] ),
    .A1(\s0.data_out[12][7] ),
    .S(net1381),
    .X(_1919_));
 sg13g2_nor2b_1 _6019_ (.A(net1375),
    .B_N(net1323),
    .Y(_1920_));
 sg13g2_a21o_1 _6020_ (.A2(_1919_),
    .A1(net1376),
    .B1(_1920_),
    .X(_1921_));
 sg13g2_nand2b_1 _6021_ (.Y(_1922_),
    .B(net522),
    .A_N(net1390));
 sg13g2_a21oi_1 _6022_ (.A1(_1778_),
    .A2(_1922_),
    .Y(_1923_),
    .B1(net1385));
 sg13g2_a21oi_1 _6023_ (.A1(net1385),
    .A2(_1921_),
    .Y(_1924_),
    .B1(_1923_));
 sg13g2_a22oi_1 _6024_ (.Y(_1925_),
    .B1(_1924_),
    .B2(net1642),
    .A2(_1917_),
    .A1(net1652));
 sg13g2_or2_1 _6025_ (.X(_1926_),
    .B(_1917_),
    .A(net1652));
 sg13g2_nor2_1 _6026_ (.A(net1642),
    .B(_1924_),
    .Y(_1927_));
 sg13g2_or2_1 _6027_ (.X(_1928_),
    .B(_1924_),
    .A(net1642));
 sg13g2_and3_1 _6028_ (.X(_1929_),
    .A(_1925_),
    .B(_1926_),
    .C(_1928_));
 sg13g2_nand3_1 _6029_ (.B(_1926_),
    .C(_1928_),
    .A(_1925_),
    .Y(_1930_));
 sg13g2_nor4_1 _6030_ (.A(_1907_),
    .B(_1909_),
    .C(_1910_),
    .D(_1930_),
    .Y(_1931_));
 sg13g2_o21ai_1 _6031_ (.B1(_1908_),
    .Y(_1932_),
    .A1(_1899_),
    .A2(_1907_));
 sg13g2_o21ai_1 _6032_ (.B1(_1852_),
    .Y(_1933_),
    .A1(_1925_),
    .A2(_1927_));
 sg13g2_a221oi_1 _6033_ (.B2(_1929_),
    .C1(_1933_),
    .B1(_1932_),
    .A1(_1891_),
    .Y(_1934_),
    .A2(_1931_));
 sg13g2_nor3_1 _6034_ (.A(net375),
    .B(net1557),
    .C(_1934_),
    .Y(_0280_));
 sg13g2_a21oi_1 _6035_ (.A1(net1369),
    .A2(\s0.data_out[12][0] ),
    .Y(_1935_),
    .B1(_1874_));
 sg13g2_a21oi_1 _6036_ (.A1(net1185),
    .A2(_1876_),
    .Y(_1936_),
    .B1(net1614));
 sg13g2_o21ai_1 _6037_ (.B1(_1936_),
    .Y(_1937_),
    .A1(net1185),
    .A2(_1935_));
 sg13g2_o21ai_1 _6038_ (.B1(_1937_),
    .Y(_1938_),
    .A1(net1729),
    .A2(net685));
 sg13g2_inv_1 _6039_ (.Y(_0281_),
    .A(net686));
 sg13g2_a21oi_1 _6040_ (.A1(net1369),
    .A2(\s0.data_out[12][1] ),
    .Y(_1939_),
    .B1(_1867_));
 sg13g2_a21oi_1 _6041_ (.A1(net1185),
    .A2(_1870_),
    .Y(_1940_),
    .B1(net1614));
 sg13g2_o21ai_1 _6042_ (.B1(_1940_),
    .Y(_1941_),
    .A1(net1185),
    .A2(_1939_));
 sg13g2_o21ai_1 _6043_ (.B1(_1941_),
    .Y(_1942_),
    .A1(net1729),
    .A2(net587));
 sg13g2_inv_1 _6044_ (.Y(_0282_),
    .A(net588));
 sg13g2_a21oi_1 _6045_ (.A1(net1370),
    .A2(\s0.data_out[12][2] ),
    .Y(_1943_),
    .B1(_1860_));
 sg13g2_a21oi_1 _6046_ (.A1(net1186),
    .A2(_1862_),
    .Y(_1944_),
    .B1(net1614));
 sg13g2_o21ai_1 _6047_ (.B1(_1944_),
    .Y(_1945_),
    .A1(net1186),
    .A2(_1943_));
 sg13g2_o21ai_1 _6048_ (.B1(_1945_),
    .Y(_1946_),
    .A1(net1729),
    .A2(net687));
 sg13g2_inv_1 _6049_ (.Y(_0283_),
    .A(net688));
 sg13g2_and2_1 _6050_ (.A(net1372),
    .B(net580),
    .X(_1947_));
 sg13g2_o21ai_1 _6051_ (.B1(net1383),
    .Y(_1948_),
    .A1(_1884_),
    .A2(_1947_));
 sg13g2_nor2_1 _6052_ (.A(net1615),
    .B(_1887_),
    .Y(_1949_));
 sg13g2_a22oi_1 _6053_ (.Y(_0284_),
    .B1(_1948_),
    .B2(_1949_),
    .A2(_3485_),
    .A1(net1615));
 sg13g2_and2_1 _6054_ (.A(net1376),
    .B(net453),
    .X(_1950_));
 sg13g2_o21ai_1 _6055_ (.B1(net1384),
    .Y(_1951_),
    .A1(_1894_),
    .A2(_1950_));
 sg13g2_nor2_1 _6056_ (.A(net1615),
    .B(_1897_),
    .Y(_1952_));
 sg13g2_a22oi_1 _6057_ (.Y(_0285_),
    .B1(_1951_),
    .B2(_1952_),
    .A2(_3484_),
    .A1(net1615));
 sg13g2_and2_1 _6058_ (.A(net1376),
    .B(\s0.data_out[12][5] ),
    .X(_1953_));
 sg13g2_o21ai_1 _6059_ (.B1(net1384),
    .Y(_1954_),
    .A1(_1902_),
    .A2(_1953_));
 sg13g2_nor2_1 _6060_ (.A(net1615),
    .B(_1905_),
    .Y(_1955_));
 sg13g2_a22oi_1 _6061_ (.Y(_0286_),
    .B1(_1954_),
    .B2(_1955_),
    .A2(_3483_),
    .A1(net1615));
 sg13g2_and2_1 _6062_ (.A(net1375),
    .B(\s0.data_out[12][6] ),
    .X(_1956_));
 sg13g2_o21ai_1 _6063_ (.B1(net1385),
    .Y(_1957_),
    .A1(_1913_),
    .A2(_1956_));
 sg13g2_nand3b_1 _6064_ (.B(_1957_),
    .C(net1738),
    .Y(_1958_),
    .A_N(_1916_));
 sg13g2_o21ai_1 _6065_ (.B1(_1958_),
    .Y(_1959_),
    .A1(net1738),
    .A2(net760));
 sg13g2_inv_1 _6066_ (.Y(_0287_),
    .A(net761));
 sg13g2_and2_1 _6067_ (.A(net1375),
    .B(net522),
    .X(_1960_));
 sg13g2_o21ai_1 _6068_ (.B1(net1385),
    .Y(_1961_),
    .A1(_1920_),
    .A2(_1960_));
 sg13g2_nor2_1 _6069_ (.A(net1615),
    .B(_1923_),
    .Y(_1962_));
 sg13g2_a22oi_1 _6070_ (.Y(_0288_),
    .B1(_1961_),
    .B2(_1962_),
    .A2(_3482_),
    .A1(net1615));
 sg13g2_o21ai_1 _6071_ (.B1(net1373),
    .Y(_1963_),
    .A1(net1630),
    .A2(net1362));
 sg13g2_nor2b_1 _6072_ (.A(net1631),
    .B_N(net1367),
    .Y(_1964_));
 sg13g2_nor2_1 _6073_ (.A(_1963_),
    .B(_1964_),
    .Y(_1965_));
 sg13g2_inv_1 _6074_ (.Y(_1966_),
    .A(_1965_));
 sg13g2_o21ai_1 _6075_ (.B1(_1966_),
    .Y(_1967_),
    .A1(net1375),
    .A2(_1849_));
 sg13g2_nor2_1 _6076_ (.A(net462),
    .B(_1967_),
    .Y(_1968_));
 sg13g2_o21ai_1 _6077_ (.B1(_1965_),
    .Y(_1969_),
    .A1(net445),
    .A2(net1366));
 sg13g2_nor2_1 _6078_ (.A(net1362),
    .B(_1963_),
    .Y(_1970_));
 sg13g2_nor2_1 _6079_ (.A(net445),
    .B(net1380),
    .Y(_1971_));
 sg13g2_o21ai_1 _6080_ (.B1(_1969_),
    .Y(_1972_),
    .A1(net1373),
    .A2(_1971_));
 sg13g2_o21ai_1 _6081_ (.B1(net1728),
    .Y(_1973_),
    .A1(_1970_),
    .A2(_1972_));
 sg13g2_nor2_1 _6082_ (.A(_1968_),
    .B(_1973_),
    .Y(_0289_));
 sg13g2_nor2_1 _6083_ (.A(net1616),
    .B(_1967_),
    .Y(_0290_));
 sg13g2_and2_1 _6084_ (.A(net1728),
    .B(net385),
    .X(_0291_));
 sg13g2_nand2_1 _6085_ (.Y(_1974_),
    .A(net1364),
    .B(net571));
 sg13g2_mux2_1 _6086_ (.A0(\s0.data_out[12][2] ),
    .A1(\s0.data_out[11][2] ),
    .S(net1365),
    .X(_1975_));
 sg13g2_nor2b_1 _6087_ (.A(net1359),
    .B_N(net1342),
    .Y(_1976_));
 sg13g2_a21o_1 _6088_ (.A2(_1975_),
    .A1(net1359),
    .B1(_1976_),
    .X(_1977_));
 sg13g2_nand2b_1 _6089_ (.Y(_1978_),
    .B(net571),
    .A_N(net1378));
 sg13g2_a21oi_1 _6090_ (.A1(_1858_),
    .A2(_1978_),
    .Y(_1979_),
    .B1(net1370));
 sg13g2_a21oi_1 _6091_ (.A1(net1368),
    .A2(_1977_),
    .Y(_1980_),
    .B1(_1979_));
 sg13g2_or2_1 _6092_ (.X(_1981_),
    .B(_1980_),
    .A(net1687));
 sg13g2_nor2b_1 _6093_ (.A(net1359),
    .B_N(net1346),
    .Y(_1982_));
 sg13g2_nand2_1 _6094_ (.Y(_1983_),
    .A(net1364),
    .B(net753));
 sg13g2_o21ai_1 _6095_ (.B1(_1983_),
    .Y(_1984_),
    .A1(net1365),
    .A2(_3491_));
 sg13g2_a21o_1 _6096_ (.A2(_1984_),
    .A1(net1359),
    .B1(_1982_),
    .X(_1985_));
 sg13g2_nand2b_1 _6097_ (.Y(_1986_),
    .B(net753),
    .A_N(net1378));
 sg13g2_a21oi_1 _6098_ (.A1(_1865_),
    .A2(_1986_),
    .Y(_1987_),
    .B1(net1368));
 sg13g2_a21oi_1 _6099_ (.A1(net1368),
    .A2(_1985_),
    .Y(_1988_),
    .B1(_1987_));
 sg13g2_mux2_1 _6100_ (.A0(\s0.data_out[12][0] ),
    .A1(\s0.data_out[11][0] ),
    .S(net1365),
    .X(_1989_));
 sg13g2_nor2b_1 _6101_ (.A(\s0.shift_out[11] [0]),
    .B_N(\s0.data_new_delayed[0] ),
    .Y(_1990_));
 sg13g2_a21oi_1 _6102_ (.A1(net1359),
    .A2(_1989_),
    .Y(_1991_),
    .B1(_1990_));
 sg13g2_nand2b_1 _6103_ (.Y(_1992_),
    .B(net1368),
    .A_N(_1991_));
 sg13g2_mux2_1 _6104_ (.A0(\s0.data_out[11][0] ),
    .A1(\s0.data_out[12][0] ),
    .S(net1378),
    .X(_1993_));
 sg13g2_nand2b_1 _6105_ (.Y(_1994_),
    .B(_1993_),
    .A_N(net1368));
 sg13g2_o21ai_1 _6106_ (.B1(_1981_),
    .Y(_1995_),
    .A1(net1697),
    .A2(_1988_));
 sg13g2_a221oi_1 _6107_ (.B2(_1994_),
    .C1(net1702),
    .B1(_1992_),
    .A1(net1697),
    .Y(_1996_),
    .A2(_1988_));
 sg13g2_nand2_1 _6108_ (.Y(_1997_),
    .A(net1364),
    .B(\s0.data_out[11][3] ));
 sg13g2_o21ai_1 _6109_ (.B1(_1997_),
    .Y(_1998_),
    .A1(net1365),
    .A2(_3489_));
 sg13g2_nor2_1 _6110_ (.A(net1359),
    .B(net1162),
    .Y(_1999_));
 sg13g2_a21o_1 _6111_ (.A2(_1998_),
    .A1(net1359),
    .B1(_1999_),
    .X(_2000_));
 sg13g2_nand2b_1 _6112_ (.Y(_2001_),
    .B(\s0.data_out[11][3] ),
    .A_N(net1379));
 sg13g2_a21oi_1 _6113_ (.A1(_1882_),
    .A2(_2001_),
    .Y(_2002_),
    .B1(net1371));
 sg13g2_a21oi_1 _6114_ (.A1(net1371),
    .A2(_2000_),
    .Y(_2003_),
    .B1(_2002_));
 sg13g2_a22oi_1 _6115_ (.Y(_2004_),
    .B1(_2003_),
    .B2(net1681),
    .A2(_1980_),
    .A1(net1687));
 sg13g2_o21ai_1 _6116_ (.B1(_2004_),
    .Y(_2005_),
    .A1(_1995_),
    .A2(_1996_));
 sg13g2_nand2_1 _6117_ (.Y(_2006_),
    .A(net1366),
    .B(net718));
 sg13g2_mux2_1 _6118_ (.A0(\s0.data_out[12][6] ),
    .A1(\s0.data_out[11][6] ),
    .S(net1367),
    .X(_2007_));
 sg13g2_nor2b_1 _6119_ (.A(net1363),
    .B_N(net1327),
    .Y(_2008_));
 sg13g2_a21o_1 _6120_ (.A2(_2007_),
    .A1(net1362),
    .B1(_2008_),
    .X(_2009_));
 sg13g2_nand2b_1 _6121_ (.Y(_2010_),
    .B(\s0.data_out[11][6] ),
    .A_N(net1380));
 sg13g2_a21oi_1 _6122_ (.A1(_1911_),
    .A2(_2010_),
    .Y(_2011_),
    .B1(net1374));
 sg13g2_a21oi_1 _6123_ (.A1(net1374),
    .A2(_2009_),
    .Y(_2012_),
    .B1(_2011_));
 sg13g2_nand2_1 _6124_ (.Y(_2013_),
    .A(net1366),
    .B(net568));
 sg13g2_mux2_1 _6125_ (.A0(\s0.data_out[12][7] ),
    .A1(\s0.data_out[11][7] ),
    .S(net1367),
    .X(_2014_));
 sg13g2_nor2b_1 _6126_ (.A(net1363),
    .B_N(net1322),
    .Y(_2015_));
 sg13g2_a21o_1 _6127_ (.A2(_2014_),
    .A1(net1362),
    .B1(_2015_),
    .X(_2016_));
 sg13g2_nand2b_1 _6128_ (.Y(_2017_),
    .B(\s0.data_out[11][7] ),
    .A_N(net1380));
 sg13g2_a21oi_1 _6129_ (.A1(_1918_),
    .A2(_2017_),
    .Y(_2018_),
    .B1(net1374));
 sg13g2_a21oi_1 _6130_ (.A1(net1374),
    .A2(_2016_),
    .Y(_2019_),
    .B1(_2018_));
 sg13g2_a22oi_1 _6131_ (.Y(_2020_),
    .B1(_2019_),
    .B2(net1642),
    .A2(_2012_),
    .A1(net1652));
 sg13g2_nor2_1 _6132_ (.A(net1652),
    .B(_2012_),
    .Y(_2021_));
 sg13g2_or2_1 _6133_ (.X(_2022_),
    .B(_2019_),
    .A(net1642));
 sg13g2_nand3b_1 _6134_ (.B(_2022_),
    .C(_2020_),
    .Y(_2023_),
    .A_N(_2021_));
 sg13g2_nand2_1 _6135_ (.Y(_2024_),
    .A(net1366),
    .B(net605));
 sg13g2_mux2_1 _6136_ (.A0(\s0.data_out[12][5] ),
    .A1(\s0.data_out[11][5] ),
    .S(net1367),
    .X(_2025_));
 sg13g2_nor2b_1 _6137_ (.A(net1362),
    .B_N(net1332),
    .Y(_2026_));
 sg13g2_a21o_1 _6138_ (.A2(_2025_),
    .A1(net1362),
    .B1(_2026_),
    .X(_2027_));
 sg13g2_nand2b_1 _6139_ (.Y(_2028_),
    .B(net605),
    .A_N(net1380));
 sg13g2_a21oi_1 _6140_ (.A1(_1900_),
    .A2(_2028_),
    .Y(_2029_),
    .B1(net1373));
 sg13g2_a21oi_1 _6141_ (.A1(net1373),
    .A2(_2027_),
    .Y(_2030_),
    .B1(_2029_));
 sg13g2_nand2_1 _6142_ (.Y(_2031_),
    .A(net1662),
    .B(_2030_));
 sg13g2_o21ai_1 _6143_ (.B1(_2031_),
    .Y(_2032_),
    .A1(net1681),
    .A2(_2003_));
 sg13g2_nand2_1 _6144_ (.Y(_2033_),
    .A(net1364),
    .B(net788));
 sg13g2_mux2_1 _6145_ (.A0(\s0.data_out[12][4] ),
    .A1(\s0.data_out[11][4] ),
    .S(net1367),
    .X(_2034_));
 sg13g2_nor2b_1 _6146_ (.A(net1362),
    .B_N(net1337),
    .Y(_2035_));
 sg13g2_a21oi_1 _6147_ (.A1(net1362),
    .A2(_2034_),
    .Y(_2036_),
    .B1(_2035_));
 sg13g2_nand2b_1 _6148_ (.Y(_2037_),
    .B(net1373),
    .A_N(_2036_));
 sg13g2_o21ai_1 _6149_ (.B1(_1892_),
    .Y(_2038_),
    .A1(net1380),
    .A2(_3497_));
 sg13g2_nand2b_1 _6150_ (.Y(_2039_),
    .B(_2038_),
    .A_N(net1373));
 sg13g2_a21o_1 _6151_ (.A2(_2039_),
    .A1(_2037_),
    .B1(net1672),
    .X(_2040_));
 sg13g2_nand3_1 _6152_ (.B(_2037_),
    .C(_2039_),
    .A(net1673),
    .Y(_2041_));
 sg13g2_nor2_1 _6153_ (.A(net1662),
    .B(_2030_),
    .Y(_2042_));
 sg13g2_nor3_1 _6154_ (.A(_2023_),
    .B(_2032_),
    .C(_2042_),
    .Y(_2043_));
 sg13g2_nand4_1 _6155_ (.B(_2040_),
    .C(_2041_),
    .A(_2005_),
    .Y(_2044_),
    .D(_2043_));
 sg13g2_o21ai_1 _6156_ (.B1(_2031_),
    .Y(_2045_),
    .A1(_2041_),
    .A2(_2042_));
 sg13g2_nor2b_1 _6157_ (.A(_2023_),
    .B_N(_2045_),
    .Y(_2046_));
 sg13g2_nor2b_1 _6158_ (.A(_2020_),
    .B_N(_2022_),
    .Y(_2047_));
 sg13g2_nor3_1 _6159_ (.A(_1967_),
    .B(_2046_),
    .C(_2047_),
    .Y(_2048_));
 sg13g2_or2_1 _6160_ (.X(_2049_),
    .B(net1558),
    .A(net386));
 sg13g2_a21oi_1 _6161_ (.A1(_2044_),
    .A2(_2048_),
    .Y(_0292_),
    .B1(_2049_));
 sg13g2_and2_1 _6162_ (.A(net1358),
    .B(\s0.data_out[11][0] ),
    .X(_2050_));
 sg13g2_o21ai_1 _6163_ (.B1(net1368),
    .Y(_2051_),
    .A1(_1990_),
    .A2(_2050_));
 sg13g2_nand3_1 _6164_ (.B(_1994_),
    .C(_2051_),
    .A(net1729),
    .Y(_2052_));
 sg13g2_o21ai_1 _6165_ (.B1(_2052_),
    .Y(_2053_),
    .A1(net1729),
    .A2(net728));
 sg13g2_inv_1 _6166_ (.Y(_0293_),
    .A(_2053_));
 sg13g2_nor2_1 _6167_ (.A(_3383_),
    .B(_3492_),
    .Y(_2054_));
 sg13g2_o21ai_1 _6168_ (.B1(net1368),
    .Y(_2055_),
    .A1(_1982_),
    .A2(_2054_));
 sg13g2_nor2_1 _6169_ (.A(net1600),
    .B(_1987_),
    .Y(_2056_));
 sg13g2_a22oi_1 _6170_ (.Y(_0294_),
    .B1(_2055_),
    .B2(_2056_),
    .A2(_3491_),
    .A1(net1600));
 sg13g2_nor2_1 _6171_ (.A(_3383_),
    .B(_3494_),
    .Y(_2057_));
 sg13g2_o21ai_1 _6172_ (.B1(net1368),
    .Y(_2058_),
    .A1(_1976_),
    .A2(_2057_));
 sg13g2_nor2_1 _6173_ (.A(net1599),
    .B(_1979_),
    .Y(_2059_));
 sg13g2_a22oi_1 _6174_ (.Y(_0295_),
    .B1(_2058_),
    .B2(_2059_),
    .A2(_3490_),
    .A1(net1599));
 sg13g2_nor2_1 _6175_ (.A(_3383_),
    .B(_3493_),
    .Y(_2060_));
 sg13g2_o21ai_1 _6176_ (.B1(net1371),
    .Y(_2061_),
    .A1(_1999_),
    .A2(_2060_));
 sg13g2_nor2_1 _6177_ (.A(net1600),
    .B(_2002_),
    .Y(_2062_));
 sg13g2_a22oi_1 _6178_ (.Y(_0296_),
    .B1(_2061_),
    .B2(_2062_),
    .A2(_3489_),
    .A1(net1600));
 sg13g2_nor2_1 _6179_ (.A(_3383_),
    .B(_3497_),
    .Y(_2063_));
 sg13g2_o21ai_1 _6180_ (.B1(net1373),
    .Y(_2064_),
    .A1(_2035_),
    .A2(_2063_));
 sg13g2_nand3_1 _6181_ (.B(_2039_),
    .C(_2064_),
    .A(net1728),
    .Y(_2065_));
 sg13g2_o21ai_1 _6182_ (.B1(_2065_),
    .Y(_2066_),
    .A1(net1728),
    .A2(net453));
 sg13g2_inv_1 _6183_ (.Y(_0297_),
    .A(_2066_));
 sg13g2_nor2_1 _6184_ (.A(_3383_),
    .B(_3496_),
    .Y(_2067_));
 sg13g2_o21ai_1 _6185_ (.B1(net1373),
    .Y(_2068_),
    .A1(_2026_),
    .A2(_2067_));
 sg13g2_nor2_1 _6186_ (.A(net1602),
    .B(_2029_),
    .Y(_2069_));
 sg13g2_a22oi_1 _6187_ (.Y(_0298_),
    .B1(_2068_),
    .B2(_2069_),
    .A2(_3488_),
    .A1(net1601));
 sg13g2_and2_1 _6188_ (.A(net1363),
    .B(\s0.data_out[11][6] ),
    .X(_2070_));
 sg13g2_o21ai_1 _6189_ (.B1(net1374),
    .Y(_2071_),
    .A1(_2008_),
    .A2(_2070_));
 sg13g2_nand3b_1 _6190_ (.B(_2071_),
    .C(net1730),
    .Y(_2072_),
    .A_N(_2011_));
 sg13g2_o21ai_1 _6191_ (.B1(_2072_),
    .Y(_2073_),
    .A1(net1728),
    .A2(net709));
 sg13g2_inv_1 _6192_ (.Y(_0299_),
    .A(_2073_));
 sg13g2_nor2_1 _6193_ (.A(_3383_),
    .B(_3495_),
    .Y(_2074_));
 sg13g2_o21ai_1 _6194_ (.B1(net1374),
    .Y(_2075_),
    .A1(_2015_),
    .A2(_2074_));
 sg13g2_nor2_1 _6195_ (.A(net1602),
    .B(_2018_),
    .Y(_2076_));
 sg13g2_a22oi_1 _6196_ (.Y(_0300_),
    .B1(_2075_),
    .B2(_2076_),
    .A2(_3487_),
    .A1(net1602));
 sg13g2_o21ai_1 _6197_ (.B1(net1361),
    .Y(_2077_),
    .A1(net1318),
    .A2(net1630));
 sg13g2_nor2b_1 _6198_ (.A(net1630),
    .B_N(net1355),
    .Y(_2078_));
 sg13g2_or2_1 _6199_ (.X(_2079_),
    .B(_2078_),
    .A(_2077_));
 sg13g2_o21ai_1 _6200_ (.B1(_2079_),
    .Y(_2080_),
    .A1(net1361),
    .A2(_1964_));
 sg13g2_nor2_1 _6201_ (.A(net445),
    .B(_2080_),
    .Y(_2081_));
 sg13g2_nor2_1 _6202_ (.A(\s0.was_valid_out[10] [0]),
    .B(net1355),
    .Y(_2082_));
 sg13g2_nor2_1 _6203_ (.A(net1318),
    .B(_2077_),
    .Y(_2083_));
 sg13g2_o21ai_1 _6204_ (.B1(_3383_),
    .Y(_2084_),
    .A1(\s0.was_valid_out[10] [0]),
    .A2(net1366));
 sg13g2_o21ai_1 _6205_ (.B1(_2084_),
    .Y(_2085_),
    .A1(_2079_),
    .A2(_2082_));
 sg13g2_o21ai_1 _6206_ (.B1(net1728),
    .Y(_2086_),
    .A1(_2083_),
    .A2(_2085_));
 sg13g2_nor2_1 _6207_ (.A(_2081_),
    .B(_2086_),
    .Y(_0301_));
 sg13g2_nor2_1 _6208_ (.A(net1601),
    .B(_2080_),
    .Y(_0302_));
 sg13g2_and2_1 _6209_ (.A(net373),
    .B(net1726),
    .X(_0303_));
 sg13g2_nand2_1 _6210_ (.Y(_2087_),
    .A(net1352),
    .B(net479));
 sg13g2_mux2_1 _6211_ (.A0(\s0.data_out[11][2] ),
    .A1(\s0.data_out[10][2] ),
    .S(net1352),
    .X(_2088_));
 sg13g2_nor2b_1 _6212_ (.A(net1313),
    .B_N(net1343),
    .Y(_2089_));
 sg13g2_a21o_1 _6213_ (.A2(_2088_),
    .A1(net1313),
    .B1(_2089_),
    .X(_2090_));
 sg13g2_nand2b_1 _6214_ (.Y(_2091_),
    .B(net479),
    .A_N(net1364));
 sg13g2_a21oi_1 _6215_ (.A1(_1974_),
    .A2(_2091_),
    .Y(_2092_),
    .B1(net1357));
 sg13g2_a21oi_1 _6216_ (.A1(net1357),
    .A2(_2090_),
    .Y(_2093_),
    .B1(_2092_));
 sg13g2_or2_1 _6217_ (.X(_2094_),
    .B(_2093_),
    .A(net1686));
 sg13g2_nand2_1 _6218_ (.Y(_2095_),
    .A(net1352),
    .B(net659));
 sg13g2_o21ai_1 _6219_ (.B1(_2095_),
    .Y(_2096_),
    .A1(net1353),
    .A2(_3492_));
 sg13g2_nor2b_1 _6220_ (.A(net1313),
    .B_N(net1346),
    .Y(_2097_));
 sg13g2_a21o_1 _6221_ (.A2(_2096_),
    .A1(net1313),
    .B1(_2097_),
    .X(_2098_));
 sg13g2_nand2b_1 _6222_ (.Y(_2099_),
    .B(net659),
    .A_N(net1364));
 sg13g2_a21oi_1 _6223_ (.A1(_1983_),
    .A2(_2099_),
    .Y(_2100_),
    .B1(net1357));
 sg13g2_a21oi_1 _6224_ (.A1(net1357),
    .A2(_2098_),
    .Y(_2101_),
    .B1(_2100_));
 sg13g2_mux2_1 _6225_ (.A0(\s0.data_out[11][0] ),
    .A1(\s0.data_out[10][0] ),
    .S(net1353),
    .X(_2102_));
 sg13g2_nor2b_1 _6226_ (.A(net1313),
    .B_N(net1350),
    .Y(_2103_));
 sg13g2_a21oi_1 _6227_ (.A1(net1314),
    .A2(_2102_),
    .Y(_2104_),
    .B1(_2103_));
 sg13g2_nand2b_1 _6228_ (.Y(_2105_),
    .B(net1357),
    .A_N(_2104_));
 sg13g2_mux2_1 _6229_ (.A0(\s0.data_out[10][0] ),
    .A1(\s0.data_out[11][0] ),
    .S(net1364),
    .X(_2106_));
 sg13g2_nand2_1 _6230_ (.Y(_2107_),
    .A(_3383_),
    .B(_2106_));
 sg13g2_a221oi_1 _6231_ (.B2(_2107_),
    .C1(net1701),
    .B1(_2105_),
    .A1(net1697),
    .Y(_2108_),
    .A2(_2101_));
 sg13g2_o21ai_1 _6232_ (.B1(_2094_),
    .Y(_2109_),
    .A1(net1697),
    .A2(_2101_));
 sg13g2_nand2_1 _6233_ (.Y(_2110_),
    .A(net1353),
    .B(net436));
 sg13g2_o21ai_1 _6234_ (.B1(_2110_),
    .Y(_2111_),
    .A1(net1353),
    .A2(_3493_));
 sg13g2_nor2_1 _6235_ (.A(net1314),
    .B(net1161),
    .Y(_2112_));
 sg13g2_a21o_1 _6236_ (.A2(_2111_),
    .A1(net1314),
    .B1(_2112_),
    .X(_2113_));
 sg13g2_nand2b_1 _6237_ (.Y(_2114_),
    .B(net436),
    .A_N(net1365));
 sg13g2_a21oi_1 _6238_ (.A1(_1997_),
    .A2(_2114_),
    .Y(_2115_),
    .B1(net1358));
 sg13g2_a21oi_1 _6239_ (.A1(net1358),
    .A2(_2113_),
    .Y(_2116_),
    .B1(_2115_));
 sg13g2_a22oi_1 _6240_ (.Y(_2117_),
    .B1(_2116_),
    .B2(net1678),
    .A2(_2093_),
    .A1(net1686));
 sg13g2_o21ai_1 _6241_ (.B1(_2117_),
    .Y(_2118_),
    .A1(_2108_),
    .A2(_2109_));
 sg13g2_nand2_1 _6242_ (.Y(_2119_),
    .A(net1354),
    .B(net626));
 sg13g2_mux2_1 _6243_ (.A0(\s0.data_out[11][6] ),
    .A1(\s0.data_out[10][6] ),
    .S(net1354),
    .X(_2120_));
 sg13g2_nor2b_1 _6244_ (.A(net1318),
    .B_N(net1327),
    .Y(_2121_));
 sg13g2_a21o_1 _6245_ (.A2(_2120_),
    .A1(net1317),
    .B1(_2121_),
    .X(_2122_));
 sg13g2_nand2b_1 _6246_ (.Y(_2123_),
    .B(net626),
    .A_N(net1366));
 sg13g2_a21oi_1 _6247_ (.A1(_2006_),
    .A2(_2123_),
    .Y(_2124_),
    .B1(net1360));
 sg13g2_a21oi_1 _6248_ (.A1(net1360),
    .A2(_2122_),
    .Y(_2125_),
    .B1(_2124_));
 sg13g2_nand2_1 _6249_ (.Y(_2126_),
    .A(net1354),
    .B(net514));
 sg13g2_mux2_1 _6250_ (.A0(\s0.data_out[11][7] ),
    .A1(\s0.data_out[10][7] ),
    .S(net1355),
    .X(_2127_));
 sg13g2_nor2b_1 _6251_ (.A(net1318),
    .B_N(net1322),
    .Y(_2128_));
 sg13g2_a21o_1 _6252_ (.A2(_2127_),
    .A1(net1318),
    .B1(_2128_),
    .X(_2129_));
 sg13g2_nand2b_1 _6253_ (.Y(_2130_),
    .B(net514),
    .A_N(net1366));
 sg13g2_a21oi_1 _6254_ (.A1(_2013_),
    .A2(_2130_),
    .Y(_2131_),
    .B1(net1360));
 sg13g2_a21oi_1 _6255_ (.A1(net1360),
    .A2(_2129_),
    .Y(_2132_),
    .B1(_2131_));
 sg13g2_a22oi_1 _6256_ (.Y(_2133_),
    .B1(_2132_),
    .B2(net1641),
    .A2(_2125_),
    .A1(net1651));
 sg13g2_inv_1 _6257_ (.Y(_2134_),
    .A(_2133_));
 sg13g2_nor2_1 _6258_ (.A(net1651),
    .B(_2125_),
    .Y(_2135_));
 sg13g2_or2_1 _6259_ (.X(_2136_),
    .B(_2132_),
    .A(net1641));
 sg13g2_nand3b_1 _6260_ (.B(_2136_),
    .C(_2133_),
    .Y(_2137_),
    .A_N(_2135_));
 sg13g2_mux2_1 _6261_ (.A0(\s0.data_out[11][4] ),
    .A1(\s0.data_out[10][4] ),
    .S(net1353),
    .X(_2138_));
 sg13g2_nor2b_1 _6262_ (.A(net1317),
    .B_N(net1338),
    .Y(_2139_));
 sg13g2_a21o_1 _6263_ (.A2(_2138_),
    .A1(net1317),
    .B1(_2139_),
    .X(_2140_));
 sg13g2_nand2b_1 _6264_ (.Y(_2141_),
    .B(net402),
    .A_N(net1364));
 sg13g2_a21oi_1 _6265_ (.A1(_2033_),
    .A2(_2141_),
    .Y(_2142_),
    .B1(net1358));
 sg13g2_a21oi_1 _6266_ (.A1(net1360),
    .A2(_2140_),
    .Y(_2143_),
    .B1(_2142_));
 sg13g2_and2_1 _6267_ (.A(net1670),
    .B(_2143_),
    .X(_2144_));
 sg13g2_nand2_1 _6268_ (.Y(_2145_),
    .A(net1354),
    .B(net497));
 sg13g2_mux2_1 _6269_ (.A0(\s0.data_out[11][5] ),
    .A1(\s0.data_out[10][5] ),
    .S(net1355),
    .X(_2146_));
 sg13g2_nor2b_1 _6270_ (.A(net1317),
    .B_N(net1332),
    .Y(_2147_));
 sg13g2_a21o_1 _6271_ (.A2(_2146_),
    .A1(net1317),
    .B1(_2147_),
    .X(_2148_));
 sg13g2_nand2b_1 _6272_ (.Y(_2149_),
    .B(net497),
    .A_N(net1366));
 sg13g2_a21oi_1 _6273_ (.A1(_2024_),
    .A2(_2149_),
    .Y(_2150_),
    .B1(net1360));
 sg13g2_a21oi_1 _6274_ (.A1(net1360),
    .A2(_2148_),
    .Y(_2151_),
    .B1(_2150_));
 sg13g2_a21o_1 _6275_ (.A2(_2151_),
    .A1(net1660),
    .B1(_2144_),
    .X(_2152_));
 sg13g2_or2_1 _6276_ (.X(_2153_),
    .B(_2151_),
    .A(net1660));
 sg13g2_o21ai_1 _6277_ (.B1(_2153_),
    .Y(_2154_),
    .A1(net1670),
    .A2(_2143_));
 sg13g2_nor2_1 _6278_ (.A(net1681),
    .B(_2116_),
    .Y(_2155_));
 sg13g2_nor4_1 _6279_ (.A(_2137_),
    .B(_2152_),
    .C(_2154_),
    .D(_2155_),
    .Y(_2156_));
 sg13g2_nand2_1 _6280_ (.Y(_2157_),
    .A(_2118_),
    .B(_2156_));
 sg13g2_nor2b_1 _6281_ (.A(_2137_),
    .B_N(_2152_),
    .Y(_2158_));
 sg13g2_a221oi_1 _6282_ (.B2(_2158_),
    .C1(_2080_),
    .B1(_2153_),
    .A1(_2134_),
    .Y(_2159_),
    .A2(_2136_));
 sg13g2_or2_1 _6283_ (.X(_2160_),
    .B(net1558),
    .A(net385));
 sg13g2_a21oi_1 _6284_ (.A1(_2157_),
    .A2(_2159_),
    .Y(_0304_),
    .B1(_2160_));
 sg13g2_and2_1 _6285_ (.A(net1313),
    .B(net840),
    .X(_2161_));
 sg13g2_o21ai_1 _6286_ (.B1(net1357),
    .Y(_2162_),
    .A1(_2103_),
    .A2(_2161_));
 sg13g2_nand3_1 _6287_ (.B(_2107_),
    .C(_2162_),
    .A(net1729),
    .Y(_2163_));
 sg13g2_o21ai_1 _6288_ (.B1(_2163_),
    .Y(_2164_),
    .A1(net1729),
    .A2(net650));
 sg13g2_inv_1 _6289_ (.Y(_0305_),
    .A(_2164_));
 sg13g2_and2_1 _6290_ (.A(net1313),
    .B(net659),
    .X(_2165_));
 sg13g2_o21ai_1 _6291_ (.B1(net1357),
    .Y(_2166_),
    .A1(_2097_),
    .A2(_2165_));
 sg13g2_nor2_1 _6292_ (.A(net1599),
    .B(_2100_),
    .Y(_2167_));
 sg13g2_a22oi_1 _6293_ (.Y(_0306_),
    .B1(_2166_),
    .B2(_2167_),
    .A2(_3492_),
    .A1(net1599));
 sg13g2_and2_1 _6294_ (.A(net1313),
    .B(net479),
    .X(_2168_));
 sg13g2_o21ai_1 _6295_ (.B1(net1357),
    .Y(_2169_),
    .A1(_2089_),
    .A2(_2168_));
 sg13g2_nor2_1 _6296_ (.A(net1599),
    .B(_2092_),
    .Y(_2170_));
 sg13g2_a22oi_1 _6297_ (.Y(_0307_),
    .B1(_2169_),
    .B2(_2170_),
    .A2(_3494_),
    .A1(net1599));
 sg13g2_and2_1 _6298_ (.A(net1314),
    .B(net436),
    .X(_2171_));
 sg13g2_o21ai_1 _6299_ (.B1(net1358),
    .Y(_2172_),
    .A1(_2112_),
    .A2(_2171_));
 sg13g2_nor2_1 _6300_ (.A(net1599),
    .B(net437),
    .Y(_2173_));
 sg13g2_a22oi_1 _6301_ (.Y(_0308_),
    .B1(_2172_),
    .B2(_2173_),
    .A2(_3493_),
    .A1(net1599));
 sg13g2_and2_1 _6302_ (.A(net1314),
    .B(net402),
    .X(_2174_));
 sg13g2_o21ai_1 _6303_ (.B1(net1358),
    .Y(_2175_),
    .A1(_2139_),
    .A2(_2174_));
 sg13g2_nor2_1 _6304_ (.A(net1601),
    .B(_2142_),
    .Y(_2176_));
 sg13g2_a22oi_1 _6305_ (.Y(_0309_),
    .B1(_2175_),
    .B2(_2176_),
    .A2(_3497_),
    .A1(net1601));
 sg13g2_and2_1 _6306_ (.A(net1317),
    .B(net497),
    .X(_2177_));
 sg13g2_o21ai_1 _6307_ (.B1(net1360),
    .Y(_2178_),
    .A1(_2147_),
    .A2(_2177_));
 sg13g2_nor2_1 _6308_ (.A(net1601),
    .B(_2150_),
    .Y(_2179_));
 sg13g2_a22oi_1 _6309_ (.Y(_0310_),
    .B1(_2178_),
    .B2(_2179_),
    .A2(_3496_),
    .A1(net1601));
 sg13g2_and2_1 _6310_ (.A(net1317),
    .B(\s0.data_out[10][6] ),
    .X(_2180_));
 sg13g2_o21ai_1 _6311_ (.B1(net1361),
    .Y(_2181_),
    .A1(_2121_),
    .A2(_2180_));
 sg13g2_nand3b_1 _6312_ (.B(_2181_),
    .C(net1728),
    .Y(_2182_),
    .A_N(_2124_));
 sg13g2_o21ai_1 _6313_ (.B1(_2182_),
    .Y(_2183_),
    .A1(net1728),
    .A2(net718));
 sg13g2_inv_1 _6314_ (.Y(_0311_),
    .A(net719));
 sg13g2_and2_1 _6315_ (.A(net1317),
    .B(net514),
    .X(_2184_));
 sg13g2_o21ai_1 _6316_ (.B1(net1361),
    .Y(_2185_),
    .A1(_2128_),
    .A2(_2184_));
 sg13g2_nor2_1 _6317_ (.A(net1601),
    .B(_2131_),
    .Y(_2186_));
 sg13g2_a22oi_1 _6318_ (.Y(_0312_),
    .B1(_2185_),
    .B2(_2186_),
    .A2(_3495_),
    .A1(net1601));
 sg13g2_o21ai_1 _6319_ (.B1(net1315),
    .Y(_2187_),
    .A1(net1631),
    .A2(net1303));
 sg13g2_nor2b_1 _6320_ (.A(net1631),
    .B_N(net1308),
    .Y(_2188_));
 sg13g2_nor2_1 _6321_ (.A(_2187_),
    .B(_2188_),
    .Y(_2189_));
 sg13g2_inv_1 _6322_ (.Y(_2190_),
    .A(_2189_));
 sg13g2_o21ai_1 _6323_ (.B1(_2189_),
    .Y(_2191_),
    .A1(net447),
    .A2(net1309));
 sg13g2_nor2_1 _6324_ (.A(net1303),
    .B(_2187_),
    .Y(_2192_));
 sg13g2_nor2_1 _6325_ (.A(net447),
    .B(net1354),
    .Y(_2193_));
 sg13g2_o21ai_1 _6326_ (.B1(_2191_),
    .Y(_2194_),
    .A1(net1315),
    .A2(_2193_));
 sg13g2_o21ai_1 _6327_ (.B1(_2190_),
    .Y(_2195_),
    .A1(net1315),
    .A2(_2078_));
 sg13g2_nor2_1 _6328_ (.A(net452),
    .B(_2195_),
    .Y(_2196_));
 sg13g2_o21ai_1 _6329_ (.B1(net1727),
    .Y(_2197_),
    .A1(_2192_),
    .A2(_2194_));
 sg13g2_nor2_1 _6330_ (.A(_2196_),
    .B(_2197_),
    .Y(_0313_));
 sg13g2_nor2_1 _6331_ (.A(net1598),
    .B(_2195_),
    .Y(_0314_));
 sg13g2_nor2_1 _6332_ (.A(net1626),
    .B(net1348),
    .Y(_2198_));
 sg13g2_a21oi_1 _6333_ (.A1(net1626),
    .A2(net1559),
    .Y(_0315_),
    .B1(_2198_));
 sg13g2_nor2_1 _6334_ (.A(net1626),
    .B(net1344),
    .Y(_2199_));
 sg13g2_a21oi_1 _6335_ (.A1(net1626),
    .A2(_3415_),
    .Y(_0316_),
    .B1(_2199_));
 sg13g2_nor2_1 _6336_ (.A(net1625),
    .B(net1340),
    .Y(_2200_));
 sg13g2_a21oi_1 _6337_ (.A1(net1625),
    .A2(net1560),
    .Y(_0317_),
    .B1(_2200_));
 sg13g2_nand2_1 _6338_ (.Y(_2201_),
    .A(net1625),
    .B(net1677));
 sg13g2_o21ai_1 _6339_ (.B1(_2201_),
    .Y(_0318_),
    .A1(net1625),
    .A2(net1160));
 sg13g2_nor2_1 _6340_ (.A(net1625),
    .B(net1335),
    .Y(_2202_));
 sg13g2_a21oi_1 _6341_ (.A1(net1625),
    .A2(_3406_),
    .Y(_0319_),
    .B1(_2202_));
 sg13g2_nor2_1 _6342_ (.A(net1625),
    .B(net1330),
    .Y(_2203_));
 sg13g2_a21oi_1 _6343_ (.A1(net1625),
    .A2(_3403_),
    .Y(_0320_),
    .B1(_2203_));
 sg13g2_nor2_1 _6344_ (.A(net1626),
    .B(net1325),
    .Y(_2204_));
 sg13g2_a21oi_1 _6345_ (.A1(net1626),
    .A2(_3402_),
    .Y(_0321_),
    .B1(_2204_));
 sg13g2_mux2_1 _6346_ (.A0(net1320),
    .A1(net1636),
    .S(net1),
    .X(_0322_));
 sg13g2_nand2_1 _6347_ (.Y(_2205_),
    .A(net1306),
    .B(net490));
 sg13g2_mux2_1 _6348_ (.A0(\s0.data_out[10][2] ),
    .A1(\s0.data_out[9][2] ),
    .S(net1307),
    .X(_2206_));
 sg13g2_nor2b_1 _6349_ (.A(net1300),
    .B_N(net1343),
    .Y(_2207_));
 sg13g2_a21o_1 _6350_ (.A2(_2206_),
    .A1(net1300),
    .B1(_2207_),
    .X(_2208_));
 sg13g2_nand2b_1 _6351_ (.Y(_2209_),
    .B(\s0.data_out[9][2] ),
    .A_N(net1352));
 sg13g2_a21oi_1 _6352_ (.A1(_2087_),
    .A2(_2209_),
    .Y(_2210_),
    .B1(net1311));
 sg13g2_a21oi_1 _6353_ (.A1(net1311),
    .A2(_2208_),
    .Y(_2211_),
    .B1(_2210_));
 sg13g2_or2_1 _6354_ (.X(_2212_),
    .B(_2211_),
    .A(net1688));
 sg13g2_nor2b_1 _6355_ (.A(net1300),
    .B_N(net1347),
    .Y(_2213_));
 sg13g2_nand2_1 _6356_ (.Y(_2214_),
    .A(net1306),
    .B(net475));
 sg13g2_o21ai_1 _6357_ (.B1(_2214_),
    .Y(_2215_),
    .A1(net1307),
    .A2(_3498_));
 sg13g2_a21o_1 _6358_ (.A2(_2215_),
    .A1(net1300),
    .B1(_2213_),
    .X(_2216_));
 sg13g2_nand2b_1 _6359_ (.Y(_2217_),
    .B(net475),
    .A_N(net1352));
 sg13g2_a21oi_1 _6360_ (.A1(_2095_),
    .A2(_2217_),
    .Y(_2218_),
    .B1(net1311));
 sg13g2_a21oi_1 _6361_ (.A1(net1311),
    .A2(_2216_),
    .Y(_2219_),
    .B1(_2218_));
 sg13g2_mux2_1 _6362_ (.A0(\s0.data_out[10][0] ),
    .A1(\s0.data_out[9][0] ),
    .S(net1307),
    .X(_2220_));
 sg13g2_nor2b_1 _6363_ (.A(net1301),
    .B_N(net1351),
    .Y(_2221_));
 sg13g2_a21oi_1 _6364_ (.A1(net1300),
    .A2(_2220_),
    .Y(_2222_),
    .B1(_2221_));
 sg13g2_nand2b_1 _6365_ (.Y(_2223_),
    .B(net1311),
    .A_N(_2222_));
 sg13g2_mux2_1 _6366_ (.A0(\s0.data_out[9][0] ),
    .A1(\s0.data_out[10][0] ),
    .S(net1352),
    .X(_2224_));
 sg13g2_nand2b_1 _6367_ (.Y(_2225_),
    .B(_2224_),
    .A_N(net1311));
 sg13g2_o21ai_1 _6368_ (.B1(_2212_),
    .Y(_2226_),
    .A1(net1694),
    .A2(_2219_));
 sg13g2_a221oi_1 _6369_ (.B2(_2225_),
    .C1(net1701),
    .B1(_2223_),
    .A1(net1694),
    .Y(_2227_),
    .A2(_2219_));
 sg13g2_nand2_1 _6370_ (.Y(_2228_),
    .A(net1307),
    .B(net664));
 sg13g2_o21ai_1 _6371_ (.B1(_2228_),
    .Y(_2229_),
    .A1(net1307),
    .A2(_3499_));
 sg13g2_nor2_1 _6372_ (.A(net1301),
    .B(net1161),
    .Y(_2230_));
 sg13g2_a21o_1 _6373_ (.A2(_2229_),
    .A1(net1301),
    .B1(_2230_),
    .X(_2231_));
 sg13g2_nand2b_1 _6374_ (.Y(_2232_),
    .B(net664),
    .A_N(net1352));
 sg13g2_a21oi_1 _6375_ (.A1(_2110_),
    .A2(_2232_),
    .Y(_2233_),
    .B1(net1312));
 sg13g2_a21oi_1 _6376_ (.A1(net1312),
    .A2(_2231_),
    .Y(_2234_),
    .B1(_2233_));
 sg13g2_a22oi_1 _6377_ (.Y(_2235_),
    .B1(_2234_),
    .B2(net1678),
    .A2(_2211_),
    .A1(net1688));
 sg13g2_o21ai_1 _6378_ (.B1(_2235_),
    .Y(_2236_),
    .A1(_2226_),
    .A2(_2227_));
 sg13g2_nand2_1 _6379_ (.Y(_2237_),
    .A(net1308),
    .B(net534));
 sg13g2_mux2_1 _6380_ (.A0(\s0.data_out[10][7] ),
    .A1(\s0.data_out[9][7] ),
    .S(net1309),
    .X(_2238_));
 sg13g2_nor2b_1 _6381_ (.A(net1303),
    .B_N(net1322),
    .Y(_2239_));
 sg13g2_a21o_1 _6382_ (.A2(_2238_),
    .A1(net1303),
    .B1(_2239_),
    .X(_2240_));
 sg13g2_nand2b_1 _6383_ (.Y(_2241_),
    .B(\s0.data_out[9][7] ),
    .A_N(net1354));
 sg13g2_a21oi_1 _6384_ (.A1(_2126_),
    .A2(_2241_),
    .Y(_2242_),
    .B1(net1315));
 sg13g2_a21oi_1 _6385_ (.A1(net1315),
    .A2(_2240_),
    .Y(_2243_),
    .B1(_2242_));
 sg13g2_nand2_1 _6386_ (.Y(_2244_),
    .A(net1308),
    .B(net735));
 sg13g2_mux2_1 _6387_ (.A0(\s0.data_out[10][6] ),
    .A1(\s0.data_out[9][6] ),
    .S(net1309),
    .X(_2245_));
 sg13g2_nor2b_1 _6388_ (.A(net1303),
    .B_N(net1327),
    .Y(_2246_));
 sg13g2_a21o_1 _6389_ (.A2(_2245_),
    .A1(net1303),
    .B1(_2246_),
    .X(_2247_));
 sg13g2_nand2b_1 _6390_ (.Y(_2248_),
    .B(net837),
    .A_N(net1354));
 sg13g2_a21oi_1 _6391_ (.A1(_2119_),
    .A2(_2248_),
    .Y(_2249_),
    .B1(net1315));
 sg13g2_a21oi_1 _6392_ (.A1(net1316),
    .A2(_2247_),
    .Y(_2250_),
    .B1(_2249_));
 sg13g2_a22oi_1 _6393_ (.Y(_2251_),
    .B1(_2250_),
    .B2(net1651),
    .A2(_2243_),
    .A1(net1641));
 sg13g2_nor2_1 _6394_ (.A(net1651),
    .B(_2250_),
    .Y(_2252_));
 sg13g2_or2_1 _6395_ (.X(_2253_),
    .B(_2243_),
    .A(net1645));
 sg13g2_nand3b_1 _6396_ (.B(_2253_),
    .C(_2251_),
    .Y(_2254_),
    .A_N(_2252_));
 sg13g2_nand2_1 _6397_ (.Y(_2255_),
    .A(net1306),
    .B(\s0.data_out[9][4] ));
 sg13g2_mux2_1 _6398_ (.A0(\s0.data_out[10][4] ),
    .A1(\s0.data_out[9][4] ),
    .S(net1307),
    .X(_2256_));
 sg13g2_nor2b_1 _6399_ (.A(net1301),
    .B_N(net1338),
    .Y(_2257_));
 sg13g2_a21oi_1 _6400_ (.A1(net1301),
    .A2(_2256_),
    .Y(_2258_),
    .B1(_2257_));
 sg13g2_nand2b_1 _6401_ (.Y(_2259_),
    .B(net1312),
    .A_N(_2258_));
 sg13g2_mux2_1 _6402_ (.A0(\s0.data_out[9][4] ),
    .A1(\s0.data_out[10][4] ),
    .S(net1352),
    .X(_2260_));
 sg13g2_nand2b_1 _6403_ (.Y(_2261_),
    .B(_2260_),
    .A_N(net1312));
 sg13g2_nand3_1 _6404_ (.B(_2259_),
    .C(_2261_),
    .A(net1670),
    .Y(_2262_));
 sg13g2_nand2_1 _6405_ (.Y(_2263_),
    .A(net1308),
    .B(\s0.data_out[9][5] ));
 sg13g2_mux2_1 _6406_ (.A0(\s0.data_out[10][5] ),
    .A1(\s0.data_out[9][5] ),
    .S(net1309),
    .X(_2264_));
 sg13g2_nor2b_1 _6407_ (.A(net1304),
    .B_N(net1332),
    .Y(_2265_));
 sg13g2_a21o_1 _6408_ (.A2(_2264_),
    .A1(net1304),
    .B1(_2265_),
    .X(_2266_));
 sg13g2_nand2b_1 _6409_ (.Y(_2267_),
    .B(\s0.data_out[9][5] ),
    .A_N(net1354));
 sg13g2_a21oi_1 _6410_ (.A1(_2145_),
    .A2(_2267_),
    .Y(_2268_),
    .B1(net1316));
 sg13g2_a21oi_1 _6411_ (.A1(net1316),
    .A2(_2266_),
    .Y(_2269_),
    .B1(_2268_));
 sg13g2_nor2_1 _6412_ (.A(net1660),
    .B(_2269_),
    .Y(_2270_));
 sg13g2_nand2_1 _6413_ (.Y(_2271_),
    .A(net1660),
    .B(_2269_));
 sg13g2_a21o_1 _6414_ (.A2(_2261_),
    .A1(_2259_),
    .B1(net1670),
    .X(_2272_));
 sg13g2_o21ai_1 _6415_ (.B1(_2271_),
    .Y(_2273_),
    .A1(net1679),
    .A2(_2234_));
 sg13g2_nor3_1 _6416_ (.A(_2254_),
    .B(_2270_),
    .C(_2273_),
    .Y(_2274_));
 sg13g2_nand4_1 _6417_ (.B(_2262_),
    .C(_2272_),
    .A(_2236_),
    .Y(_2275_),
    .D(_2274_));
 sg13g2_o21ai_1 _6418_ (.B1(_2271_),
    .Y(_2276_),
    .A1(_2262_),
    .A2(_2270_));
 sg13g2_nor2b_1 _6419_ (.A(_2254_),
    .B_N(_2276_),
    .Y(_2277_));
 sg13g2_nor2b_1 _6420_ (.A(_2251_),
    .B_N(_2253_),
    .Y(_2278_));
 sg13g2_nor3_1 _6421_ (.A(_2195_),
    .B(_2277_),
    .C(_2278_),
    .Y(_2279_));
 sg13g2_or2_1 _6422_ (.X(_2280_),
    .B(net1558),
    .A(net373));
 sg13g2_a21oi_1 _6423_ (.A1(_2275_),
    .A2(_2279_),
    .Y(_0323_),
    .B1(_2280_));
 sg13g2_and2_1 _6424_ (.A(net1300),
    .B(\s0.data_out[9][0] ),
    .X(_2281_));
 sg13g2_o21ai_1 _6425_ (.B1(net1311),
    .Y(_2282_),
    .A1(_2221_),
    .A2(_2281_));
 sg13g2_nand3_1 _6426_ (.B(_2225_),
    .C(_2282_),
    .A(net1726),
    .Y(_2283_));
 sg13g2_o21ai_1 _6427_ (.B1(_2283_),
    .Y(_2284_),
    .A1(net1726),
    .A2(net705));
 sg13g2_inv_1 _6428_ (.Y(_0324_),
    .A(_2284_));
 sg13g2_and2_1 _6429_ (.A(net1300),
    .B(net475),
    .X(_2285_));
 sg13g2_o21ai_1 _6430_ (.B1(net1311),
    .Y(_2286_),
    .A1(_2213_),
    .A2(_2285_));
 sg13g2_nor2_1 _6431_ (.A(net1597),
    .B(_2218_),
    .Y(_2287_));
 sg13g2_a22oi_1 _6432_ (.Y(_0325_),
    .B1(_2286_),
    .B2(_2287_),
    .A2(_3498_),
    .A1(net1597));
 sg13g2_and2_1 _6433_ (.A(net1300),
    .B(\s0.data_out[9][2] ),
    .X(_2288_));
 sg13g2_o21ai_1 _6434_ (.B1(net1312),
    .Y(_2289_),
    .A1(_2207_),
    .A2(_2288_));
 sg13g2_nor2_1 _6435_ (.A(net1596),
    .B(_2210_),
    .Y(_2290_));
 sg13g2_a22oi_1 _6436_ (.Y(_0326_),
    .B1(_2289_),
    .B2(_2290_),
    .A2(_3500_),
    .A1(net1596));
 sg13g2_and2_1 _6437_ (.A(net1301),
    .B(net664),
    .X(_2291_));
 sg13g2_o21ai_1 _6438_ (.B1(net1312),
    .Y(_2292_),
    .A1(_2230_),
    .A2(net665));
 sg13g2_nor2_1 _6439_ (.A(net1597),
    .B(_2233_),
    .Y(_2293_));
 sg13g2_a22oi_1 _6440_ (.Y(_0327_),
    .B1(net666),
    .B2(_2293_),
    .A2(_3499_),
    .A1(net1597));
 sg13g2_and2_1 _6441_ (.A(net1301),
    .B(\s0.data_out[9][4] ),
    .X(_2294_));
 sg13g2_o21ai_1 _6442_ (.B1(net1312),
    .Y(_2295_),
    .A1(_2257_),
    .A2(_2294_));
 sg13g2_nand3_1 _6443_ (.B(_2261_),
    .C(_2295_),
    .A(net1726),
    .Y(_2296_));
 sg13g2_o21ai_1 _6444_ (.B1(_2296_),
    .Y(_2297_),
    .A1(net1726),
    .A2(net402));
 sg13g2_inv_1 _6445_ (.Y(_0328_),
    .A(_2297_));
 sg13g2_and2_1 _6446_ (.A(net1304),
    .B(\s0.data_out[9][5] ),
    .X(_2298_));
 sg13g2_o21ai_1 _6447_ (.B1(net1316),
    .Y(_2299_),
    .A1(_2265_),
    .A2(_2298_));
 sg13g2_nor2_1 _6448_ (.A(net1598),
    .B(_2268_),
    .Y(_2300_));
 sg13g2_a22oi_1 _6449_ (.Y(_0329_),
    .B1(_2299_),
    .B2(_2300_),
    .A2(_3502_),
    .A1(net1598));
 sg13g2_and2_1 _6450_ (.A(net1304),
    .B(\s0.data_out[9][6] ),
    .X(_2301_));
 sg13g2_o21ai_1 _6451_ (.B1(net1315),
    .Y(_2302_),
    .A1(_2246_),
    .A2(_2301_));
 sg13g2_nand3b_1 _6452_ (.B(_2302_),
    .C(net1727),
    .Y(_2303_),
    .A_N(_2249_));
 sg13g2_o21ai_1 _6453_ (.B1(_2303_),
    .Y(_2304_),
    .A1(net1726),
    .A2(net626));
 sg13g2_inv_1 _6454_ (.Y(_0330_),
    .A(_2304_));
 sg13g2_and2_1 _6455_ (.A(net1303),
    .B(\s0.data_out[9][7] ),
    .X(_2305_));
 sg13g2_o21ai_1 _6456_ (.B1(net1315),
    .Y(_2306_),
    .A1(_2239_),
    .A2(_2305_));
 sg13g2_nor2_1 _6457_ (.A(net1598),
    .B(_2242_),
    .Y(_2307_));
 sg13g2_a22oi_1 _6458_ (.Y(_0331_),
    .B1(_2306_),
    .B2(_2307_),
    .A2(_3501_),
    .A1(net1598));
 sg13g2_o21ai_1 _6459_ (.B1(net1305),
    .Y(_2308_),
    .A1(net1631),
    .A2(net1292));
 sg13g2_nor2b_1 _6460_ (.A(net1629),
    .B_N(net1296),
    .Y(_2309_));
 sg13g2_nor2_1 _6461_ (.A(_2308_),
    .B(_2309_),
    .Y(_2310_));
 sg13g2_inv_1 _6462_ (.Y(_2311_),
    .A(_2310_));
 sg13g2_o21ai_1 _6463_ (.B1(_2311_),
    .Y(_2312_),
    .A1(net1303),
    .A2(_2188_));
 sg13g2_nor2_1 _6464_ (.A(net447),
    .B(_2312_),
    .Y(_2313_));
 sg13g2_o21ai_1 _6465_ (.B1(_2310_),
    .Y(_2314_),
    .A1(\s0.was_valid_out[8] [0]),
    .A2(net1297));
 sg13g2_nor2_1 _6466_ (.A(net1292),
    .B(_2308_),
    .Y(_2315_));
 sg13g2_nor2_1 _6467_ (.A(\s0.was_valid_out[8] [0]),
    .B(net1308),
    .Y(_2316_));
 sg13g2_o21ai_1 _6468_ (.B1(_2314_),
    .Y(_2317_),
    .A1(net1305),
    .A2(_2316_));
 sg13g2_o21ai_1 _6469_ (.B1(net1727),
    .Y(_2318_),
    .A1(_2315_),
    .A2(_2317_));
 sg13g2_nor2_1 _6470_ (.A(_2313_),
    .B(_2318_),
    .Y(_0332_));
 sg13g2_nor2_1 _6471_ (.A(net1603),
    .B(_2312_),
    .Y(_0333_));
 sg13g2_and2_1 _6472_ (.A(net1720),
    .B(net391),
    .X(_0334_));
 sg13g2_nand2_1 _6473_ (.Y(_2319_),
    .A(net1294),
    .B(net562));
 sg13g2_mux2_1 _6474_ (.A0(\s0.data_out[9][2] ),
    .A1(\s0.data_out[8][2] ),
    .S(net1294),
    .X(_2320_));
 sg13g2_nor2b_1 _6475_ (.A(net1288),
    .B_N(net1343),
    .Y(_2321_));
 sg13g2_a21o_1 _6476_ (.A2(_2320_),
    .A1(net1288),
    .B1(_2321_),
    .X(_2322_));
 sg13g2_nand2b_1 _6477_ (.Y(_2323_),
    .B(\s0.data_out[8][2] ),
    .A_N(net1306));
 sg13g2_a21oi_1 _6478_ (.A1(_2205_),
    .A2(_2323_),
    .Y(_2324_),
    .B1(net1298));
 sg13g2_a21oi_1 _6479_ (.A1(net1298),
    .A2(_2322_),
    .Y(_2325_),
    .B1(_2324_));
 sg13g2_nor2_1 _6480_ (.A(net1688),
    .B(_2325_),
    .Y(_2326_));
 sg13g2_nand2_1 _6481_ (.Y(_2327_),
    .A(net1294),
    .B(net594));
 sg13g2_mux2_1 _6482_ (.A0(\s0.data_out[9][1] ),
    .A1(\s0.data_out[8][1] ),
    .S(net1294),
    .X(_2328_));
 sg13g2_nor2b_1 _6483_ (.A(net1288),
    .B_N(net1347),
    .Y(_2329_));
 sg13g2_a21o_1 _6484_ (.A2(_2328_),
    .A1(net1288),
    .B1(_2329_),
    .X(_2330_));
 sg13g2_nand2b_1 _6485_ (.Y(_2331_),
    .B(\s0.data_out[8][1] ),
    .A_N(net1306));
 sg13g2_a21oi_1 _6486_ (.A1(_2214_),
    .A2(_2331_),
    .Y(_2332_),
    .B1(net1298));
 sg13g2_a21oi_1 _6487_ (.A1(net1299),
    .A2(_2330_),
    .Y(_2333_),
    .B1(_2332_));
 sg13g2_mux2_1 _6488_ (.A0(\s0.data_out[9][0] ),
    .A1(\s0.data_out[8][0] ),
    .S(net1294),
    .X(_2334_));
 sg13g2_nor2b_1 _6489_ (.A(net1288),
    .B_N(net1351),
    .Y(_2335_));
 sg13g2_a21oi_1 _6490_ (.A1(net1288),
    .A2(_2334_),
    .Y(_2336_),
    .B1(_2335_));
 sg13g2_nand2b_1 _6491_ (.Y(_2337_),
    .B(net1298),
    .A_N(_2336_));
 sg13g2_mux2_1 _6492_ (.A0(\s0.data_out[8][0] ),
    .A1(\s0.data_out[9][0] ),
    .S(net1306),
    .X(_2338_));
 sg13g2_nand2b_1 _6493_ (.Y(_2339_),
    .B(_2338_),
    .A_N(net1298));
 sg13g2_nor2_1 _6494_ (.A(net1694),
    .B(_2333_),
    .Y(_2340_));
 sg13g2_a221oi_1 _6495_ (.B2(_2339_),
    .C1(net1701),
    .B1(_2337_),
    .A1(net1694),
    .Y(_2341_),
    .A2(_2333_));
 sg13g2_nor3_1 _6496_ (.A(_2326_),
    .B(_2340_),
    .C(_2341_),
    .Y(_2342_));
 sg13g2_nand2_1 _6497_ (.Y(_2343_),
    .A(net1295),
    .B(net610));
 sg13g2_o21ai_1 _6498_ (.B1(_2343_),
    .Y(_2344_),
    .A1(net1295),
    .A2(_3504_));
 sg13g2_nor2_1 _6499_ (.A(net1289),
    .B(net1161),
    .Y(_2345_));
 sg13g2_a21o_1 _6500_ (.A2(_2344_),
    .A1(net1289),
    .B1(_2345_),
    .X(_2346_));
 sg13g2_nand2b_1 _6501_ (.Y(_2347_),
    .B(net610),
    .A_N(net1306));
 sg13g2_a21oi_1 _6502_ (.A1(_2228_),
    .A2(_2347_),
    .Y(_2348_),
    .B1(net1299));
 sg13g2_a21oi_1 _6503_ (.A1(net1299),
    .A2(_2346_),
    .Y(_2349_),
    .B1(_2348_));
 sg13g2_a221oi_1 _6504_ (.B2(net1679),
    .C1(_2342_),
    .B1(_2349_),
    .A1(net1688),
    .Y(_2350_),
    .A2(_2325_));
 sg13g2_nand2_1 _6505_ (.Y(_2351_),
    .A(net1296),
    .B(net553));
 sg13g2_mux2_1 _6506_ (.A0(\s0.data_out[9][7] ),
    .A1(\s0.data_out[8][7] ),
    .S(net1296),
    .X(_2352_));
 sg13g2_nor2b_1 _6507_ (.A(net1292),
    .B_N(net1321),
    .Y(_2353_));
 sg13g2_a21o_1 _6508_ (.A2(_2352_),
    .A1(net1292),
    .B1(_2353_),
    .X(_2354_));
 sg13g2_nand2b_1 _6509_ (.Y(_2355_),
    .B(\s0.data_out[8][7] ),
    .A_N(net1308));
 sg13g2_a21oi_1 _6510_ (.A1(_2237_),
    .A2(_2355_),
    .Y(_2356_),
    .B1(net1302));
 sg13g2_a21oi_1 _6511_ (.A1(net1302),
    .A2(_2354_),
    .Y(_2357_),
    .B1(_2356_));
 sg13g2_nand2_1 _6512_ (.Y(_2358_),
    .A(net1296),
    .B(net640));
 sg13g2_mux2_1 _6513_ (.A0(\s0.data_out[9][6] ),
    .A1(\s0.data_out[8][6] ),
    .S(net1296),
    .X(_2359_));
 sg13g2_nor2b_1 _6514_ (.A(net1292),
    .B_N(net1326),
    .Y(_2360_));
 sg13g2_a21o_1 _6515_ (.A2(_2359_),
    .A1(net1292),
    .B1(_2360_),
    .X(_2361_));
 sg13g2_nand2b_1 _6516_ (.Y(_2362_),
    .B(net640),
    .A_N(net1308));
 sg13g2_a21oi_1 _6517_ (.A1(_2244_),
    .A2(_2362_),
    .Y(_2363_),
    .B1(net1302));
 sg13g2_a21oi_1 _6518_ (.A1(net1302),
    .A2(_2361_),
    .Y(_2364_),
    .B1(_2363_));
 sg13g2_a22oi_1 _6519_ (.Y(_2365_),
    .B1(_2364_),
    .B2(net1654),
    .A2(_2357_),
    .A1(net1641));
 sg13g2_or2_1 _6520_ (.X(_2366_),
    .B(_2357_),
    .A(net1645));
 sg13g2_nor2_1 _6521_ (.A(net1654),
    .B(_2364_),
    .Y(_2367_));
 sg13g2_nand3b_1 _6522_ (.B(_2365_),
    .C(_2366_),
    .Y(_2368_),
    .A_N(_2367_));
 sg13g2_nand2_1 _6523_ (.Y(_2369_),
    .A(net1297),
    .B(net813));
 sg13g2_mux2_1 _6524_ (.A0(\s0.data_out[9][5] ),
    .A1(\s0.data_out[8][5] ),
    .S(net1297),
    .X(_2370_));
 sg13g2_nor2b_1 _6525_ (.A(net1290),
    .B_N(net1331),
    .Y(_2371_));
 sg13g2_a21oi_1 _6526_ (.A1(net1293),
    .A2(_2370_),
    .Y(_2372_),
    .B1(_2371_));
 sg13g2_nand2b_1 _6527_ (.Y(_2373_),
    .B(net1302),
    .A_N(_2372_));
 sg13g2_o21ai_1 _6528_ (.B1(_2263_),
    .Y(_2374_),
    .A1(net1308),
    .A2(_3509_));
 sg13g2_nand2b_2 _6529_ (.Y(_2375_),
    .B(_2374_),
    .A_N(net1302));
 sg13g2_nand2_1 _6530_ (.Y(_2376_),
    .A(_2373_),
    .B(_2375_));
 sg13g2_nand3_1 _6531_ (.B(_2373_),
    .C(_2375_),
    .A(net1664),
    .Y(_2377_));
 sg13g2_nor2b_1 _6532_ (.A(net470),
    .B_N(net1336),
    .Y(_2378_));
 sg13g2_nand2_1 _6533_ (.Y(_2379_),
    .A(net1297),
    .B(net773));
 sg13g2_mux2_1 _6534_ (.A0(\s0.data_out[9][4] ),
    .A1(\s0.data_out[8][4] ),
    .S(net1295),
    .X(_2380_));
 sg13g2_a21oi_1 _6535_ (.A1(net1290),
    .A2(_2380_),
    .Y(_2381_),
    .B1(_2378_));
 sg13g2_nand2b_1 _6536_ (.Y(_2382_),
    .B(net1299),
    .A_N(_2381_));
 sg13g2_o21ai_1 _6537_ (.B1(_2255_),
    .Y(_2383_),
    .A1(net1306),
    .A2(_3510_));
 sg13g2_nand2b_1 _6538_ (.Y(_2384_),
    .B(_2383_),
    .A_N(net1299));
 sg13g2_nand3_1 _6539_ (.B(_2382_),
    .C(_2384_),
    .A(net1673),
    .Y(_2385_));
 sg13g2_nand2_1 _6540_ (.Y(_2386_),
    .A(_2377_),
    .B(_2385_));
 sg13g2_a21oi_1 _6541_ (.A1(_2382_),
    .A2(_2384_),
    .Y(_2387_),
    .B1(net1673));
 sg13g2_a21oi_1 _6542_ (.A1(_2373_),
    .A2(_2375_),
    .Y(_2388_),
    .B1(net1664));
 sg13g2_nor2_1 _6543_ (.A(net1679),
    .B(_2349_),
    .Y(_2389_));
 sg13g2_or3_1 _6544_ (.A(_2387_),
    .B(_2388_),
    .C(_2389_),
    .X(_2390_));
 sg13g2_or4_1 _6545_ (.A(_2350_),
    .B(_2368_),
    .C(_2386_),
    .D(_2390_),
    .X(_2391_));
 sg13g2_a21o_1 _6546_ (.A2(_2376_),
    .A1(_3403_),
    .B1(_2385_),
    .X(_2392_));
 sg13g2_a21oi_1 _6547_ (.A1(_2377_),
    .A2(_2392_),
    .Y(_2393_),
    .B1(_2368_));
 sg13g2_nor2b_1 _6548_ (.A(_2365_),
    .B_N(_2366_),
    .Y(_2394_));
 sg13g2_nor3_1 _6549_ (.A(_2312_),
    .B(_2393_),
    .C(_2394_),
    .Y(_2395_));
 sg13g2_or2_1 _6550_ (.X(_2396_),
    .B(net1558),
    .A(net388));
 sg13g2_a21oi_1 _6551_ (.A1(_2391_),
    .A2(_2395_),
    .Y(_0335_),
    .B1(_2396_));
 sg13g2_and2_1 _6552_ (.A(net1289),
    .B(\s0.data_out[8][0] ),
    .X(_2397_));
 sg13g2_o21ai_1 _6553_ (.B1(net1298),
    .Y(_2398_),
    .A1(_2335_),
    .A2(_2397_));
 sg13g2_nand3_1 _6554_ (.B(_2339_),
    .C(_2398_),
    .A(net1726),
    .Y(_2399_));
 sg13g2_o21ai_1 _6555_ (.B1(_2399_),
    .Y(_2400_),
    .A1(net1726),
    .A2(net607));
 sg13g2_inv_1 _6556_ (.Y(_0336_),
    .A(_2400_));
 sg13g2_nor2_1 _6557_ (.A(_3394_),
    .B(_3513_),
    .Y(_2401_));
 sg13g2_o21ai_1 _6558_ (.B1(net1298),
    .Y(_2402_),
    .A1(_2329_),
    .A2(_2401_));
 sg13g2_nor2_1 _6559_ (.A(net1596),
    .B(_2332_),
    .Y(_2403_));
 sg13g2_a22oi_1 _6560_ (.Y(_0337_),
    .B1(_2402_),
    .B2(_2403_),
    .A2(_3506_),
    .A1(net1596));
 sg13g2_nor2_1 _6561_ (.A(_3394_),
    .B(_3512_),
    .Y(_2404_));
 sg13g2_o21ai_1 _6562_ (.B1(net1298),
    .Y(_2405_),
    .A1(_2321_),
    .A2(_2404_));
 sg13g2_nor2_1 _6563_ (.A(net1596),
    .B(_2324_),
    .Y(_2406_));
 sg13g2_a22oi_1 _6564_ (.Y(_0338_),
    .B1(_2405_),
    .B2(_2406_),
    .A2(_3505_),
    .A1(net1596));
 sg13g2_nor2_1 _6565_ (.A(_3394_),
    .B(_3511_),
    .Y(_2407_));
 sg13g2_o21ai_1 _6566_ (.B1(net1299),
    .Y(_2408_),
    .A1(_2345_),
    .A2(_2407_));
 sg13g2_nor2_1 _6567_ (.A(net1596),
    .B(_2348_),
    .Y(_2409_));
 sg13g2_a22oi_1 _6568_ (.Y(_0339_),
    .B1(_2408_),
    .B2(_2409_),
    .A2(_3504_),
    .A1(net1596));
 sg13g2_nor2_1 _6569_ (.A(_3394_),
    .B(_3510_),
    .Y(_2410_));
 sg13g2_o21ai_1 _6570_ (.B1(net1299),
    .Y(_2411_),
    .A1(_2378_),
    .A2(_2410_));
 sg13g2_nand3_1 _6571_ (.B(_2384_),
    .C(_2411_),
    .A(net1719),
    .Y(_2412_));
 sg13g2_o21ai_1 _6572_ (.B1(_2412_),
    .Y(_2413_),
    .A1(net1719),
    .A2(net672));
 sg13g2_inv_1 _6573_ (.Y(_0340_),
    .A(_2413_));
 sg13g2_nor2_1 _6574_ (.A(_3394_),
    .B(_3509_),
    .Y(_2414_));
 sg13g2_o21ai_1 _6575_ (.B1(net1302),
    .Y(_2415_),
    .A1(_2371_),
    .A2(_2414_));
 sg13g2_nand3_1 _6576_ (.B(_2375_),
    .C(_2415_),
    .A(net1719),
    .Y(_2416_));
 sg13g2_o21ai_1 _6577_ (.B1(_2416_),
    .Y(_2417_),
    .A1(net1719),
    .A2(net633));
 sg13g2_inv_1 _6578_ (.Y(_0341_),
    .A(_2417_));
 sg13g2_nor2_1 _6579_ (.A(_3394_),
    .B(_3508_),
    .Y(_2418_));
 sg13g2_o21ai_1 _6580_ (.B1(net1305),
    .Y(_2419_),
    .A1(_2360_),
    .A2(_2418_));
 sg13g2_nand3b_1 _6581_ (.B(_2419_),
    .C(net1719),
    .Y(_2420_),
    .A_N(_2363_));
 sg13g2_o21ai_1 _6582_ (.B1(_2420_),
    .Y(_2421_),
    .A1(net1727),
    .A2(net735));
 sg13g2_inv_1 _6583_ (.Y(_0342_),
    .A(_2421_));
 sg13g2_nor2_1 _6584_ (.A(_3394_),
    .B(_3507_),
    .Y(_2422_));
 sg13g2_o21ai_1 _6585_ (.B1(net1302),
    .Y(_2423_),
    .A1(_2353_),
    .A2(_2422_));
 sg13g2_nor2_1 _6586_ (.A(net1603),
    .B(_2356_),
    .Y(_2424_));
 sg13g2_a22oi_1 _6587_ (.Y(_0343_),
    .B1(_2423_),
    .B2(_2424_),
    .A2(_3503_),
    .A1(net1598));
 sg13g2_o21ai_1 _6588_ (.B1(net1291),
    .Y(_2425_),
    .A1(net1629),
    .A2(net1281));
 sg13g2_nor2b_1 _6589_ (.A(net1629),
    .B_N(net1284),
    .Y(_2426_));
 sg13g2_or2_1 _6590_ (.X(_2427_),
    .B(_2426_),
    .A(_2425_));
 sg13g2_o21ai_1 _6591_ (.B1(_2427_),
    .Y(_2428_),
    .A1(net1291),
    .A2(_2309_));
 sg13g2_nor2_1 _6592_ (.A(net459),
    .B(net1285),
    .Y(_2429_));
 sg13g2_nor2_1 _6593_ (.A(_2427_),
    .B(_2429_),
    .Y(_2430_));
 sg13g2_o21ai_1 _6594_ (.B1(_3394_),
    .Y(_2431_),
    .A1(net459),
    .A2(net1296));
 sg13g2_o21ai_1 _6595_ (.B1(_2431_),
    .Y(_2432_),
    .A1(net1281),
    .A2(_2425_));
 sg13g2_nor2_1 _6596_ (.A(_2430_),
    .B(_2432_),
    .Y(_2433_));
 sg13g2_o21ai_1 _6597_ (.B1(net1719),
    .Y(_2434_),
    .A1(net689),
    .A2(_2428_));
 sg13g2_nor2_1 _6598_ (.A(_2433_),
    .B(_2434_),
    .Y(_0000_));
 sg13g2_nor2_1 _6599_ (.A(net1590),
    .B(_2428_),
    .Y(_0001_));
 sg13g2_and2_1 _6600_ (.A(net1720),
    .B(net393),
    .X(_0002_));
 sg13g2_nand2_1 _6601_ (.Y(_2435_),
    .A(net1283),
    .B(net590));
 sg13g2_mux2_1 _6602_ (.A0(\s0.data_out[8][2] ),
    .A1(\s0.data_out[7][2] ),
    .S(net1286),
    .X(_2436_));
 sg13g2_nor2b_1 _6603_ (.A(net1276),
    .B_N(net1341),
    .Y(_2437_));
 sg13g2_a21o_1 _6604_ (.A2(_2436_),
    .A1(net1276),
    .B1(_2437_),
    .X(_2438_));
 sg13g2_nand2b_1 _6605_ (.Y(_2439_),
    .B(\s0.data_out[7][2] ),
    .A_N(net1294));
 sg13g2_a21oi_1 _6606_ (.A1(_2319_),
    .A2(_2439_),
    .Y(_2440_),
    .B1(net1287));
 sg13g2_a21oi_1 _6607_ (.A1(net1287),
    .A2(_2438_),
    .Y(_2441_),
    .B1(_2440_));
 sg13g2_nor2_1 _6608_ (.A(net1688),
    .B(_2441_),
    .Y(_2442_));
 sg13g2_nand2_1 _6609_ (.Y(_2443_),
    .A(net1283),
    .B(net796));
 sg13g2_mux2_1 _6610_ (.A0(\s0.data_out[8][1] ),
    .A1(\s0.data_out[7][1] ),
    .S(net1283),
    .X(_2444_));
 sg13g2_nor2b_1 _6611_ (.A(net1276),
    .B_N(net1347),
    .Y(_2445_));
 sg13g2_a21o_1 _6612_ (.A2(_2444_),
    .A1(net1276),
    .B1(_2445_),
    .X(_2446_));
 sg13g2_nand2b_1 _6613_ (.Y(_2447_),
    .B(\s0.data_out[7][1] ),
    .A_N(net1294));
 sg13g2_a21oi_1 _6614_ (.A1(_2327_),
    .A2(_2447_),
    .Y(_2448_),
    .B1(net1287));
 sg13g2_a21oi_1 _6615_ (.A1(net1287),
    .A2(_2446_),
    .Y(_2449_),
    .B1(_2448_));
 sg13g2_mux2_1 _6616_ (.A0(\s0.data_out[8][0] ),
    .A1(\s0.data_out[7][0] ),
    .S(net1286),
    .X(_2450_));
 sg13g2_nor2b_1 _6617_ (.A(net1277),
    .B_N(net1351),
    .Y(_2451_));
 sg13g2_a21oi_1 _6618_ (.A1(net1276),
    .A2(_2450_),
    .Y(_2452_),
    .B1(_2451_));
 sg13g2_nand2b_1 _6619_ (.Y(_2453_),
    .B(net1287),
    .A_N(_2452_));
 sg13g2_mux2_1 _6620_ (.A0(\s0.data_out[7][0] ),
    .A1(\s0.data_out[8][0] ),
    .S(net1294),
    .X(_2454_));
 sg13g2_nand2b_1 _6621_ (.Y(_2455_),
    .B(_2454_),
    .A_N(net1287));
 sg13g2_nor2_1 _6622_ (.A(net1699),
    .B(_2449_),
    .Y(_2456_));
 sg13g2_a221oi_1 _6623_ (.B2(_2455_),
    .C1(net1701),
    .B1(_2453_),
    .A1(net1699),
    .Y(_2457_),
    .A2(_2449_));
 sg13g2_nor3_1 _6624_ (.A(_2442_),
    .B(_2456_),
    .C(_2457_),
    .Y(_2458_));
 sg13g2_nand2_1 _6625_ (.Y(_2459_),
    .A(net1283),
    .B(net576));
 sg13g2_mux2_1 _6626_ (.A0(\s0.data_out[8][3] ),
    .A1(\s0.data_out[7][3] ),
    .S(net1283),
    .X(_2460_));
 sg13g2_nor2b_1 _6627_ (.A(net1277),
    .B_N(net1339),
    .Y(_2461_));
 sg13g2_a21o_1 _6628_ (.A2(_2460_),
    .A1(net1277),
    .B1(_2461_),
    .X(_2462_));
 sg13g2_nand2b_1 _6629_ (.Y(_2463_),
    .B(net576),
    .A_N(net1295));
 sg13g2_a21oi_1 _6630_ (.A1(_2343_),
    .A2(_2463_),
    .Y(_2464_),
    .B1(net1289));
 sg13g2_a21oi_1 _6631_ (.A1(net1289),
    .A2(_2462_),
    .Y(_2465_),
    .B1(_2464_));
 sg13g2_a221oi_1 _6632_ (.B2(net1679),
    .C1(_2458_),
    .B1(_2465_),
    .A1(net1688),
    .Y(_2466_),
    .A2(_2441_));
 sg13g2_nand2_1 _6633_ (.Y(_2467_),
    .A(net1284),
    .B(\s0.data_out[7][6] ));
 sg13g2_mux2_1 _6634_ (.A0(\s0.data_out[8][6] ),
    .A1(\s0.data_out[7][6] ),
    .S(net1285),
    .X(_2468_));
 sg13g2_nor2b_1 _6635_ (.A(net1281),
    .B_N(net1326),
    .Y(_2469_));
 sg13g2_a21o_1 _6636_ (.A2(_2468_),
    .A1(net1280),
    .B1(_2469_),
    .X(_2470_));
 sg13g2_nand2b_1 _6637_ (.Y(_2471_),
    .B(\s0.data_out[7][6] ),
    .A_N(net1296));
 sg13g2_a21oi_1 _6638_ (.A1(_2358_),
    .A2(_2471_),
    .Y(_2472_),
    .B1(net1291));
 sg13g2_a21oi_1 _6639_ (.A1(net1291),
    .A2(_2470_),
    .Y(_2473_),
    .B1(_2472_));
 sg13g2_nand2_1 _6640_ (.Y(_2474_),
    .A(net1284),
    .B(net460));
 sg13g2_mux2_1 _6641_ (.A0(\s0.data_out[8][7] ),
    .A1(\s0.data_out[7][7] ),
    .S(net1285),
    .X(_2475_));
 sg13g2_nor2b_1 _6642_ (.A(net1280),
    .B_N(net1321),
    .Y(_2476_));
 sg13g2_a21o_1 _6643_ (.A2(_2475_),
    .A1(net1280),
    .B1(_2476_),
    .X(_2477_));
 sg13g2_nand2b_1 _6644_ (.Y(_2478_),
    .B(net460),
    .A_N(net1296));
 sg13g2_a21oi_1 _6645_ (.A1(_2351_),
    .A2(_2478_),
    .Y(_2479_),
    .B1(net1291));
 sg13g2_a21oi_1 _6646_ (.A1(net1291),
    .A2(_2477_),
    .Y(_2480_),
    .B1(_2479_));
 sg13g2_a22oi_1 _6647_ (.Y(_2481_),
    .B1(_2480_),
    .B2(net1639),
    .A2(_2473_),
    .A1(net1649));
 sg13g2_or2_1 _6648_ (.X(_2482_),
    .B(_2473_),
    .A(net1649));
 sg13g2_or2_1 _6649_ (.X(_2483_),
    .B(_2480_),
    .A(net1639));
 sg13g2_nand3_1 _6650_ (.B(_2482_),
    .C(_2483_),
    .A(_2481_),
    .Y(_2484_));
 sg13g2_mux2_1 _6651_ (.A0(\s0.data_out[8][4] ),
    .A1(\s0.data_out[7][4] ),
    .S(net1285),
    .X(_2485_));
 sg13g2_nor2b_1 _6652_ (.A(net1280),
    .B_N(net1336),
    .Y(_2486_));
 sg13g2_a21o_1 _6653_ (.A2(_2485_),
    .A1(net1280),
    .B1(_2486_),
    .X(_2487_));
 sg13g2_nand2b_1 _6654_ (.Y(_2488_),
    .B(net740),
    .A_N(net1297));
 sg13g2_a21oi_1 _6655_ (.A1(_2379_),
    .A2(_2488_),
    .Y(_2489_),
    .B1(net1290));
 sg13g2_a21oi_1 _6656_ (.A1(net1290),
    .A2(_2487_),
    .Y(_2490_),
    .B1(_2489_));
 sg13g2_mux2_1 _6657_ (.A0(\s0.data_out[8][5] ),
    .A1(\s0.data_out[7][5] ),
    .S(net1285),
    .X(_2491_));
 sg13g2_nor2b_1 _6658_ (.A(net1280),
    .B_N(net1331),
    .Y(_2492_));
 sg13g2_a21o_1 _6659_ (.A2(_2491_),
    .A1(net1280),
    .B1(_2492_),
    .X(_2493_));
 sg13g2_nand2b_1 _6660_ (.Y(_2494_),
    .B(net758),
    .A_N(net1297));
 sg13g2_a21oi_1 _6661_ (.A1(_2369_),
    .A2(_2494_),
    .Y(_2495_),
    .B1(net1290));
 sg13g2_a21oi_1 _6662_ (.A1(net1290),
    .A2(_2493_),
    .Y(_2496_),
    .B1(_2495_));
 sg13g2_a22oi_1 _6663_ (.Y(_2497_),
    .B1(_2496_),
    .B2(net1657),
    .A2(_2490_),
    .A1(net1668));
 sg13g2_nor2_1 _6664_ (.A(net1668),
    .B(_2490_),
    .Y(_2498_));
 sg13g2_nor2_1 _6665_ (.A(net1659),
    .B(_2496_),
    .Y(_2499_));
 sg13g2_nor2_1 _6666_ (.A(net1679),
    .B(_2465_),
    .Y(_2500_));
 sg13g2_nor3_1 _6667_ (.A(_2498_),
    .B(_2499_),
    .C(_2500_),
    .Y(_2501_));
 sg13g2_nand2_1 _6668_ (.Y(_2502_),
    .A(_2497_),
    .B(_2501_));
 sg13g2_or3_1 _6669_ (.A(_2466_),
    .B(_2484_),
    .C(_2502_),
    .X(_2503_));
 sg13g2_nor3_1 _6670_ (.A(_2484_),
    .B(_2497_),
    .C(_2499_),
    .Y(_2504_));
 sg13g2_nor2b_1 _6671_ (.A(_2481_),
    .B_N(_2483_),
    .Y(_2505_));
 sg13g2_nor3_1 _6672_ (.A(_2428_),
    .B(_2504_),
    .C(_2505_),
    .Y(_2506_));
 sg13g2_or2_1 _6673_ (.X(_2507_),
    .B(net1556),
    .A(net391));
 sg13g2_a21oi_1 _6674_ (.A1(_2503_),
    .A2(_2506_),
    .Y(_0003_),
    .B1(_2507_));
 sg13g2_and2_1 _6675_ (.A(net1277),
    .B(\s0.data_out[7][0] ),
    .X(_2508_));
 sg13g2_o21ai_1 _6676_ (.B1(net1287),
    .Y(_2509_),
    .A1(_2451_),
    .A2(_2508_));
 sg13g2_nand3_1 _6677_ (.B(_2455_),
    .C(_2509_),
    .A(net1719),
    .Y(_2510_));
 sg13g2_o21ai_1 _6678_ (.B1(_2510_),
    .Y(_2511_),
    .A1(net1717),
    .A2(net742));
 sg13g2_inv_1 _6679_ (.Y(_0004_),
    .A(_2511_));
 sg13g2_nor2_1 _6680_ (.A(net1170),
    .B(_3514_),
    .Y(_2512_));
 sg13g2_o21ai_1 _6681_ (.B1(net1287),
    .Y(_2513_),
    .A1(_2445_),
    .A2(_2512_));
 sg13g2_nor2_1 _6682_ (.A(net1587),
    .B(_2448_),
    .Y(_2514_));
 sg13g2_a22oi_1 _6683_ (.Y(_0005_),
    .B1(_2513_),
    .B2(_2514_),
    .A2(_3513_),
    .A1(net1588));
 sg13g2_nor2_1 _6684_ (.A(net1170),
    .B(_3516_),
    .Y(_2515_));
 sg13g2_o21ai_1 _6685_ (.B1(net1288),
    .Y(_2516_),
    .A1(_2437_),
    .A2(_2515_));
 sg13g2_nor2_1 _6686_ (.A(net1588),
    .B(_2440_),
    .Y(_2517_));
 sg13g2_a22oi_1 _6687_ (.Y(_0006_),
    .B1(_2516_),
    .B2(_2517_),
    .A2(_3512_),
    .A1(net1588));
 sg13g2_nor2_1 _6688_ (.A(net1170),
    .B(_3515_),
    .Y(_2518_));
 sg13g2_o21ai_1 _6689_ (.B1(net1289),
    .Y(_2519_),
    .A1(_2461_),
    .A2(_2518_));
 sg13g2_nor2_1 _6690_ (.A(net1587),
    .B(_2464_),
    .Y(_2520_));
 sg13g2_a22oi_1 _6691_ (.Y(_0007_),
    .B1(_2519_),
    .B2(_2520_),
    .A2(_3511_),
    .A1(net1588));
 sg13g2_nor2_1 _6692_ (.A(net1169),
    .B(_3518_),
    .Y(_2521_));
 sg13g2_o21ai_1 _6693_ (.B1(net1290),
    .Y(_2522_),
    .A1(_2486_),
    .A2(_2521_));
 sg13g2_nor2_1 _6694_ (.A(net1589),
    .B(_2489_),
    .Y(_2523_));
 sg13g2_a22oi_1 _6695_ (.Y(_0008_),
    .B1(_2522_),
    .B2(_2523_),
    .A2(_3510_),
    .A1(net1589));
 sg13g2_and2_1 _6696_ (.A(net1280),
    .B(net758),
    .X(_2524_));
 sg13g2_o21ai_1 _6697_ (.B1(net1290),
    .Y(_2525_),
    .A1(_2492_),
    .A2(_2524_));
 sg13g2_nor2_1 _6698_ (.A(net1589),
    .B(_2495_),
    .Y(_2526_));
 sg13g2_a22oi_1 _6699_ (.Y(_0009_),
    .B1(_2525_),
    .B2(_2526_),
    .A2(_3509_),
    .A1(net1589));
 sg13g2_and2_1 _6700_ (.A(net1281),
    .B(\s0.data_out[7][6] ),
    .X(_2527_));
 sg13g2_o21ai_1 _6701_ (.B1(net1291),
    .Y(_2528_),
    .A1(_2469_),
    .A2(_2527_));
 sg13g2_nor2_1 _6702_ (.A(net1589),
    .B(_2472_),
    .Y(_2529_));
 sg13g2_a22oi_1 _6703_ (.Y(_0010_),
    .B1(_2528_),
    .B2(_2529_),
    .A2(_3508_),
    .A1(net1589));
 sg13g2_nor2_1 _6704_ (.A(net1169),
    .B(_3517_),
    .Y(_2530_));
 sg13g2_o21ai_1 _6705_ (.B1(net1291),
    .Y(_2531_),
    .A1(_2476_),
    .A2(_2530_));
 sg13g2_nor2_1 _6706_ (.A(net1589),
    .B(_2479_),
    .Y(_2532_));
 sg13g2_a22oi_1 _6707_ (.Y(_0011_),
    .B1(_2531_),
    .B2(_2532_),
    .A2(_3507_),
    .A1(net1589));
 sg13g2_o21ai_1 _6708_ (.B1(net1282),
    .Y(_2533_),
    .A1(net1634),
    .A2(net1270));
 sg13g2_nand2_1 _6709_ (.Y(_2534_),
    .A(net1622),
    .B(net1275));
 sg13g2_nand2b_1 _6710_ (.Y(_2535_),
    .B(_2534_),
    .A_N(_2533_));
 sg13g2_o21ai_1 _6711_ (.B1(_2535_),
    .Y(_2536_),
    .A1(net1279),
    .A2(_2426_));
 sg13g2_nor2_1 _6712_ (.A(net459),
    .B(_2536_),
    .Y(_2537_));
 sg13g2_nor2_1 _6713_ (.A(net422),
    .B(net1275),
    .Y(_2538_));
 sg13g2_nor2_1 _6714_ (.A(net1270),
    .B(_2533_),
    .Y(_2539_));
 sg13g2_o21ai_1 _6715_ (.B1(net1169),
    .Y(_2540_),
    .A1(net422),
    .A2(net1284));
 sg13g2_o21ai_1 _6716_ (.B1(_2540_),
    .Y(_2541_),
    .A1(_2535_),
    .A2(_2538_));
 sg13g2_o21ai_1 _6717_ (.B1(net1719),
    .Y(_2542_),
    .A1(_2539_),
    .A2(_2541_));
 sg13g2_nor2_1 _6718_ (.A(_2537_),
    .B(_2542_),
    .Y(_0012_));
 sg13g2_nor2_1 _6719_ (.A(net1590),
    .B(_2536_),
    .Y(_0013_));
 sg13g2_and2_1 _6720_ (.A(net1718),
    .B(net397),
    .X(_0014_));
 sg13g2_nand2_1 _6721_ (.Y(_2543_),
    .A(net1272),
    .B(net549));
 sg13g2_mux2_1 _6722_ (.A0(\s0.data_out[7][2] ),
    .A1(\s0.data_out[6][2] ),
    .S(net1272),
    .X(_2544_));
 sg13g2_nor2b_1 _6723_ (.A(net1265),
    .B_N(net1341),
    .Y(_2545_));
 sg13g2_a21o_1 _6724_ (.A2(_2544_),
    .A1(net1266),
    .B1(_2545_),
    .X(_2546_));
 sg13g2_nand2b_1 _6725_ (.Y(_2547_),
    .B(net549),
    .A_N(net1283));
 sg13g2_a21oi_1 _6726_ (.A1(_2435_),
    .A2(_2547_),
    .Y(_2548_),
    .B1(net1276));
 sg13g2_a21oi_1 _6727_ (.A1(net1278),
    .A2(_2546_),
    .Y(_2549_),
    .B1(_2548_));
 sg13g2_or2_1 _6728_ (.X(_2550_),
    .B(_2549_),
    .A(net1685));
 sg13g2_nand2_1 _6729_ (.Y(_2551_),
    .A(net1272),
    .B(net737));
 sg13g2_o21ai_1 _6730_ (.B1(_2551_),
    .Y(_2552_),
    .A1(net1272),
    .A2(_3514_));
 sg13g2_nor2b_1 _6731_ (.A(net1265),
    .B_N(net1345),
    .Y(_2553_));
 sg13g2_a21o_1 _6732_ (.A2(_2552_),
    .A1(net1266),
    .B1(_2553_),
    .X(_2554_));
 sg13g2_nand2b_1 _6733_ (.Y(_2555_),
    .B(net737),
    .A_N(net1286));
 sg13g2_a21oi_1 _6734_ (.A1(_2443_),
    .A2(_2555_),
    .Y(_2556_),
    .B1(net1276));
 sg13g2_a21oi_1 _6735_ (.A1(net1276),
    .A2(_2554_),
    .Y(_2557_),
    .B1(_2556_));
 sg13g2_mux2_1 _6736_ (.A0(\s0.data_out[7][0] ),
    .A1(\s0.data_out[6][0] ),
    .S(net1272),
    .X(_2558_));
 sg13g2_nor2b_1 _6737_ (.A(net1265),
    .B_N(net1349),
    .Y(_2559_));
 sg13g2_a21oi_1 _6738_ (.A1(net1266),
    .A2(_2558_),
    .Y(_2560_),
    .B1(_2559_));
 sg13g2_nand2b_1 _6739_ (.Y(_2561_),
    .B(net1278),
    .A_N(_2560_));
 sg13g2_mux2_1 _6740_ (.A0(\s0.data_out[6][0] ),
    .A1(\s0.data_out[7][0] ),
    .S(net1283),
    .X(_2562_));
 sg13g2_nand2_1 _6741_ (.Y(_2563_),
    .A(net1170),
    .B(_2562_));
 sg13g2_a221oi_1 _6742_ (.B2(_2563_),
    .C1(net1700),
    .B1(_2561_),
    .A1(net1692),
    .Y(_2564_),
    .A2(_2557_));
 sg13g2_o21ai_1 _6743_ (.B1(_2550_),
    .Y(_2565_),
    .A1(net1693),
    .A2(_2557_));
 sg13g2_nand2_1 _6744_ (.Y(_2566_),
    .A(net1273),
    .B(\s0.data_out[6][3] ));
 sg13g2_mux2_1 _6745_ (.A0(\s0.data_out[7][3] ),
    .A1(\s0.data_out[6][3] ),
    .S(net1273),
    .X(_2567_));
 sg13g2_nor2b_1 _6746_ (.A(net1267),
    .B_N(net1339),
    .Y(_2568_));
 sg13g2_a21o_1 _6747_ (.A2(_2567_),
    .A1(net1267),
    .B1(_2568_),
    .X(_2569_));
 sg13g2_nand2b_1 _6748_ (.Y(_2570_),
    .B(\s0.data_out[6][3] ),
    .A_N(net1283));
 sg13g2_a21oi_1 _6749_ (.A1(_2459_),
    .A2(_2570_),
    .Y(_2571_),
    .B1(net1278));
 sg13g2_a21oi_1 _6750_ (.A1(net1278),
    .A2(_2569_),
    .Y(_2572_),
    .B1(_2571_));
 sg13g2_a22oi_1 _6751_ (.Y(_2573_),
    .B1(_2572_),
    .B2(net1677),
    .A2(_2549_),
    .A1(net1689));
 sg13g2_o21ai_1 _6752_ (.B1(_2573_),
    .Y(_2574_),
    .A1(_2564_),
    .A2(_2565_));
 sg13g2_nand2_1 _6753_ (.Y(_2575_),
    .A(net1274),
    .B(net668));
 sg13g2_mux2_1 _6754_ (.A0(\s0.data_out[7][7] ),
    .A1(\s0.data_out[6][7] ),
    .S(net1275),
    .X(_2576_));
 sg13g2_nor2b_1 _6755_ (.A(net1270),
    .B_N(net1324),
    .Y(_2577_));
 sg13g2_a21o_1 _6756_ (.A2(_2576_),
    .A1(net1270),
    .B1(_2577_),
    .X(_2578_));
 sg13g2_nand2b_1 _6757_ (.Y(_2579_),
    .B(\s0.data_out[6][7] ),
    .A_N(net1284));
 sg13g2_a21oi_1 _6758_ (.A1(_2474_),
    .A2(_2579_),
    .Y(_2580_),
    .B1(net1279));
 sg13g2_a21oi_1 _6759_ (.A1(net1279),
    .A2(_2578_),
    .Y(_2581_),
    .B1(_2580_));
 sg13g2_nand2_1 _6760_ (.Y(_2582_),
    .A(net1274),
    .B(net779));
 sg13g2_mux2_1 _6761_ (.A0(\s0.data_out[7][6] ),
    .A1(\s0.data_out[6][6] ),
    .S(net1274),
    .X(_2583_));
 sg13g2_nor2b_1 _6762_ (.A(net1269),
    .B_N(net1326),
    .Y(_2584_));
 sg13g2_a21o_1 _6763_ (.A2(_2583_),
    .A1(net1270),
    .B1(_2584_),
    .X(_2585_));
 sg13g2_nand2b_1 _6764_ (.Y(_2586_),
    .B(\s0.data_out[6][6] ),
    .A_N(net1284));
 sg13g2_a21oi_1 _6765_ (.A1(_2467_),
    .A2(_2586_),
    .Y(_2587_),
    .B1(net1279));
 sg13g2_a21oi_1 _6766_ (.A1(net1279),
    .A2(_2585_),
    .Y(_2588_),
    .B1(_2587_));
 sg13g2_a22oi_1 _6767_ (.Y(_2589_),
    .B1(_2588_),
    .B2(net1648),
    .A2(_2581_),
    .A1(net1639));
 sg13g2_or2_1 _6768_ (.X(_2590_),
    .B(_2581_),
    .A(net1639));
 sg13g2_or2_1 _6769_ (.X(_2591_),
    .B(_2588_),
    .A(net1648));
 sg13g2_and3_1 _6770_ (.X(_2592_),
    .A(_2589_),
    .B(_2590_),
    .C(_2591_));
 sg13g2_nor2b_1 _6771_ (.A(net1270),
    .B_N(\s0.data_new_delayed[4] ),
    .Y(_2593_));
 sg13g2_nand2_1 _6772_ (.Y(_2594_),
    .A(net1275),
    .B(\s0.data_out[6][4] ));
 sg13g2_o21ai_1 _6773_ (.B1(_2594_),
    .Y(_2595_),
    .A1(net1275),
    .A2(_3518_));
 sg13g2_a21oi_1 _6774_ (.A1(net1270),
    .A2(_2595_),
    .Y(_2596_),
    .B1(_2593_));
 sg13g2_mux2_1 _6775_ (.A0(\s0.data_out[6][4] ),
    .A1(\s0.data_out[7][4] ),
    .S(net1284),
    .X(_2597_));
 sg13g2_nand2_1 _6776_ (.Y(_2598_),
    .A(net1169),
    .B(_2597_));
 sg13g2_o21ai_1 _6777_ (.B1(_2598_),
    .Y(_2599_),
    .A1(net1169),
    .A2(_2596_));
 sg13g2_or2_1 _6778_ (.X(_2600_),
    .B(_2599_),
    .A(_3406_));
 sg13g2_nand2_1 _6779_ (.Y(_2601_),
    .A(net1274),
    .B(\s0.data_out[6][5] ));
 sg13g2_mux2_1 _6780_ (.A0(\s0.data_out[7][5] ),
    .A1(\s0.data_out[6][5] ),
    .S(net1275),
    .X(_2602_));
 sg13g2_nor2b_1 _6781_ (.A(net1271),
    .B_N(net1334),
    .Y(_2603_));
 sg13g2_a21oi_1 _6782_ (.A1(net1271),
    .A2(_2602_),
    .Y(_2604_),
    .B1(_2603_));
 sg13g2_nand2b_1 _6783_ (.Y(_2605_),
    .B(net1279),
    .A_N(_2604_));
 sg13g2_mux2_1 _6784_ (.A0(\s0.data_out[6][5] ),
    .A1(\s0.data_out[7][5] ),
    .S(net1284),
    .X(_2606_));
 sg13g2_nand2_1 _6785_ (.Y(_2607_),
    .A(_3395_),
    .B(_2606_));
 sg13g2_nand3_1 _6786_ (.B(_2605_),
    .C(_2607_),
    .A(net1657),
    .Y(_2608_));
 sg13g2_nor2_1 _6787_ (.A(net1677),
    .B(_2572_),
    .Y(_2609_));
 sg13g2_a21oi_1 _6788_ (.A1(_2605_),
    .A2(_2607_),
    .Y(_2610_),
    .B1(net1657));
 sg13g2_nor2_1 _6789_ (.A(_2609_),
    .B(_2610_),
    .Y(_2611_));
 sg13g2_xnor2_1 _6790_ (.Y(_2612_),
    .A(net1668),
    .B(_2599_));
 sg13g2_and4_1 _6791_ (.A(_2592_),
    .B(_2608_),
    .C(_2611_),
    .D(_2612_),
    .X(_2613_));
 sg13g2_o21ai_1 _6792_ (.B1(_2608_),
    .Y(_2614_),
    .A1(_2600_),
    .A2(_2610_));
 sg13g2_nand2b_1 _6793_ (.Y(_2615_),
    .B(_2590_),
    .A_N(_2589_));
 sg13g2_a221oi_1 _6794_ (.B2(_2592_),
    .C1(_2536_),
    .B1(_2614_),
    .A1(_2574_),
    .Y(_2616_),
    .A2(_2613_));
 sg13g2_or2_1 _6795_ (.X(_2617_),
    .B(net1556),
    .A(net393));
 sg13g2_a21oi_1 _6796_ (.A1(_2615_),
    .A2(_2616_),
    .Y(_0015_),
    .B1(_2617_));
 sg13g2_a21oi_1 _6797_ (.A1(net1266),
    .A2(\s0.data_out[6][0] ),
    .Y(_2618_),
    .B1(_2559_));
 sg13g2_a21oi_1 _6798_ (.A1(net1170),
    .A2(_2562_),
    .Y(_2619_),
    .B1(net1587));
 sg13g2_o21ai_1 _6799_ (.B1(_2619_),
    .Y(_2620_),
    .A1(net1170),
    .A2(_2618_));
 sg13g2_o21ai_1 _6800_ (.B1(_2620_),
    .Y(_2621_),
    .A1(net1717),
    .A2(net629));
 sg13g2_inv_1 _6801_ (.Y(_0016_),
    .A(net630));
 sg13g2_nor2_1 _6802_ (.A(net1168),
    .B(_3523_),
    .Y(_2622_));
 sg13g2_o21ai_1 _6803_ (.B1(net1278),
    .Y(_2623_),
    .A1(_2553_),
    .A2(_2622_));
 sg13g2_nor2_1 _6804_ (.A(net1587),
    .B(_2556_),
    .Y(_2624_));
 sg13g2_a22oi_1 _6805_ (.Y(_0017_),
    .B1(_2623_),
    .B2(_2624_),
    .A2(_3514_),
    .A1(net1582));
 sg13g2_nor2_1 _6806_ (.A(net1168),
    .B(_3522_),
    .Y(_2625_));
 sg13g2_o21ai_1 _6807_ (.B1(net1278),
    .Y(_2626_),
    .A1(_2545_),
    .A2(_2625_));
 sg13g2_nor2_1 _6808_ (.A(net1587),
    .B(_2548_),
    .Y(_2627_));
 sg13g2_a22oi_1 _6809_ (.Y(_0018_),
    .B1(_2626_),
    .B2(_2627_),
    .A2(_3516_),
    .A1(net1587));
 sg13g2_nor2_1 _6810_ (.A(net1168),
    .B(_3521_),
    .Y(_2628_));
 sg13g2_o21ai_1 _6811_ (.B1(net1278),
    .Y(_2629_),
    .A1(_2568_),
    .A2(_2628_));
 sg13g2_nor2_1 _6812_ (.A(net1587),
    .B(_2571_),
    .Y(_2630_));
 sg13g2_a22oi_1 _6813_ (.Y(_0019_),
    .B1(_2629_),
    .B2(_2630_),
    .A2(_3515_),
    .A1(net1587));
 sg13g2_a21oi_1 _6814_ (.A1(net1270),
    .A2(net654),
    .Y(_2631_),
    .B1(_2593_));
 sg13g2_a21oi_1 _6815_ (.A1(net1169),
    .A2(_2597_),
    .Y(_2632_),
    .B1(net1590));
 sg13g2_o21ai_1 _6816_ (.B1(_2632_),
    .Y(_2633_),
    .A1(net1169),
    .A2(_2631_));
 sg13g2_o21ai_1 _6817_ (.B1(_2633_),
    .Y(_2634_),
    .A1(net1720),
    .A2(net740));
 sg13g2_inv_1 _6818_ (.Y(_0020_),
    .A(net741));
 sg13g2_a21oi_1 _6819_ (.A1(net1271),
    .A2(\s0.data_out[6][5] ),
    .Y(_2635_),
    .B1(_2603_));
 sg13g2_a21oi_1 _6820_ (.A1(net1170),
    .A2(_2606_),
    .Y(_2636_),
    .B1(net1590));
 sg13g2_o21ai_1 _6821_ (.B1(_2636_),
    .Y(_2637_),
    .A1(net1169),
    .A2(_2635_));
 sg13g2_o21ai_1 _6822_ (.B1(_2637_),
    .Y(_2638_),
    .A1(net1718),
    .A2(net758));
 sg13g2_inv_1 _6823_ (.Y(_0021_),
    .A(net759));
 sg13g2_nor2_1 _6824_ (.A(net1167),
    .B(_3520_),
    .Y(_2639_));
 sg13g2_o21ai_1 _6825_ (.B1(net1279),
    .Y(_2640_),
    .A1(_2584_),
    .A2(_2639_));
 sg13g2_nand3b_1 _6826_ (.B(_2640_),
    .C(net1718),
    .Y(_2641_),
    .A_N(_2587_));
 sg13g2_o21ai_1 _6827_ (.B1(_2641_),
    .Y(_2642_),
    .A1(net1718),
    .A2(net810));
 sg13g2_inv_1 _6828_ (.Y(_0022_),
    .A(net811));
 sg13g2_nor2_1 _6829_ (.A(_3396_),
    .B(_3519_),
    .Y(_2643_));
 sg13g2_o21ai_1 _6830_ (.B1(net1279),
    .Y(_2644_),
    .A1(_2577_),
    .A2(_2643_));
 sg13g2_nor2_1 _6831_ (.A(net1585),
    .B(net461),
    .Y(_2645_));
 sg13g2_a22oi_1 _6832_ (.Y(_0023_),
    .B1(net669),
    .B2(_2645_),
    .A2(_3517_),
    .A1(net1585));
 sg13g2_o21ai_1 _6833_ (.B1(net1268),
    .Y(_2646_),
    .A1(net1634),
    .A2(net1258));
 sg13g2_a21oi_1 _6834_ (.A1(net1622),
    .A2(net1264),
    .Y(_2647_),
    .B1(_2646_));
 sg13g2_a21oi_1 _6835_ (.A1(_3396_),
    .A2(_2534_),
    .Y(_2648_),
    .B1(_2647_));
 sg13g2_o21ai_1 _6836_ (.B1(_2647_),
    .Y(_2649_),
    .A1(\s0.was_valid_out[5] [0]),
    .A2(net1263));
 sg13g2_nor2_1 _6837_ (.A(net1258),
    .B(_2646_),
    .Y(_2650_));
 sg13g2_o21ai_1 _6838_ (.B1(net1167),
    .Y(_2651_),
    .A1(\s0.was_valid_out[5] [0]),
    .A2(net1274));
 sg13g2_nand2_1 _6839_ (.Y(_2652_),
    .A(_2649_),
    .B(_2651_));
 sg13g2_o21ai_1 _6840_ (.B1(net1718),
    .Y(_2653_),
    .A1(_2650_),
    .A2(_2652_));
 sg13g2_a21oi_1 _6841_ (.A1(_3363_),
    .A2(_2648_),
    .Y(_0024_),
    .B1(_2653_));
 sg13g2_and2_1 _6842_ (.A(net1718),
    .B(_2648_),
    .X(_0025_));
 sg13g2_and2_1 _6843_ (.A(net1717),
    .B(net396),
    .X(_0026_));
 sg13g2_nand2_1 _6844_ (.Y(_2654_),
    .A(net1260),
    .B(net546));
 sg13g2_o21ai_1 _6845_ (.B1(_2654_),
    .Y(_2655_),
    .A1(net1260),
    .A2(_3523_));
 sg13g2_nor2b_1 _6846_ (.A(net1253),
    .B_N(net1345),
    .Y(_2656_));
 sg13g2_a21o_1 _6847_ (.A2(_2655_),
    .A1(net1253),
    .B1(_2656_),
    .X(_2657_));
 sg13g2_nand2b_1 _6848_ (.Y(_2658_),
    .B(net546),
    .A_N(net1272));
 sg13g2_a21oi_1 _6849_ (.A1(_2551_),
    .A2(_2658_),
    .Y(_2659_),
    .B1(net1265));
 sg13g2_a21oi_1 _6850_ (.A1(net1265),
    .A2(_2657_),
    .Y(_2660_),
    .B1(_2659_));
 sg13g2_mux2_1 _6851_ (.A0(\s0.data_out[5][0] ),
    .A1(\s0.data_out[6][0] ),
    .S(net1272),
    .X(_2661_));
 sg13g2_nand2_1 _6852_ (.Y(_2662_),
    .A(net1168),
    .B(_2661_));
 sg13g2_nor2b_1 _6853_ (.A(net1253),
    .B_N(net1349),
    .Y(_2663_));
 sg13g2_mux2_1 _6854_ (.A0(\s0.data_out[6][0] ),
    .A1(\s0.data_out[5][0] ),
    .S(net1260),
    .X(_2664_));
 sg13g2_a21oi_1 _6855_ (.A1(net1253),
    .A2(_2664_),
    .Y(_2665_),
    .B1(_2663_));
 sg13g2_nand2b_1 _6856_ (.Y(_2666_),
    .B(net1265),
    .A_N(_2665_));
 sg13g2_a221oi_1 _6857_ (.B2(_2666_),
    .C1(net1703),
    .B1(_2662_),
    .A1(net1692),
    .Y(_2667_),
    .A2(_2660_));
 sg13g2_nand2_1 _6858_ (.Y(_2668_),
    .A(net1260),
    .B(net646));
 sg13g2_o21ai_1 _6859_ (.B1(_2668_),
    .Y(_2669_),
    .A1(net1261),
    .A2(_3522_));
 sg13g2_nor2b_1 _6860_ (.A(net1253),
    .B_N(net1341),
    .Y(_2670_));
 sg13g2_a21oi_1 _6861_ (.A1(net1254),
    .A2(_2669_),
    .Y(_2671_),
    .B1(_2670_));
 sg13g2_o21ai_1 _6862_ (.B1(_2543_),
    .Y(_2672_),
    .A1(net1272),
    .A2(_3529_));
 sg13g2_nand2_1 _6863_ (.Y(_2673_),
    .A(net1168),
    .B(_2672_));
 sg13g2_o21ai_1 _6864_ (.B1(_2673_),
    .Y(_2674_),
    .A1(net1168),
    .A2(_2671_));
 sg13g2_or2_1 _6865_ (.X(_2675_),
    .B(_2674_),
    .A(net1561));
 sg13g2_xnor2_1 _6866_ (.Y(_2676_),
    .A(net1561),
    .B(_2674_));
 sg13g2_nand2_1 _6867_ (.Y(_2677_),
    .A(net1262),
    .B(\s0.data_out[5][3] ));
 sg13g2_o21ai_1 _6868_ (.B1(_2677_),
    .Y(_2678_),
    .A1(net1262),
    .A2(_3521_));
 sg13g2_nor2_1 _6869_ (.A(net1255),
    .B(net1162),
    .Y(_2679_));
 sg13g2_a21o_1 _6870_ (.A2(_2678_),
    .A1(net1255),
    .B1(_2679_),
    .X(_2680_));
 sg13g2_nand2b_1 _6871_ (.Y(_2681_),
    .B(\s0.data_out[5][3] ),
    .A_N(net1273));
 sg13g2_a21oi_1 _6872_ (.A1(_2566_),
    .A2(_2681_),
    .Y(_2682_),
    .B1(net1267));
 sg13g2_a21oi_1 _6873_ (.A1(net1267),
    .A2(_2680_),
    .Y(_2683_),
    .B1(_2682_));
 sg13g2_nor2_1 _6874_ (.A(net1676),
    .B(_2683_),
    .Y(_2684_));
 sg13g2_nor2_1 _6875_ (.A(net1692),
    .B(_2660_),
    .Y(_2685_));
 sg13g2_nor4_1 _6876_ (.A(_2667_),
    .B(_2676_),
    .C(_2684_),
    .D(_2685_),
    .Y(_2686_));
 sg13g2_nand2_1 _6877_ (.Y(_2687_),
    .A(net1676),
    .B(_2683_));
 sg13g2_o21ai_1 _6878_ (.B1(_2687_),
    .Y(_2688_),
    .A1(_2675_),
    .A2(_2684_));
 sg13g2_nand2_1 _6879_ (.Y(_2689_),
    .A(net1260),
    .B(net596));
 sg13g2_mux2_1 _6880_ (.A0(\s0.data_out[6][6] ),
    .A1(\s0.data_out[5][6] ),
    .S(net1263),
    .X(_2690_));
 sg13g2_nor2b_1 _6881_ (.A(net1256),
    .B_N(net1329),
    .Y(_2691_));
 sg13g2_a21o_1 _6882_ (.A2(_2690_),
    .A1(net1256),
    .B1(_2691_),
    .X(_2692_));
 sg13g2_nand2b_1 _6883_ (.Y(_2693_),
    .B(net596),
    .A_N(net1274));
 sg13g2_a21oi_1 _6884_ (.A1(_2582_),
    .A2(_2693_),
    .Y(_2694_),
    .B1(net1268));
 sg13g2_a21oi_1 _6885_ (.A1(net1268),
    .A2(_2692_),
    .Y(_2695_),
    .B1(_2694_));
 sg13g2_nand2_1 _6886_ (.Y(_2696_),
    .A(net1262),
    .B(net528));
 sg13g2_mux2_1 _6887_ (.A0(\s0.data_out[6][7] ),
    .A1(\s0.data_out[5][7] ),
    .S(net1263),
    .X(_2697_));
 sg13g2_nor2b_1 _6888_ (.A(net1256),
    .B_N(net1320),
    .Y(_2698_));
 sg13g2_a21o_1 _6889_ (.A2(_2697_),
    .A1(net1258),
    .B1(_2698_),
    .X(_2699_));
 sg13g2_nand2b_1 _6890_ (.Y(_2700_),
    .B(net528),
    .A_N(net1274));
 sg13g2_a21oi_1 _6891_ (.A1(_2575_),
    .A2(_2700_),
    .Y(_2701_),
    .B1(net1268));
 sg13g2_a21oi_1 _6892_ (.A1(net1268),
    .A2(_2699_),
    .Y(_2702_),
    .B1(_2701_));
 sg13g2_a22oi_1 _6893_ (.Y(_2703_),
    .B1(_2702_),
    .B2(net1638),
    .A2(_2695_),
    .A1(net1648));
 sg13g2_or2_1 _6894_ (.X(_2704_),
    .B(_2695_),
    .A(net1649));
 sg13g2_nor2_1 _6895_ (.A(net1638),
    .B(_2702_),
    .Y(_2705_));
 sg13g2_nand3b_1 _6896_ (.B(_2703_),
    .C(_2704_),
    .Y(_2706_),
    .A_N(_2705_));
 sg13g2_nand2_1 _6897_ (.Y(_2707_),
    .A(net1263),
    .B(net651));
 sg13g2_mux2_1 _6898_ (.A0(\s0.data_out[6][5] ),
    .A1(\s0.data_out[5][5] ),
    .S(net1264),
    .X(_2708_));
 sg13g2_nor2b_1 _6899_ (.A(net1258),
    .B_N(net1331),
    .Y(_2709_));
 sg13g2_a21oi_1 _6900_ (.A1(net1257),
    .A2(_2708_),
    .Y(_2710_),
    .B1(_2709_));
 sg13g2_nand2b_1 _6901_ (.Y(_2711_),
    .B(net1269),
    .A_N(_2710_));
 sg13g2_o21ai_1 _6902_ (.B1(_2601_),
    .Y(_2712_),
    .A1(net1274),
    .A2(_3526_));
 sg13g2_nand2_1 _6903_ (.Y(_2713_),
    .A(net1167),
    .B(_2712_));
 sg13g2_nand3_1 _6904_ (.B(_2711_),
    .C(_2713_),
    .A(net1657),
    .Y(_2714_));
 sg13g2_nor2b_1 _6905_ (.A(net1257),
    .B_N(net1336),
    .Y(_2715_));
 sg13g2_nand2_1 _6906_ (.Y(_2716_),
    .A(net1263),
    .B(net751));
 sg13g2_mux2_1 _6907_ (.A0(\s0.data_out[6][4] ),
    .A1(\s0.data_out[5][4] ),
    .S(net1263),
    .X(_2717_));
 sg13g2_a21oi_1 _6908_ (.A1(net1257),
    .A2(_2717_),
    .Y(_2718_),
    .B1(_2715_));
 sg13g2_nand2b_1 _6909_ (.Y(_2719_),
    .B(net1269),
    .A_N(_2718_));
 sg13g2_o21ai_1 _6910_ (.B1(_2594_),
    .Y(_2720_),
    .A1(net1275),
    .A2(_3527_));
 sg13g2_nand2_1 _6911_ (.Y(_2721_),
    .A(net1167),
    .B(_2720_));
 sg13g2_nand3_1 _6912_ (.B(_2719_),
    .C(_2721_),
    .A(net1667),
    .Y(_2722_));
 sg13g2_nand2_1 _6913_ (.Y(_2723_),
    .A(_2714_),
    .B(_2722_));
 sg13g2_a21oi_1 _6914_ (.A1(_2719_),
    .A2(_2721_),
    .Y(_2724_),
    .B1(net1667));
 sg13g2_a21oi_1 _6915_ (.A1(_2711_),
    .A2(_2713_),
    .Y(_2725_),
    .B1(net1657));
 sg13g2_a21o_1 _6916_ (.A2(_2713_),
    .A1(_2711_),
    .B1(net1657),
    .X(_2726_));
 sg13g2_nor4_1 _6917_ (.A(_2706_),
    .B(_2723_),
    .C(_2724_),
    .D(_2725_),
    .Y(_2727_));
 sg13g2_o21ai_1 _6918_ (.B1(_2727_),
    .Y(_2728_),
    .A1(_2686_),
    .A2(_2688_));
 sg13g2_a21oi_1 _6919_ (.A1(_2714_),
    .A2(_2722_),
    .Y(_2729_),
    .B1(_2706_));
 sg13g2_o21ai_1 _6920_ (.B1(_2648_),
    .Y(_2730_),
    .A1(_2703_),
    .A2(_2705_));
 sg13g2_a21oi_1 _6921_ (.A1(_2726_),
    .A2(_2729_),
    .Y(_2731_),
    .B1(_2730_));
 sg13g2_or2_1 _6922_ (.X(_2732_),
    .B(net1556),
    .A(net397));
 sg13g2_a21oi_1 _6923_ (.A1(_2728_),
    .A2(_2731_),
    .Y(_0027_),
    .B1(_2732_));
 sg13g2_and2_1 _6924_ (.A(net1253),
    .B(net839),
    .X(_2733_));
 sg13g2_o21ai_1 _6925_ (.B1(net1265),
    .Y(_2734_),
    .A1(_2663_),
    .A2(_2733_));
 sg13g2_nand3_1 _6926_ (.B(_2662_),
    .C(_2734_),
    .A(net1715),
    .Y(_2735_));
 sg13g2_o21ai_1 _6927_ (.B1(_2735_),
    .Y(_2736_),
    .A1(net1715),
    .A2(net696));
 sg13g2_inv_1 _6928_ (.Y(_0028_),
    .A(_2736_));
 sg13g2_and2_1 _6929_ (.A(net1253),
    .B(net546),
    .X(_2737_));
 sg13g2_o21ai_1 _6930_ (.B1(net1265),
    .Y(_2738_),
    .A1(_2656_),
    .A2(_2737_));
 sg13g2_nor2_1 _6931_ (.A(net1583),
    .B(_2659_),
    .Y(_2739_));
 sg13g2_a22oi_1 _6932_ (.Y(_0029_),
    .B1(_2738_),
    .B2(_2739_),
    .A2(_3523_),
    .A1(net1583));
 sg13g2_a21oi_1 _6933_ (.A1(net1253),
    .A2(\s0.data_out[5][2] ),
    .Y(_2740_),
    .B1(_2670_));
 sg13g2_a21oi_1 _6934_ (.A1(net1168),
    .A2(_2672_),
    .Y(_2741_),
    .B1(net1584));
 sg13g2_o21ai_1 _6935_ (.B1(_2741_),
    .Y(_2742_),
    .A1(net1168),
    .A2(_2740_));
 sg13g2_o21ai_1 _6936_ (.B1(_2742_),
    .Y(_2743_),
    .A1(net1715),
    .A2(net549));
 sg13g2_inv_1 _6937_ (.Y(_0030_),
    .A(net550));
 sg13g2_and2_1 _6938_ (.A(net1255),
    .B(\s0.data_out[5][3] ),
    .X(_2744_));
 sg13g2_o21ai_1 _6939_ (.B1(net426),
    .Y(_2745_),
    .A1(_2679_),
    .A2(_2744_));
 sg13g2_nor2_1 _6940_ (.A(net1586),
    .B(_2682_),
    .Y(_2746_));
 sg13g2_a22oi_1 _6941_ (.Y(_0031_),
    .B1(net427),
    .B2(_2746_),
    .A2(_3521_),
    .A1(net1586));
 sg13g2_a21oi_1 _6942_ (.A1(net1257),
    .A2(\s0.data_out[5][4] ),
    .Y(_2747_),
    .B1(_2715_));
 sg13g2_a21oi_1 _6943_ (.A1(net1167),
    .A2(_2720_),
    .Y(_2748_),
    .B1(net1585));
 sg13g2_o21ai_1 _6944_ (.B1(_2748_),
    .Y(_2749_),
    .A1(net1167),
    .A2(_2747_));
 sg13g2_o21ai_1 _6945_ (.B1(_2749_),
    .Y(_2750_),
    .A1(net1718),
    .A2(net654));
 sg13g2_inv_1 _6946_ (.Y(_0032_),
    .A(net655));
 sg13g2_a21oi_1 _6947_ (.A1(net1257),
    .A2(net651),
    .Y(_2751_),
    .B1(_2709_));
 sg13g2_a21oi_1 _6948_ (.A1(net1167),
    .A2(_2712_),
    .Y(_2752_),
    .B1(net1586));
 sg13g2_o21ai_1 _6949_ (.B1(_2752_),
    .Y(_2753_),
    .A1(net1167),
    .A2(_2751_));
 sg13g2_o21ai_1 _6950_ (.B1(_2753_),
    .Y(_2754_),
    .A1(net1718),
    .A2(net800));
 sg13g2_inv_1 _6951_ (.Y(_0033_),
    .A(_2754_));
 sg13g2_and2_1 _6952_ (.A(net1256),
    .B(net596),
    .X(_2755_));
 sg13g2_o21ai_1 _6953_ (.B1(net1268),
    .Y(_2756_),
    .A1(_2691_),
    .A2(_2755_));
 sg13g2_nor2_1 _6954_ (.A(net1585),
    .B(_2694_),
    .Y(_2757_));
 sg13g2_a22oi_1 _6955_ (.Y(_0034_),
    .B1(_2756_),
    .B2(_2757_),
    .A2(_3520_),
    .A1(net1585));
 sg13g2_and2_1 _6956_ (.A(net1256),
    .B(net528),
    .X(_2758_));
 sg13g2_o21ai_1 _6957_ (.B1(net1268),
    .Y(_2759_),
    .A1(_2698_),
    .A2(_2758_));
 sg13g2_nor2_1 _6958_ (.A(net1585),
    .B(_2701_),
    .Y(_2760_));
 sg13g2_a22oi_1 _6959_ (.Y(_0035_),
    .B1(_2759_),
    .B2(_2760_),
    .A2(_3519_),
    .A1(net1585));
 sg13g2_o21ai_1 _6960_ (.B1(net1250),
    .Y(_2761_),
    .A1(net1627),
    .A2(net1242));
 sg13g2_nor2b_1 _6961_ (.A(net1627),
    .B_N(net1247),
    .Y(_2762_));
 sg13g2_nor2_1 _6962_ (.A(_2761_),
    .B(_2762_),
    .Y(_2763_));
 sg13g2_a21oi_1 _6963_ (.A1(net1622),
    .A2(net1260),
    .Y(_2764_),
    .B1(net1250));
 sg13g2_nor2_1 _6964_ (.A(_2763_),
    .B(_2764_),
    .Y(_2765_));
 sg13g2_o21ai_1 _6965_ (.B1(_2763_),
    .Y(_2766_),
    .A1(net416),
    .A2(net1247));
 sg13g2_nor2_1 _6966_ (.A(net1242),
    .B(_2761_),
    .Y(_2767_));
 sg13g2_nor2_1 _6967_ (.A(net416),
    .B(net1260),
    .Y(_2768_));
 sg13g2_o21ai_1 _6968_ (.B1(_2766_),
    .Y(_2769_),
    .A1(net1250),
    .A2(_2768_));
 sg13g2_o21ai_1 _6969_ (.B1(net1715),
    .Y(_2770_),
    .A1(_2767_),
    .A2(_2769_));
 sg13g2_a21oi_1 _6970_ (.A1(_3362_),
    .A2(_2765_),
    .Y(_0036_),
    .B1(_2770_));
 sg13g2_nor3_1 _6971_ (.A(net1579),
    .B(_2763_),
    .C(_2764_),
    .Y(_0037_));
 sg13g2_and2_1 _6972_ (.A(net1706),
    .B(net380),
    .X(_0038_));
 sg13g2_mux2_1 _6973_ (.A0(\s0.data_out[5][2] ),
    .A1(\s0.data_out[4][2] ),
    .S(net1247),
    .X(_2771_));
 sg13g2_nor2b_1 _6974_ (.A(net1241),
    .B_N(net1341),
    .Y(_2772_));
 sg13g2_a21o_1 _6975_ (.A2(_2771_),
    .A1(net1241),
    .B1(_2772_),
    .X(_2773_));
 sg13g2_nand2b_1 _6976_ (.Y(_2774_),
    .B(\s0.data_out[4][2] ),
    .A_N(net1261));
 sg13g2_a21oi_1 _6977_ (.A1(_2668_),
    .A2(_2774_),
    .Y(_2775_),
    .B1(net1252));
 sg13g2_a21oi_1 _6978_ (.A1(net1252),
    .A2(_2773_),
    .Y(_2776_),
    .B1(_2775_));
 sg13g2_or2_1 _6979_ (.X(_2777_),
    .B(_2776_),
    .A(net1689));
 sg13g2_nand2_1 _6980_ (.Y(_2778_),
    .A(net1247),
    .B(\s0.data_out[4][1] ));
 sg13g2_o21ai_1 _6981_ (.B1(_2778_),
    .Y(_2779_),
    .A1(net1247),
    .A2(_3530_));
 sg13g2_nor2b_1 _6982_ (.A(net1241),
    .B_N(net1345),
    .Y(_2780_));
 sg13g2_a21o_1 _6983_ (.A2(_2779_),
    .A1(net1241),
    .B1(_2780_),
    .X(_2781_));
 sg13g2_nand2b_1 _6984_ (.Y(_2782_),
    .B(\s0.data_out[4][1] ),
    .A_N(net1261));
 sg13g2_a21oi_1 _6985_ (.A1(_2654_),
    .A2(_2782_),
    .Y(_2783_),
    .B1(net1254));
 sg13g2_a21oi_1 _6986_ (.A1(net1252),
    .A2(_2781_),
    .Y(_2784_),
    .B1(_2783_));
 sg13g2_mux2_1 _6987_ (.A0(\s0.data_out[5][0] ),
    .A1(\s0.data_out[4][0] ),
    .S(net1247),
    .X(_2785_));
 sg13g2_nor2b_1 _6988_ (.A(net1241),
    .B_N(net1349),
    .Y(_2786_));
 sg13g2_a21oi_1 _6989_ (.A1(net1241),
    .A2(_2785_),
    .Y(_2787_),
    .B1(_2786_));
 sg13g2_nand2b_1 _6990_ (.Y(_2788_),
    .B(net1252),
    .A_N(_2787_));
 sg13g2_mux2_1 _6991_ (.A0(\s0.data_out[4][0] ),
    .A1(\s0.data_out[5][0] ),
    .S(net1261),
    .X(_2789_));
 sg13g2_nand2b_1 _6992_ (.Y(_2790_),
    .B(_2789_),
    .A_N(net1252));
 sg13g2_a221oi_1 _6993_ (.B2(_2790_),
    .C1(net1700),
    .B1(_2788_),
    .A1(net1692),
    .Y(_2791_),
    .A2(_2784_));
 sg13g2_o21ai_1 _6994_ (.B1(_2777_),
    .Y(_2792_),
    .A1(net1692),
    .A2(_2784_));
 sg13g2_nand2_1 _6995_ (.Y(_2793_),
    .A(net1247),
    .B(net495));
 sg13g2_o21ai_1 _6996_ (.B1(_2793_),
    .Y(_2794_),
    .A1(net1248),
    .A2(_3528_));
 sg13g2_nor2_1 _6997_ (.A(net1243),
    .B(net1160),
    .Y(_2795_));
 sg13g2_a21o_1 _6998_ (.A2(_2794_),
    .A1(net1243),
    .B1(_2795_),
    .X(_2796_));
 sg13g2_nand2b_1 _6999_ (.Y(_2797_),
    .B(net495),
    .A_N(net1262));
 sg13g2_a21oi_1 _7000_ (.A1(_2677_),
    .A2(_2797_),
    .Y(_2798_),
    .B1(net1250));
 sg13g2_a21oi_1 _7001_ (.A1(net1251),
    .A2(_2796_),
    .Y(_2799_),
    .B1(_2798_));
 sg13g2_a22oi_1 _7002_ (.Y(_2800_),
    .B1(_2799_),
    .B2(net1676),
    .A2(_2776_),
    .A1(net1685));
 sg13g2_o21ai_1 _7003_ (.B1(_2800_),
    .Y(_2801_),
    .A1(_2791_),
    .A2(_2792_));
 sg13g2_nand2_1 _7004_ (.Y(_2802_),
    .A(net1245),
    .B(net624));
 sg13g2_mux2_1 _7005_ (.A0(\s0.data_out[5][7] ),
    .A1(\s0.data_out[4][7] ),
    .S(net1248),
    .X(_2803_));
 sg13g2_nor2b_1 _7006_ (.A(net1243),
    .B_N(net1320),
    .Y(_2804_));
 sg13g2_a21o_1 _7007_ (.A2(_2803_),
    .A1(net1243),
    .B1(_2804_),
    .X(_2805_));
 sg13g2_nand2b_1 _7008_ (.Y(_2806_),
    .B(\s0.data_out[4][7] ),
    .A_N(net1262));
 sg13g2_a21oi_1 _7009_ (.A1(_2696_),
    .A2(_2806_),
    .Y(_2807_),
    .B1(net1251));
 sg13g2_a21oi_1 _7010_ (.A1(net1251),
    .A2(_2805_),
    .Y(_2808_),
    .B1(_2807_));
 sg13g2_nand2_1 _7011_ (.Y(_2809_),
    .A(net1245),
    .B(net558));
 sg13g2_mux2_1 _7012_ (.A0(\s0.data_out[5][6] ),
    .A1(\s0.data_out[4][6] ),
    .S(net1247),
    .X(_2810_));
 sg13g2_nor2b_1 _7013_ (.A(net1242),
    .B_N(net1325),
    .Y(_2811_));
 sg13g2_a21o_1 _7014_ (.A2(_2810_),
    .A1(net1242),
    .B1(_2811_),
    .X(_2812_));
 sg13g2_nand2b_1 _7015_ (.Y(_2813_),
    .B(net558),
    .A_N(net1260));
 sg13g2_a21oi_1 _7016_ (.A1(_2689_),
    .A2(_2813_),
    .Y(_2814_),
    .B1(net1250));
 sg13g2_a21oi_1 _7017_ (.A1(net1250),
    .A2(_2812_),
    .Y(_2815_),
    .B1(_2814_));
 sg13g2_a22oi_1 _7018_ (.Y(_2816_),
    .B1(_2815_),
    .B2(net1648),
    .A2(_2808_),
    .A1(net1638));
 sg13g2_or2_1 _7019_ (.X(_2817_),
    .B(_2815_),
    .A(net1649));
 sg13g2_nor2_1 _7020_ (.A(net1638),
    .B(_2808_),
    .Y(_2818_));
 sg13g2_nand3b_1 _7021_ (.B(_2816_),
    .C(_2817_),
    .Y(_2819_),
    .A_N(_2818_));
 sg13g2_mux2_1 _7022_ (.A0(\s0.data_out[5][4] ),
    .A1(\s0.data_out[4][4] ),
    .S(net1248),
    .X(_2820_));
 sg13g2_nor2b_1 _7023_ (.A(net1243),
    .B_N(net1336),
    .Y(_2821_));
 sg13g2_a21o_1 _7024_ (.A2(_2820_),
    .A1(net1243),
    .B1(_2821_),
    .X(_2822_));
 sg13g2_nand2b_1 _7025_ (.Y(_2823_),
    .B(net642),
    .A_N(net1263));
 sg13g2_a21oi_1 _7026_ (.A1(_2716_),
    .A2(_2823_),
    .Y(_2824_),
    .B1(net1257));
 sg13g2_a21oi_1 _7027_ (.A1(net1257),
    .A2(_2822_),
    .Y(_2825_),
    .B1(_2824_));
 sg13g2_nand2_1 _7028_ (.Y(_2826_),
    .A(net1246),
    .B(\s0.data_out[4][5] ));
 sg13g2_mux2_1 _7029_ (.A0(\s0.data_out[5][5] ),
    .A1(\s0.data_out[4][5] ),
    .S(net1248),
    .X(_2827_));
 sg13g2_nor2b_1 _7030_ (.A(net1243),
    .B_N(net1330),
    .Y(_2828_));
 sg13g2_a21o_1 _7031_ (.A2(_2827_),
    .A1(net1243),
    .B1(_2828_),
    .X(_2829_));
 sg13g2_nand2b_1 _7032_ (.Y(_2830_),
    .B(\s0.data_out[4][5] ),
    .A_N(net1263));
 sg13g2_a21oi_1 _7033_ (.A1(_2707_),
    .A2(_2830_),
    .Y(_2831_),
    .B1(net1256));
 sg13g2_a21oi_1 _7034_ (.A1(net1256),
    .A2(_2829_),
    .Y(_2832_),
    .B1(_2831_));
 sg13g2_a22oi_1 _7035_ (.Y(_2833_),
    .B1(_2832_),
    .B2(net1657),
    .A2(_2825_),
    .A1(net1668));
 sg13g2_nor2_1 _7036_ (.A(net1676),
    .B(_2799_),
    .Y(_2834_));
 sg13g2_nor2_1 _7037_ (.A(net1657),
    .B(_2832_),
    .Y(_2835_));
 sg13g2_o21ai_1 _7038_ (.B1(_2833_),
    .Y(_2836_),
    .A1(net1668),
    .A2(_2825_));
 sg13g2_nor4_1 _7039_ (.A(_2819_),
    .B(_2834_),
    .C(_2835_),
    .D(_2836_),
    .Y(_2837_));
 sg13g2_nand2_1 _7040_ (.Y(_2838_),
    .A(_2801_),
    .B(_2837_));
 sg13g2_nor3_1 _7041_ (.A(_2819_),
    .B(_2833_),
    .C(_2835_),
    .Y(_2839_));
 sg13g2_o21ai_1 _7042_ (.B1(_2765_),
    .Y(_2840_),
    .A1(_2816_),
    .A2(_2818_));
 sg13g2_nor2_1 _7043_ (.A(_2839_),
    .B(_2840_),
    .Y(_2841_));
 sg13g2_or2_1 _7044_ (.X(_2842_),
    .B(net1556),
    .A(net396));
 sg13g2_a21oi_1 _7045_ (.A1(_2838_),
    .A2(_2841_),
    .Y(_0039_),
    .B1(_2842_));
 sg13g2_and2_1 _7046_ (.A(net1241),
    .B(\s0.data_out[4][0] ),
    .X(_2843_));
 sg13g2_o21ai_1 _7047_ (.B1(net1252),
    .Y(_2844_),
    .A1(_2786_),
    .A2(_2843_));
 sg13g2_nand3_1 _7048_ (.B(_2790_),
    .C(_2844_),
    .A(net1715),
    .Y(_2845_));
 sg13g2_o21ai_1 _7049_ (.B1(_2845_),
    .Y(_2846_),
    .A1(net1715),
    .A2(net757));
 sg13g2_inv_1 _7050_ (.Y(_0040_),
    .A(_2846_));
 sg13g2_and2_1 _7051_ (.A(net1241),
    .B(\s0.data_out[4][1] ),
    .X(_2847_));
 sg13g2_o21ai_1 _7052_ (.B1(net1252),
    .Y(_2848_),
    .A1(_2780_),
    .A2(_2847_));
 sg13g2_nor2_1 _7053_ (.A(net1583),
    .B(_2783_),
    .Y(_2849_));
 sg13g2_a22oi_1 _7054_ (.Y(_0041_),
    .B1(_2848_),
    .B2(_2849_),
    .A2(_3530_),
    .A1(net1583));
 sg13g2_and2_1 _7055_ (.A(net1242),
    .B(\s0.data_out[4][2] ),
    .X(_2850_));
 sg13g2_o21ai_1 _7056_ (.B1(net1252),
    .Y(_2851_),
    .A1(_2772_),
    .A2(_2850_));
 sg13g2_nor2_1 _7057_ (.A(net1583),
    .B(_2775_),
    .Y(_2852_));
 sg13g2_a22oi_1 _7058_ (.Y(_0042_),
    .B1(_2851_),
    .B2(_2852_),
    .A2(_3529_),
    .A1(net1579));
 sg13g2_nor2_1 _7059_ (.A(net1165),
    .B(_3533_),
    .Y(_2853_));
 sg13g2_o21ai_1 _7060_ (.B1(net1250),
    .Y(_2854_),
    .A1(_2795_),
    .A2(_2853_));
 sg13g2_nor2_1 _7061_ (.A(net1584),
    .B(net496),
    .Y(_2855_));
 sg13g2_a22oi_1 _7062_ (.Y(_0043_),
    .B1(_2854_),
    .B2(_2855_),
    .A2(_3528_),
    .A1(net1584));
 sg13g2_and2_1 _7063_ (.A(net1244),
    .B(net642),
    .X(_2856_));
 sg13g2_o21ai_1 _7064_ (.B1(net1257),
    .Y(_2857_),
    .A1(_2821_),
    .A2(_2856_));
 sg13g2_nor2_1 _7065_ (.A(net1584),
    .B(_2824_),
    .Y(_2858_));
 sg13g2_a22oi_1 _7066_ (.Y(_0044_),
    .B1(_2857_),
    .B2(_2858_),
    .A2(_3527_),
    .A1(net1586));
 sg13g2_and2_1 _7067_ (.A(net1244),
    .B(\s0.data_out[4][5] ),
    .X(_2859_));
 sg13g2_o21ai_1 _7068_ (.B1(net1256),
    .Y(_2860_),
    .A1(_2828_),
    .A2(_2859_));
 sg13g2_nor2_1 _7069_ (.A(net1584),
    .B(_2831_),
    .Y(_2861_));
 sg13g2_a22oi_1 _7070_ (.Y(_0045_),
    .B1(_2860_),
    .B2(_2861_),
    .A2(_3526_),
    .A1(net1585));
 sg13g2_nor2_1 _7071_ (.A(net1166),
    .B(_3532_),
    .Y(_2862_));
 sg13g2_o21ai_1 _7072_ (.B1(net1250),
    .Y(_2863_),
    .A1(_2811_),
    .A2(_2862_));
 sg13g2_nor2_1 _7073_ (.A(net1584),
    .B(_2814_),
    .Y(_2864_));
 sg13g2_a22oi_1 _7074_ (.Y(_0046_),
    .B1(_2863_),
    .B2(_2864_),
    .A2(_3525_),
    .A1(net1579));
 sg13g2_nor2_1 _7075_ (.A(net1165),
    .B(_3531_),
    .Y(_2865_));
 sg13g2_o21ai_1 _7076_ (.B1(net1251),
    .Y(_2866_),
    .A1(_2804_),
    .A2(_2865_));
 sg13g2_nor2_1 _7077_ (.A(net1584),
    .B(_2807_),
    .Y(_2867_));
 sg13g2_a22oi_1 _7078_ (.Y(_0047_),
    .B1(_2866_),
    .B2(_2867_),
    .A2(_3524_),
    .A1(net1584));
 sg13g2_o21ai_1 _7079_ (.B1(net1239),
    .Y(_2868_),
    .A1(net1627),
    .A2(net1231));
 sg13g2_nand2_1 _7080_ (.Y(_2869_),
    .A(net1621),
    .B(net1238));
 sg13g2_a21oi_1 _7081_ (.A1(net1621),
    .A2(net1237),
    .Y(_2870_),
    .B1(_2868_));
 sg13g2_nor2_1 _7082_ (.A(net1239),
    .B(_2762_),
    .Y(_2871_));
 sg13g2_nor2_1 _7083_ (.A(_2870_),
    .B(_2871_),
    .Y(_2872_));
 sg13g2_o21ai_1 _7084_ (.B1(_2870_),
    .Y(_2873_),
    .A1(net406),
    .A2(net1237));
 sg13g2_nor2_1 _7085_ (.A(net1231),
    .B(_2868_),
    .Y(_2874_));
 sg13g2_o21ai_1 _7086_ (.B1(net1164),
    .Y(_2875_),
    .A1(net406),
    .A2(net1245));
 sg13g2_nand2_1 _7087_ (.Y(_2876_),
    .A(_2873_),
    .B(_2875_));
 sg13g2_o21ai_1 _7088_ (.B1(net1706),
    .Y(_2877_),
    .A1(_2874_),
    .A2(_2876_));
 sg13g2_a21oi_1 _7089_ (.A1(_3361_),
    .A2(_2872_),
    .Y(_0048_),
    .B1(_2877_));
 sg13g2_nor3_1 _7090_ (.A(net1570),
    .B(_2870_),
    .C(_2871_),
    .Y(_0049_));
 sg13g2_and2_1 _7091_ (.A(net1705),
    .B(net377),
    .X(_0050_));
 sg13g2_mux2_1 _7092_ (.A0(\s0.data_out[4][2] ),
    .A1(\s0.data_out[3][2] ),
    .S(net1237),
    .X(_2878_));
 sg13g2_nor2b_1 _7093_ (.A(net1230),
    .B_N(net1340),
    .Y(_2879_));
 sg13g2_a21oi_1 _7094_ (.A1(net1231),
    .A2(_2878_),
    .Y(_2880_),
    .B1(_2879_));
 sg13g2_mux2_1 _7095_ (.A0(\s0.data_out[3][2] ),
    .A1(\s0.data_out[4][2] ),
    .S(net1245),
    .X(_2881_));
 sg13g2_nand2_1 _7096_ (.Y(_2882_),
    .A(net1163),
    .B(_2881_));
 sg13g2_o21ai_1 _7097_ (.B1(_2882_),
    .Y(_2883_),
    .A1(net1164),
    .A2(_2880_));
 sg13g2_mux2_1 _7098_ (.A0(\s0.data_out[4][1] ),
    .A1(\s0.data_out[3][1] ),
    .S(net1237),
    .X(_2884_));
 sg13g2_nor2b_1 _7099_ (.A(net1230),
    .B_N(net1344),
    .Y(_2885_));
 sg13g2_a21oi_1 _7100_ (.A1(net1230),
    .A2(_2884_),
    .Y(_2886_),
    .B1(_2885_));
 sg13g2_nand2b_1 _7101_ (.Y(_2887_),
    .B(net1239),
    .A_N(_2886_));
 sg13g2_mux2_1 _7102_ (.A0(\s0.data_out[3][1] ),
    .A1(\s0.data_out[4][1] ),
    .S(net1245),
    .X(_2888_));
 sg13g2_nand2_1 _7103_ (.Y(_2889_),
    .A(net1164),
    .B(_2888_));
 sg13g2_nand3_1 _7104_ (.B(_2887_),
    .C(_2889_),
    .A(net1690),
    .Y(_2890_));
 sg13g2_mux2_1 _7105_ (.A0(\s0.data_out[4][0] ),
    .A1(\s0.data_out[3][0] ),
    .S(net1237),
    .X(_2891_));
 sg13g2_nor2b_1 _7106_ (.A(net1230),
    .B_N(net1348),
    .Y(_2892_));
 sg13g2_a21oi_1 _7107_ (.A1(net1230),
    .A2(_2891_),
    .Y(_2893_),
    .B1(_2892_));
 sg13g2_mux2_1 _7108_ (.A0(\s0.data_out[3][0] ),
    .A1(\s0.data_out[4][0] ),
    .S(net1245),
    .X(_2894_));
 sg13g2_nand2_1 _7109_ (.Y(_2895_),
    .A(net1163),
    .B(_2894_));
 sg13g2_o21ai_1 _7110_ (.B1(_2895_),
    .Y(_2896_),
    .A1(net1163),
    .A2(_2893_));
 sg13g2_and2_1 _7111_ (.A(net1559),
    .B(_2896_),
    .X(_2897_));
 sg13g2_a21oi_1 _7112_ (.A1(_2887_),
    .A2(_2889_),
    .Y(_2898_),
    .B1(net1690));
 sg13g2_a221oi_1 _7113_ (.B2(_2897_),
    .C1(_2898_),
    .B1(_2890_),
    .A1(net1560),
    .Y(_2899_),
    .A2(_2883_));
 sg13g2_nand2_1 _7114_ (.Y(_2900_),
    .A(net1236),
    .B(net501));
 sg13g2_mux2_1 _7115_ (.A0(\s0.data_out[4][3] ),
    .A1(\s0.data_out[3][3] ),
    .S(net1236),
    .X(_2901_));
 sg13g2_nor2b_1 _7116_ (.A(net1232),
    .B_N(net1339),
    .Y(_2902_));
 sg13g2_a21o_1 _7117_ (.A2(_2901_),
    .A1(net1232),
    .B1(_2902_),
    .X(_2903_));
 sg13g2_nand2b_1 _7118_ (.Y(_2904_),
    .B(net501),
    .A_N(net1246));
 sg13g2_a21oi_1 _7119_ (.A1(_2793_),
    .A2(_2904_),
    .Y(_2905_),
    .B1(net1240));
 sg13g2_a21oi_1 _7120_ (.A1(net1240),
    .A2(_2903_),
    .Y(_2906_),
    .B1(_2905_));
 sg13g2_nand2_1 _7121_ (.Y(_2907_),
    .A(net1674),
    .B(_2906_));
 sg13g2_o21ai_1 _7122_ (.B1(_2907_),
    .Y(_2908_),
    .A1(net1560),
    .A2(_2883_));
 sg13g2_nand2_1 _7123_ (.Y(_2909_),
    .A(net1236),
    .B(net812));
 sg13g2_mux2_1 _7124_ (.A0(\s0.data_out[4][5] ),
    .A1(\s0.data_out[3][5] ),
    .S(net1236),
    .X(_2910_));
 sg13g2_nor2b_1 _7125_ (.A(net1232),
    .B_N(net1330),
    .Y(_2911_));
 sg13g2_a21oi_1 _7126_ (.A1(net1232),
    .A2(_2910_),
    .Y(_2912_),
    .B1(_2911_));
 sg13g2_nand2b_1 _7127_ (.Y(_2913_),
    .B(net1239),
    .A_N(_2912_));
 sg13g2_o21ai_1 _7128_ (.B1(_2826_),
    .Y(_2914_),
    .A1(net1246),
    .A2(_3536_));
 sg13g2_nand2_1 _7129_ (.Y(_2915_),
    .A(net1166),
    .B(_2914_));
 sg13g2_and3_1 _7130_ (.X(_2916_),
    .A(net1655),
    .B(_2913_),
    .C(_2915_));
 sg13g2_nor2_1 _7131_ (.A(net1674),
    .B(_2906_),
    .Y(_2917_));
 sg13g2_nor2_1 _7132_ (.A(_2916_),
    .B(_2917_),
    .Y(_2918_));
 sg13g2_a21o_1 _7133_ (.A2(_2915_),
    .A1(_2913_),
    .B1(net1655),
    .X(_2919_));
 sg13g2_nor2b_1 _7134_ (.A(net1232),
    .B_N(net1335),
    .Y(_2920_));
 sg13g2_nand2_1 _7135_ (.Y(_2921_),
    .A(\s0.valid_out[3] [0]),
    .B(\s0.data_out[3][4] ));
 sg13g2_mux2_1 _7136_ (.A0(\s0.data_out[4][4] ),
    .A1(\s0.data_out[3][4] ),
    .S(net1236),
    .X(_2922_));
 sg13g2_a21oi_1 _7137_ (.A1(net1232),
    .A2(_2922_),
    .Y(_2923_),
    .B1(_2920_));
 sg13g2_mux2_1 _7138_ (.A0(\s0.data_out[3][4] ),
    .A1(\s0.data_out[4][4] ),
    .S(net1245),
    .X(_2924_));
 sg13g2_nand2_1 _7139_ (.Y(_2925_),
    .A(net1165),
    .B(_2924_));
 sg13g2_o21ai_1 _7140_ (.B1(_2925_),
    .Y(_2926_),
    .A1(net1165),
    .A2(_2923_));
 sg13g2_nor2_1 _7141_ (.A(_3406_),
    .B(_2926_),
    .Y(_2927_));
 sg13g2_xnor2_1 _7142_ (.Y(_2928_),
    .A(net1665),
    .B(_2926_));
 sg13g2_nand3_1 _7143_ (.B(_2919_),
    .C(_2928_),
    .A(_2918_),
    .Y(_2929_));
 sg13g2_nand2_1 _7144_ (.Y(_2930_),
    .A(net1238),
    .B(net634));
 sg13g2_mux2_1 _7145_ (.A0(\s0.data_out[4][7] ),
    .A1(\s0.data_out[3][7] ),
    .S(net1236),
    .X(_2931_));
 sg13g2_nor2b_1 _7146_ (.A(net1231),
    .B_N(net1320),
    .Y(_2932_));
 sg13g2_a21o_1 _7147_ (.A2(_2931_),
    .A1(net1231),
    .B1(_2932_),
    .X(_2933_));
 sg13g2_nand2b_1 _7148_ (.Y(_2934_),
    .B(\s0.data_out[3][7] ),
    .A_N(net1246));
 sg13g2_a21oi_1 _7149_ (.A1(_2802_),
    .A2(_2934_),
    .Y(_2935_),
    .B1(net1240));
 sg13g2_a21oi_1 _7150_ (.A1(net1240),
    .A2(_2933_),
    .Y(_2936_),
    .B1(_2935_));
 sg13g2_mux2_1 _7151_ (.A0(\s0.data_out[4][6] ),
    .A1(\s0.data_out[3][6] ),
    .S(net1237),
    .X(_2937_));
 sg13g2_nor2b_1 _7152_ (.A(net1231),
    .B_N(net1325),
    .Y(_2938_));
 sg13g2_a21o_1 _7153_ (.A2(_2937_),
    .A1(net1231),
    .B1(_2938_),
    .X(_2939_));
 sg13g2_nand2b_1 _7154_ (.Y(_2940_),
    .B(\s0.data_out[3][6] ),
    .A_N(net1245));
 sg13g2_a21oi_1 _7155_ (.A1(_2809_),
    .A2(_2940_),
    .Y(_2941_),
    .B1(net1239));
 sg13g2_a21oi_1 _7156_ (.A1(net1239),
    .A2(_2939_),
    .Y(_2942_),
    .B1(_2941_));
 sg13g2_a22oi_1 _7157_ (.Y(_2943_),
    .B1(_2942_),
    .B2(net1646),
    .A2(_2936_),
    .A1(net1636));
 sg13g2_or2_1 _7158_ (.X(_2944_),
    .B(_2942_),
    .A(net1647));
 sg13g2_nor2_1 _7159_ (.A(net1636),
    .B(_2936_),
    .Y(_2945_));
 sg13g2_or2_1 _7160_ (.X(_2946_),
    .B(_2936_),
    .A(net1636));
 sg13g2_and3_1 _7161_ (.X(_2947_),
    .A(_2943_),
    .B(_2944_),
    .C(_2946_));
 sg13g2_o21ai_1 _7162_ (.B1(_2947_),
    .Y(_2948_),
    .A1(_2899_),
    .A2(_2908_));
 sg13g2_a21o_1 _7163_ (.A2(_2927_),
    .A1(_2919_),
    .B1(_2916_),
    .X(_2949_));
 sg13g2_o21ai_1 _7164_ (.B1(_2872_),
    .Y(_2950_),
    .A1(_2943_),
    .A2(_2945_));
 sg13g2_a21oi_1 _7165_ (.A1(_2947_),
    .A2(_2949_),
    .Y(_2951_),
    .B1(_2950_));
 sg13g2_o21ai_1 _7166_ (.B1(_2951_),
    .Y(_2952_),
    .A1(_2929_),
    .A2(_2948_));
 sg13g2_nor2_1 _7167_ (.A(net380),
    .B(net1555),
    .Y(_2953_));
 sg13g2_and2_1 _7168_ (.A(_2952_),
    .B(_2953_),
    .X(_0051_));
 sg13g2_a21oi_1 _7169_ (.A1(net1230),
    .A2(\s0.data_out[3][0] ),
    .Y(_2954_),
    .B1(_2892_));
 sg13g2_a21oi_1 _7170_ (.A1(net1163),
    .A2(_2894_),
    .Y(_2955_),
    .B1(net1570));
 sg13g2_o21ai_1 _7171_ (.B1(_2955_),
    .Y(_2956_),
    .A1(net1163),
    .A2(_2954_));
 sg13g2_o21ai_1 _7172_ (.B1(_2956_),
    .Y(_2957_),
    .A1(net1706),
    .A2(net710));
 sg13g2_inv_1 _7173_ (.Y(_0052_),
    .A(net711));
 sg13g2_a21oi_1 _7174_ (.A1(net1230),
    .A2(\s0.data_out[3][1] ),
    .Y(_2958_),
    .B1(_2885_));
 sg13g2_a21oi_1 _7175_ (.A1(net1163),
    .A2(_2888_),
    .Y(_2959_),
    .B1(net1570));
 sg13g2_o21ai_1 _7176_ (.B1(_2959_),
    .Y(_2960_),
    .A1(net1163),
    .A2(_2958_));
 sg13g2_o21ai_1 _7177_ (.B1(_2960_),
    .Y(_2961_),
    .A1(net1706),
    .A2(net723));
 sg13g2_inv_1 _7178_ (.Y(_0053_),
    .A(net724));
 sg13g2_a21oi_1 _7179_ (.A1(net1230),
    .A2(net703),
    .Y(_2962_),
    .B1(_2879_));
 sg13g2_a21oi_1 _7180_ (.A1(net1164),
    .A2(_2881_),
    .Y(_2963_),
    .B1(net1570));
 sg13g2_o21ai_1 _7181_ (.B1(_2963_),
    .Y(_2964_),
    .A1(net1163),
    .A2(_2962_));
 sg13g2_o21ai_1 _7182_ (.B1(_2964_),
    .Y(_2965_),
    .A1(net1706),
    .A2(net748));
 sg13g2_inv_1 _7183_ (.Y(_0054_),
    .A(_2965_));
 sg13g2_nor2_1 _7184_ (.A(net1184),
    .B(_3534_),
    .Y(_2966_));
 sg13g2_o21ai_1 _7185_ (.B1(net1240),
    .Y(_2967_),
    .A1(_2902_),
    .A2(_2966_));
 sg13g2_nor2_1 _7186_ (.A(net1574),
    .B(_2905_),
    .Y(_2968_));
 sg13g2_a22oi_1 _7187_ (.Y(_0055_),
    .B1(_2967_),
    .B2(_2968_),
    .A2(_3533_),
    .A1(net1574));
 sg13g2_a21oi_1 _7188_ (.A1(net1232),
    .A2(\s0.data_out[3][4] ),
    .Y(_2969_),
    .B1(_2920_));
 sg13g2_a21oi_1 _7189_ (.A1(net1165),
    .A2(_2924_),
    .Y(_2970_),
    .B1(net1574));
 sg13g2_o21ai_1 _7190_ (.B1(_2970_),
    .Y(_2971_),
    .A1(net1165),
    .A2(_2969_));
 sg13g2_o21ai_1 _7191_ (.B1(_2971_),
    .Y(_2972_),
    .A1(net1713),
    .A2(net642));
 sg13g2_inv_1 _7192_ (.Y(_0056_),
    .A(net643));
 sg13g2_a21oi_1 _7193_ (.A1(net1232),
    .A2(\s0.data_out[3][5] ),
    .Y(_2973_),
    .B1(_2911_));
 sg13g2_a21oi_1 _7194_ (.A1(net1165),
    .A2(_2914_),
    .Y(_2974_),
    .B1(net1575));
 sg13g2_o21ai_1 _7195_ (.B1(_2974_),
    .Y(_2975_),
    .A1(net1165),
    .A2(_2973_));
 sg13g2_o21ai_1 _7196_ (.B1(_2975_),
    .Y(_2976_),
    .A1(net1713),
    .A2(net675));
 sg13g2_inv_1 _7197_ (.Y(_0057_),
    .A(net676));
 sg13g2_and2_1 _7198_ (.A(net1231),
    .B(\s0.data_out[3][6] ),
    .X(_2977_));
 sg13g2_o21ai_1 _7199_ (.B1(net1239),
    .Y(_2978_),
    .A1(_2938_),
    .A2(_2977_));
 sg13g2_nor2_1 _7200_ (.A(net1574),
    .B(_2941_),
    .Y(_2979_));
 sg13g2_a22oi_1 _7201_ (.Y(_0058_),
    .B1(_2978_),
    .B2(_2979_),
    .A2(_3532_),
    .A1(net1570));
 sg13g2_nor2_1 _7202_ (.A(net1184),
    .B(_3535_),
    .Y(_2980_));
 sg13g2_o21ai_1 _7203_ (.B1(net1240),
    .Y(_2981_),
    .A1(_2932_),
    .A2(_2980_));
 sg13g2_nor2_1 _7204_ (.A(net1574),
    .B(_2935_),
    .Y(_2982_));
 sg13g2_a22oi_1 _7205_ (.Y(_0059_),
    .B1(_2981_),
    .B2(_2982_),
    .A2(_3531_),
    .A1(net1574));
 sg13g2_o21ai_1 _7206_ (.B1(net1235),
    .Y(_2983_),
    .A1(net1628),
    .A2(net1220));
 sg13g2_nor2b_1 _7207_ (.A(net1628),
    .B_N(net1227),
    .Y(_2984_));
 sg13g2_nor2_1 _7208_ (.A(_2983_),
    .B(_2984_),
    .Y(_2985_));
 sg13g2_a21oi_1 _7209_ (.A1(net1183),
    .A2(_2869_),
    .Y(_2986_),
    .B1(_2985_));
 sg13g2_o21ai_1 _7210_ (.B1(_2985_),
    .Y(_2987_),
    .A1(\s0.was_valid_out[2] [0]),
    .A2(net1227));
 sg13g2_nor2_1 _7211_ (.A(net1220),
    .B(_2983_),
    .Y(_2988_));
 sg13g2_o21ai_1 _7212_ (.B1(net1184),
    .Y(_2989_),
    .A1(\s0.was_valid_out[2] [0]),
    .A2(net1238));
 sg13g2_nand2_1 _7213_ (.Y(_2990_),
    .A(_2987_),
    .B(_2989_));
 sg13g2_o21ai_1 _7214_ (.B1(net1708),
    .Y(_2991_),
    .A1(_2988_),
    .A2(_2990_));
 sg13g2_a21oi_1 _7215_ (.A1(_3360_),
    .A2(_2986_),
    .Y(_0060_),
    .B1(_2991_));
 sg13g2_and2_1 _7216_ (.A(net1704),
    .B(_2986_),
    .X(_0061_));
 sg13g2_and2_1 _7217_ (.A(net1709),
    .B(net372),
    .X(_0062_));
 sg13g2_nand2_1 _7218_ (.Y(_2992_),
    .A(net1226),
    .B(\s0.data_out[2][1] ));
 sg13g2_mux2_1 _7219_ (.A0(\s0.data_out[3][1] ),
    .A1(\s0.data_out[2][1] ),
    .S(net1227),
    .X(_2993_));
 sg13g2_nor2b_1 _7220_ (.A(net1219),
    .B_N(net1344),
    .Y(_2994_));
 sg13g2_a21oi_1 _7221_ (.A1(net1219),
    .A2(_2993_),
    .Y(_2995_),
    .B1(_2994_));
 sg13g2_mux2_1 _7222_ (.A0(\s0.data_out[2][1] ),
    .A1(\s0.data_out[3][1] ),
    .S(net1238),
    .X(_2996_));
 sg13g2_nand2_1 _7223_ (.Y(_2997_),
    .A(net1183),
    .B(_2996_));
 sg13g2_o21ai_1 _7224_ (.B1(_2997_),
    .Y(_2998_),
    .A1(net1183),
    .A2(_2995_));
 sg13g2_nor2_1 _7225_ (.A(_3415_),
    .B(_2998_),
    .Y(_2999_));
 sg13g2_mux2_1 _7226_ (.A0(\s0.data_out[3][0] ),
    .A1(\s0.data_out[2][0] ),
    .S(net1227),
    .X(_3000_));
 sg13g2_nor2b_1 _7227_ (.A(net1219),
    .B_N(net1348),
    .Y(_3001_));
 sg13g2_a21oi_1 _7228_ (.A1(net1219),
    .A2(_3000_),
    .Y(_3002_),
    .B1(_3001_));
 sg13g2_mux2_1 _7229_ (.A0(\s0.data_out[2][0] ),
    .A1(\s0.data_out[3][0] ),
    .S(net1238),
    .X(_3003_));
 sg13g2_nand2_1 _7230_ (.Y(_3004_),
    .A(net1183),
    .B(_3003_));
 sg13g2_o21ai_1 _7231_ (.B1(_3004_),
    .Y(_3005_),
    .A1(net1183),
    .A2(_3002_));
 sg13g2_mux2_1 _7232_ (.A0(\s0.data_out[3][2] ),
    .A1(\s0.data_out[2][2] ),
    .S(net1229),
    .X(_3006_));
 sg13g2_nor2b_1 _7233_ (.A(net1221),
    .B_N(net1340),
    .Y(_3007_));
 sg13g2_a21oi_1 _7234_ (.A1(net1221),
    .A2(_3006_),
    .Y(_3008_),
    .B1(_3007_));
 sg13g2_nor2_1 _7235_ (.A(net1184),
    .B(_3008_),
    .Y(_3009_));
 sg13g2_mux2_1 _7236_ (.A0(\s0.data_out[2][2] ),
    .A1(\s0.data_out[3][2] ),
    .S(net1238),
    .X(_3010_));
 sg13g2_a21oi_1 _7237_ (.A1(net1184),
    .A2(_3010_),
    .Y(_3011_),
    .B1(_3009_));
 sg13g2_nor2_1 _7238_ (.A(net1685),
    .B(_3011_),
    .Y(_3012_));
 sg13g2_a22oi_1 _7239_ (.Y(_3013_),
    .B1(_3005_),
    .B2(net1559),
    .A2(_2998_),
    .A1(_3415_));
 sg13g2_nor2_1 _7240_ (.A(_2999_),
    .B(_3013_),
    .Y(_3014_));
 sg13g2_nand2_1 _7241_ (.Y(_3015_),
    .A(net1228),
    .B(net784));
 sg13g2_o21ai_1 _7242_ (.B1(_3015_),
    .Y(_3016_),
    .A1(net1228),
    .A2(_3534_));
 sg13g2_nor2_1 _7243_ (.A(net1223),
    .B(net1160),
    .Y(_3017_));
 sg13g2_a21o_1 _7244_ (.A2(_3016_),
    .A1(net1221),
    .B1(_3017_),
    .X(_3018_));
 sg13g2_nand2b_1 _7245_ (.Y(_3019_),
    .B(net784),
    .A_N(net1236));
 sg13g2_a21oi_1 _7246_ (.A1(_2900_),
    .A2(_3019_),
    .Y(_3020_),
    .B1(net1233));
 sg13g2_a21oi_1 _7247_ (.A1(net1233),
    .A2(_3018_),
    .Y(_3021_),
    .B1(_3020_));
 sg13g2_a22oi_1 _7248_ (.Y(_3022_),
    .B1(_3021_),
    .B2(net1675),
    .A2(_3011_),
    .A1(net1685));
 sg13g2_o21ai_1 _7249_ (.B1(_3022_),
    .Y(_3023_),
    .A1(_3012_),
    .A2(_3014_));
 sg13g2_nand2_1 _7250_ (.Y(_3024_),
    .A(net1226),
    .B(\s0.data_out[2][6] ));
 sg13g2_mux2_1 _7251_ (.A0(\s0.data_out[3][6] ),
    .A1(\s0.data_out[2][6] ),
    .S(net1227),
    .X(_3025_));
 sg13g2_nor2b_1 _7252_ (.A(net1220),
    .B_N(net1326),
    .Y(_3026_));
 sg13g2_a21oi_1 _7253_ (.A1(net1219),
    .A2(_3025_),
    .Y(_3027_),
    .B1(_3026_));
 sg13g2_nand2b_1 _7254_ (.Y(_3028_),
    .B(net1235),
    .A_N(_3027_));
 sg13g2_mux2_1 _7255_ (.A0(\s0.data_out[2][6] ),
    .A1(\s0.data_out[3][6] ),
    .S(net1238),
    .X(_3029_));
 sg13g2_nand2_1 _7256_ (.Y(_3030_),
    .A(net1183),
    .B(_3029_));
 sg13g2_and2_1 _7257_ (.A(_3028_),
    .B(_3030_),
    .X(_3031_));
 sg13g2_nand2_1 _7258_ (.Y(_3032_),
    .A(net1226),
    .B(net542));
 sg13g2_mux2_1 _7259_ (.A0(\s0.data_out[3][7] ),
    .A1(\s0.data_out[2][7] ),
    .S(net1227),
    .X(_3033_));
 sg13g2_nor2b_1 _7260_ (.A(net1220),
    .B_N(net1321),
    .Y(_3034_));
 sg13g2_a21o_1 _7261_ (.A2(_3033_),
    .A1(net1220),
    .B1(_3034_),
    .X(_3035_));
 sg13g2_nand2b_1 _7262_ (.Y(_3036_),
    .B(net542),
    .A_N(net1238));
 sg13g2_a21oi_1 _7263_ (.A1(_2930_),
    .A2(_3036_),
    .Y(_3037_),
    .B1(net1235));
 sg13g2_a21oi_1 _7264_ (.A1(net1235),
    .A2(_3035_),
    .Y(_3038_),
    .B1(_3037_));
 sg13g2_a22oi_1 _7265_ (.Y(_3039_),
    .B1(_3038_),
    .B2(net1635),
    .A2(_3031_),
    .A1(net1647));
 sg13g2_nor2_1 _7266_ (.A(net1635),
    .B(_3038_),
    .Y(_3040_));
 sg13g2_a21oi_1 _7267_ (.A1(_3028_),
    .A2(_3030_),
    .Y(_3041_),
    .B1(net1647));
 sg13g2_nand2_1 _7268_ (.Y(_3042_),
    .A(net1228),
    .B(\s0.data_out[2][5] ));
 sg13g2_o21ai_1 _7269_ (.B1(_3042_),
    .Y(_3043_),
    .A1(net1228),
    .A2(_3536_));
 sg13g2_nor2b_1 _7270_ (.A(net1223),
    .B_N(net1331),
    .Y(_3044_));
 sg13g2_a21o_1 _7271_ (.A2(_3043_),
    .A1(net1223),
    .B1(_3044_),
    .X(_3045_));
 sg13g2_nand2b_1 _7272_ (.Y(_3046_),
    .B(net622),
    .A_N(net1236));
 sg13g2_a21oi_1 _7273_ (.A1(_2909_),
    .A2(_3046_),
    .Y(_3047_),
    .B1(net1233));
 sg13g2_a21oi_1 _7274_ (.A1(net1233),
    .A2(_3045_),
    .Y(_3048_),
    .B1(_3047_));
 sg13g2_nor2_1 _7275_ (.A(net1655),
    .B(_3048_),
    .Y(_3049_));
 sg13g2_nor2_1 _7276_ (.A(_3040_),
    .B(_3041_),
    .Y(_3050_));
 sg13g2_and2_1 _7277_ (.A(_3039_),
    .B(_3050_),
    .X(_3051_));
 sg13g2_nand2_1 _7278_ (.Y(_3052_),
    .A(net1228),
    .B(net424));
 sg13g2_o21ai_1 _7279_ (.B1(_3052_),
    .Y(_3053_),
    .A1(net1228),
    .A2(_3537_));
 sg13g2_nor2b_1 _7280_ (.A(net1223),
    .B_N(net1335),
    .Y(_3054_));
 sg13g2_a21o_1 _7281_ (.A2(_3053_),
    .A1(net1223),
    .B1(_3054_),
    .X(_3055_));
 sg13g2_nand2b_1 _7282_ (.Y(_3056_),
    .B(net424),
    .A_N(net1237));
 sg13g2_a21oi_1 _7283_ (.A1(_2921_),
    .A2(_3056_),
    .Y(_3057_),
    .B1(net1234));
 sg13g2_a21oi_1 _7284_ (.A1(net1233),
    .A2(_3055_),
    .Y(_3058_),
    .B1(_3057_));
 sg13g2_a22oi_1 _7285_ (.Y(_3059_),
    .B1(_3058_),
    .B2(net1666),
    .A2(_3048_),
    .A1(net1655));
 sg13g2_nor2_1 _7286_ (.A(net1675),
    .B(_3021_),
    .Y(_3060_));
 sg13g2_nor2_1 _7287_ (.A(net1666),
    .B(_3058_),
    .Y(_3061_));
 sg13g2_nor3_1 _7288_ (.A(_3049_),
    .B(_3060_),
    .C(_3061_),
    .Y(_3062_));
 sg13g2_nand4_1 _7289_ (.B(_3051_),
    .C(_3059_),
    .A(_3023_),
    .Y(_3063_),
    .D(_3062_));
 sg13g2_nor2_1 _7290_ (.A(_3049_),
    .B(_3059_),
    .Y(_3064_));
 sg13g2_o21ai_1 _7291_ (.B1(_2986_),
    .Y(_3065_),
    .A1(_3039_),
    .A2(_3040_));
 sg13g2_a21oi_1 _7292_ (.A1(_3051_),
    .A2(_3064_),
    .Y(_3066_),
    .B1(_3065_));
 sg13g2_or2_1 _7293_ (.X(_3067_),
    .B(net1555),
    .A(net377));
 sg13g2_a21oi_1 _7294_ (.A1(_3063_),
    .A2(_3066_),
    .Y(_0063_),
    .B1(_3067_));
 sg13g2_a21oi_1 _7295_ (.A1(net1219),
    .A2(net706),
    .Y(_3068_),
    .B1(_3001_));
 sg13g2_a21oi_1 _7296_ (.A1(net1183),
    .A2(_3003_),
    .Y(_3069_),
    .B1(net1566));
 sg13g2_o21ai_1 _7297_ (.B1(_3069_),
    .Y(_3070_),
    .A1(net1183),
    .A2(_3068_));
 sg13g2_o21ai_1 _7298_ (.B1(_3070_),
    .Y(_3071_),
    .A1(net1705),
    .A2(net782));
 sg13g2_inv_1 _7299_ (.Y(_0064_),
    .A(_3071_));
 sg13g2_and2_1 _7300_ (.A(net1219),
    .B(\s0.data_out[2][1] ),
    .X(_3072_));
 sg13g2_o21ai_1 _7301_ (.B1(net1235),
    .Y(_3073_),
    .A1(_2994_),
    .A2(_3072_));
 sg13g2_nand3_1 _7302_ (.B(_2997_),
    .C(_3073_),
    .A(net1705),
    .Y(_3074_));
 sg13g2_o21ai_1 _7303_ (.B1(_3074_),
    .Y(_3075_),
    .A1(net1704),
    .A2(net771));
 sg13g2_inv_1 _7304_ (.Y(_0065_),
    .A(net772));
 sg13g2_a21oi_1 _7305_ (.A1(net1221),
    .A2(\s0.data_out[2][2] ),
    .Y(_3076_),
    .B1(_3007_));
 sg13g2_a21oi_1 _7306_ (.A1(net1184),
    .A2(_3010_),
    .Y(_3077_),
    .B1(net1571));
 sg13g2_o21ai_1 _7307_ (.B1(_3077_),
    .Y(_3078_),
    .A1(net1184),
    .A2(_3076_));
 sg13g2_o21ai_1 _7308_ (.B1(_3078_),
    .Y(_3079_),
    .A1(net1705),
    .A2(net703));
 sg13g2_inv_1 _7309_ (.Y(_0066_),
    .A(net704));
 sg13g2_nor2_1 _7310_ (.A(net1181),
    .B(_3540_),
    .Y(_3080_));
 sg13g2_o21ai_1 _7311_ (.B1(net1233),
    .Y(_3081_),
    .A1(_3017_),
    .A2(_3080_));
 sg13g2_nor2_1 _7312_ (.A(net1573),
    .B(_3020_),
    .Y(_3082_));
 sg13g2_a22oi_1 _7313_ (.Y(_0067_),
    .B1(_3081_),
    .B2(_3082_),
    .A2(_3534_),
    .A1(net1573));
 sg13g2_nor2_1 _7314_ (.A(net1181),
    .B(_3539_),
    .Y(_3083_));
 sg13g2_o21ai_1 _7315_ (.B1(net1233),
    .Y(_3084_),
    .A1(_3054_),
    .A2(_3083_));
 sg13g2_nor2_1 _7316_ (.A(net1573),
    .B(net425),
    .Y(_3085_));
 sg13g2_a22oi_1 _7317_ (.Y(_0068_),
    .B1(_3084_),
    .B2(_3085_),
    .A2(_3537_),
    .A1(net1574));
 sg13g2_and2_1 _7318_ (.A(net1223),
    .B(net622),
    .X(_3086_));
 sg13g2_o21ai_1 _7319_ (.B1(net1233),
    .Y(_3087_),
    .A1(_3044_),
    .A2(_3086_));
 sg13g2_nor2_1 _7320_ (.A(net1573),
    .B(_3047_),
    .Y(_3088_));
 sg13g2_a22oi_1 _7321_ (.Y(_0069_),
    .B1(_3087_),
    .B2(_3088_),
    .A2(_3536_),
    .A1(net1573));
 sg13g2_and2_1 _7322_ (.A(net1219),
    .B(\s0.data_out[2][6] ),
    .X(_3089_));
 sg13g2_o21ai_1 _7323_ (.B1(net1235),
    .Y(_3090_),
    .A1(_3026_),
    .A2(_3089_));
 sg13g2_nand3_1 _7324_ (.B(_3030_),
    .C(_3090_),
    .A(net1708),
    .Y(_3091_));
 sg13g2_o21ai_1 _7325_ (.B1(_3091_),
    .Y(_3092_),
    .A1(net1708),
    .A2(net816));
 sg13g2_inv_1 _7326_ (.Y(_0070_),
    .A(_3092_));
 sg13g2_nor2_1 _7327_ (.A(net1182),
    .B(_3538_),
    .Y(_3093_));
 sg13g2_o21ai_1 _7328_ (.B1(net1235),
    .Y(_3094_),
    .A1(_3034_),
    .A2(_3093_));
 sg13g2_nor2_1 _7329_ (.A(net1571),
    .B(_3037_),
    .Y(_3095_));
 sg13g2_a22oi_1 _7330_ (.Y(_0071_),
    .B1(_3094_),
    .B2(_3095_),
    .A2(_3535_),
    .A1(net1571));
 sg13g2_o21ai_1 _7331_ (.B1(net1222),
    .Y(_3096_),
    .A1(net1628),
    .A2(net1209));
 sg13g2_nor2b_1 _7332_ (.A(net1628),
    .B_N(net1216),
    .Y(_3097_));
 sg13g2_nor2_1 _7333_ (.A(_3096_),
    .B(_3097_),
    .Y(_3098_));
 sg13g2_nor2_1 _7334_ (.A(net1222),
    .B(_2984_),
    .Y(_3099_));
 sg13g2_nor2_1 _7335_ (.A(_3098_),
    .B(_3099_),
    .Y(_3100_));
 sg13g2_o21ai_1 _7336_ (.B1(_3098_),
    .Y(_3101_),
    .A1(\s0.was_valid_out[1] [0]),
    .A2(net1215));
 sg13g2_nor2_1 _7337_ (.A(net1209),
    .B(_3096_),
    .Y(_3102_));
 sg13g2_o21ai_1 _7338_ (.B1(net1180),
    .Y(_3103_),
    .A1(\s0.was_valid_out[1] [0]),
    .A2(net1226));
 sg13g2_nand2_1 _7339_ (.Y(_3104_),
    .A(_3101_),
    .B(_3103_));
 sg13g2_o21ai_1 _7340_ (.B1(net1708),
    .Y(_3105_),
    .A1(_3102_),
    .A2(_3104_));
 sg13g2_a21oi_1 _7341_ (.A1(_3359_),
    .A2(_3100_),
    .Y(_0072_),
    .B1(_3105_));
 sg13g2_nor3_1 _7342_ (.A(net1571),
    .B(_3098_),
    .C(_3099_),
    .Y(_0073_));
 sg13g2_and2_1 _7343_ (.A(net1704),
    .B(net383),
    .X(_0074_));
 sg13g2_mux2_1 _7344_ (.A0(\s0.data_out[2][2] ),
    .A1(\s0.data_out[1][2] ),
    .S(net1217),
    .X(_3106_));
 sg13g2_nor2b_1 _7345_ (.A(net1213),
    .B_N(net1340),
    .Y(_3107_));
 sg13g2_a21oi_1 _7346_ (.A1(net1213),
    .A2(_3106_),
    .Y(_3108_),
    .B1(_3107_));
 sg13g2_mux2_1 _7347_ (.A0(\s0.data_out[1][2] ),
    .A1(\s0.data_out[2][2] ),
    .S(net1226),
    .X(_3109_));
 sg13g2_nand2_1 _7348_ (.Y(_3110_),
    .A(net1181),
    .B(_3109_));
 sg13g2_o21ai_1 _7349_ (.B1(_3110_),
    .Y(_3111_),
    .A1(net1182),
    .A2(_3108_));
 sg13g2_nand2_1 _7350_ (.Y(_3112_),
    .A(net1215),
    .B(net736));
 sg13g2_mux2_1 _7351_ (.A0(\s0.data_out[2][1] ),
    .A1(\s0.data_out[1][1] ),
    .S(net1215),
    .X(_3113_));
 sg13g2_nor2b_1 _7352_ (.A(net1210),
    .B_N(net1344),
    .Y(_3114_));
 sg13g2_a21oi_1 _7353_ (.A1(net1210),
    .A2(_3113_),
    .Y(_3115_),
    .B1(_3114_));
 sg13g2_nand2b_1 _7354_ (.Y(_3116_),
    .B(net1222),
    .A_N(_3115_));
 sg13g2_o21ai_1 _7355_ (.B1(_2992_),
    .Y(_3117_),
    .A1(net1226),
    .A2(_3542_));
 sg13g2_nand2_1 _7356_ (.Y(_3118_),
    .A(net1180),
    .B(_3117_));
 sg13g2_nand3_1 _7357_ (.B(_3116_),
    .C(_3118_),
    .A(net1691),
    .Y(_3119_));
 sg13g2_mux2_1 _7358_ (.A0(\s0.data_out[2][0] ),
    .A1(\s0.data_out[1][0] ),
    .S(net1215),
    .X(_3120_));
 sg13g2_nor2b_1 _7359_ (.A(net1210),
    .B_N(net1349),
    .Y(_3121_));
 sg13g2_a21oi_1 _7360_ (.A1(net1210),
    .A2(_3120_),
    .Y(_3122_),
    .B1(_3121_));
 sg13g2_mux2_1 _7361_ (.A0(\s0.data_out[1][0] ),
    .A1(\s0.data_out[2][0] ),
    .S(net1226),
    .X(_3123_));
 sg13g2_nand2_1 _7362_ (.Y(_3124_),
    .A(net1180),
    .B(_3123_));
 sg13g2_o21ai_1 _7363_ (.B1(_3124_),
    .Y(_3125_),
    .A1(net1180),
    .A2(_3122_));
 sg13g2_and2_1 _7364_ (.A(net1559),
    .B(_3125_),
    .X(_3126_));
 sg13g2_a21oi_1 _7365_ (.A1(_3116_),
    .A2(_3118_),
    .Y(_3127_),
    .B1(net1691));
 sg13g2_a221oi_1 _7366_ (.B2(_3126_),
    .C1(_3127_),
    .B1(_3119_),
    .A1(net1560),
    .Y(_3128_),
    .A2(_3111_));
 sg13g2_or2_1 _7367_ (.X(_3129_),
    .B(_3111_),
    .A(net1560));
 sg13g2_nand2_1 _7368_ (.Y(_3130_),
    .A(net1217),
    .B(\s0.data_out[1][3] ));
 sg13g2_o21ai_1 _7369_ (.B1(_3130_),
    .Y(_3131_),
    .A1(net1217),
    .A2(_3540_));
 sg13g2_nor2_1 _7370_ (.A(net1213),
    .B(net1160),
    .Y(_3132_));
 sg13g2_a21o_1 _7371_ (.A2(_3131_),
    .A1(net1213),
    .B1(_3132_),
    .X(_3133_));
 sg13g2_nand2b_1 _7372_ (.Y(_3134_),
    .B(net602),
    .A_N(net1228));
 sg13g2_a21oi_1 _7373_ (.A1(_3015_),
    .A2(_3134_),
    .Y(_3135_),
    .B1(net1223));
 sg13g2_a21oi_1 _7374_ (.A1(net1224),
    .A2(_3133_),
    .Y(_3136_),
    .B1(_3135_));
 sg13g2_nand2_1 _7375_ (.Y(_3137_),
    .A(net1674),
    .B(_3136_));
 sg13g2_nand3b_1 _7376_ (.B(_3129_),
    .C(_3137_),
    .Y(_3138_),
    .A_N(_3128_));
 sg13g2_mux2_1 _7377_ (.A0(\s0.data_out[2][6] ),
    .A1(\s0.data_out[1][6] ),
    .S(net1215),
    .X(_3139_));
 sg13g2_nor2b_1 _7378_ (.A(net1209),
    .B_N(net1325),
    .Y(_3140_));
 sg13g2_a21o_1 _7379_ (.A2(_3139_),
    .A1(net1209),
    .B1(_3140_),
    .X(_3141_));
 sg13g2_nand2b_1 _7380_ (.Y(_3142_),
    .B(\s0.data_out[1][6] ),
    .A_N(net1226));
 sg13g2_a21oi_1 _7381_ (.A1(_3024_),
    .A2(_3142_),
    .Y(_3143_),
    .B1(net1222));
 sg13g2_a21oi_1 _7382_ (.A1(net1225),
    .A2(_3141_),
    .Y(_3144_),
    .B1(_3143_));
 sg13g2_mux2_1 _7383_ (.A0(\s0.data_out[2][7] ),
    .A1(\s0.data_out[1][7] ),
    .S(net1215),
    .X(_3145_));
 sg13g2_nor2b_1 _7384_ (.A(net1211),
    .B_N(net1320),
    .Y(_3146_));
 sg13g2_a21o_1 _7385_ (.A2(_3145_),
    .A1(net1211),
    .B1(_3146_),
    .X(_3147_));
 sg13g2_nand2b_1 _7386_ (.Y(_3148_),
    .B(\s0.data_out[1][7] ),
    .A_N(net1227));
 sg13g2_a21oi_1 _7387_ (.A1(_3032_),
    .A2(_3148_),
    .Y(_3149_),
    .B1(net1222));
 sg13g2_a21oi_1 _7388_ (.A1(net1222),
    .A2(_3147_),
    .Y(_3150_),
    .B1(_3149_));
 sg13g2_a22oi_1 _7389_ (.Y(_3151_),
    .B1(_3150_),
    .B2(net1636),
    .A2(_3144_),
    .A1(net1647));
 sg13g2_nor2_1 _7390_ (.A(net1647),
    .B(_3144_),
    .Y(_3152_));
 sg13g2_nor2_1 _7391_ (.A(net1635),
    .B(_3150_),
    .Y(_3153_));
 sg13g2_or2_1 _7392_ (.X(_3154_),
    .B(_3150_),
    .A(net1635));
 sg13g2_mux2_1 _7393_ (.A0(\s0.data_out[2][5] ),
    .A1(\s0.data_out[1][5] ),
    .S(net1217),
    .X(_3155_));
 sg13g2_nor2b_1 _7394_ (.A(net1213),
    .B_N(net1331),
    .Y(_3156_));
 sg13g2_a21oi_1 _7395_ (.A1(net1214),
    .A2(_3155_),
    .Y(_3157_),
    .B1(_3156_));
 sg13g2_o21ai_1 _7396_ (.B1(_3042_),
    .Y(_3158_),
    .A1(net1229),
    .A2(_3541_));
 sg13g2_nand2_1 _7397_ (.Y(_3159_),
    .A(net1181),
    .B(_3158_));
 sg13g2_o21ai_1 _7398_ (.B1(_3159_),
    .Y(_3160_),
    .A1(net1181),
    .A2(_3157_));
 sg13g2_and2_1 _7399_ (.A(_3403_),
    .B(_3160_),
    .X(_3161_));
 sg13g2_nand3b_1 _7400_ (.B(_3154_),
    .C(_3151_),
    .Y(_3162_),
    .A_N(_3152_));
 sg13g2_nor2_1 _7401_ (.A(_3161_),
    .B(_3162_),
    .Y(_3163_));
 sg13g2_mux2_1 _7402_ (.A0(\s0.data_out[2][4] ),
    .A1(\s0.data_out[1][4] ),
    .S(net1217),
    .X(_3164_));
 sg13g2_nor2b_1 _7403_ (.A(net1214),
    .B_N(net1336),
    .Y(_3165_));
 sg13g2_a21o_1 _7404_ (.A2(_3164_),
    .A1(net1213),
    .B1(_3165_),
    .X(_3166_));
 sg13g2_nand2b_1 _7405_ (.Y(_3167_),
    .B(net566),
    .A_N(net1228));
 sg13g2_a21oi_1 _7406_ (.A1(_3052_),
    .A2(_3167_),
    .Y(_3168_),
    .B1(net1224));
 sg13g2_a21oi_1 _7407_ (.A1(net1224),
    .A2(_3166_),
    .Y(_3169_),
    .B1(_3168_));
 sg13g2_nand2_1 _7408_ (.Y(_3170_),
    .A(net1666),
    .B(_3169_));
 sg13g2_o21ai_1 _7409_ (.B1(_3170_),
    .Y(_3171_),
    .A1(_3403_),
    .A2(_3160_));
 sg13g2_or2_1 _7410_ (.X(_3172_),
    .B(_3169_),
    .A(net1666));
 sg13g2_o21ai_1 _7411_ (.B1(_3172_),
    .Y(_3173_),
    .A1(net1674),
    .A2(_3136_));
 sg13g2_nor4_1 _7412_ (.A(_3161_),
    .B(_3162_),
    .C(_3171_),
    .D(_3173_),
    .Y(_3174_));
 sg13g2_o21ai_1 _7413_ (.B1(_3100_),
    .Y(_3175_),
    .A1(_3151_),
    .A2(_3153_));
 sg13g2_a221oi_1 _7414_ (.B2(_3138_),
    .C1(_3175_),
    .B1(_3174_),
    .A1(_3163_),
    .Y(_3176_),
    .A2(_3171_));
 sg13g2_nor3_1 _7415_ (.A(net372),
    .B(net1555),
    .C(_3176_),
    .Y(_0075_));
 sg13g2_a21oi_1 _7416_ (.A1(net1210),
    .A2(\s0.data_out[1][0] ),
    .Y(_3177_),
    .B1(_3121_));
 sg13g2_a21oi_1 _7417_ (.A1(net1180),
    .A2(_3123_),
    .Y(_3178_),
    .B1(net1571));
 sg13g2_o21ai_1 _7418_ (.B1(_3178_),
    .Y(_3179_),
    .A1(net1180),
    .A2(_3177_));
 sg13g2_o21ai_1 _7419_ (.B1(_3179_),
    .Y(_3180_),
    .A1(net1708),
    .A2(net706));
 sg13g2_inv_1 _7420_ (.Y(_0076_),
    .A(net707));
 sg13g2_a21oi_1 _7421_ (.A1(net1210),
    .A2(\s0.data_out[1][1] ),
    .Y(_3181_),
    .B1(_3114_));
 sg13g2_a21oi_1 _7422_ (.A1(net1180),
    .A2(_3117_),
    .Y(_3182_),
    .B1(net1571));
 sg13g2_o21ai_1 _7423_ (.B1(_3182_),
    .Y(_3183_),
    .A1(net1180),
    .A2(_3181_));
 sg13g2_o21ai_1 _7424_ (.B1(_3183_),
    .Y(_3184_),
    .A1(net1708),
    .A2(net698));
 sg13g2_inv_1 _7425_ (.Y(_0077_),
    .A(net699));
 sg13g2_a21oi_1 _7426_ (.A1(net1213),
    .A2(net762),
    .Y(_3185_),
    .B1(_3107_));
 sg13g2_a21oi_1 _7427_ (.A1(net1181),
    .A2(_3109_),
    .Y(_3186_),
    .B1(net1572));
 sg13g2_o21ai_1 _7428_ (.B1(_3186_),
    .Y(_3187_),
    .A1(net1181),
    .A2(_3185_));
 sg13g2_o21ai_1 _7429_ (.B1(_3187_),
    .Y(_3188_),
    .A1(net1711),
    .A2(net774));
 sg13g2_inv_1 _7430_ (.Y(_0078_),
    .A(_3188_));
 sg13g2_and2_1 _7431_ (.A(net1213),
    .B(net602),
    .X(_3189_));
 sg13g2_o21ai_1 _7432_ (.B1(net1223),
    .Y(_3190_),
    .A1(_3132_),
    .A2(_3189_));
 sg13g2_nor2_1 _7433_ (.A(net1573),
    .B(_3135_),
    .Y(_3191_));
 sg13g2_a22oi_1 _7434_ (.Y(_0079_),
    .B1(_3190_),
    .B2(_3191_),
    .A2(_3540_),
    .A1(net1573));
 sg13g2_and2_1 _7435_ (.A(net1214),
    .B(net566),
    .X(_3192_));
 sg13g2_o21ai_1 _7436_ (.B1(net1224),
    .Y(_3193_),
    .A1(_3165_),
    .A2(_3192_));
 sg13g2_nor2_1 _7437_ (.A(net1575),
    .B(_3168_),
    .Y(_3194_));
 sg13g2_a22oi_1 _7438_ (.Y(_0080_),
    .B1(net567),
    .B2(_3194_),
    .A2(_3539_),
    .A1(net1575));
 sg13g2_a21oi_1 _7439_ (.A1(net1214),
    .A2(\s0.data_out[1][5] ),
    .Y(_3195_),
    .B1(_3156_));
 sg13g2_a21oi_1 _7440_ (.A1(net1182),
    .A2(_3158_),
    .Y(_3196_),
    .B1(net1573));
 sg13g2_o21ai_1 _7441_ (.B1(_3196_),
    .Y(_3197_),
    .A1(net1181),
    .A2(_3195_));
 sg13g2_o21ai_1 _7442_ (.B1(_3197_),
    .Y(_3198_),
    .A1(net1713),
    .A2(net622));
 sg13g2_inv_1 _7443_ (.Y(_0081_),
    .A(net623));
 sg13g2_and2_1 _7444_ (.A(net1209),
    .B(\s0.data_out[1][6] ),
    .X(_3199_));
 sg13g2_o21ai_1 _7445_ (.B1(net1225),
    .Y(_3200_),
    .A1(_3140_),
    .A2(_3199_));
 sg13g2_nand3b_1 _7446_ (.B(_3200_),
    .C(net1708),
    .Y(_3201_),
    .A_N(_3143_));
 sg13g2_o21ai_1 _7447_ (.B1(_3201_),
    .Y(_3202_),
    .A1(net1708),
    .A2(net793));
 sg13g2_inv_1 _7448_ (.Y(_0082_),
    .A(net794));
 sg13g2_and2_1 _7449_ (.A(net1211),
    .B(\s0.data_out[1][7] ),
    .X(_3203_));
 sg13g2_o21ai_1 _7450_ (.B1(net1222),
    .Y(_3204_),
    .A1(_3146_),
    .A2(_3203_));
 sg13g2_nor2_1 _7451_ (.A(net1571),
    .B(_3149_),
    .Y(_3205_));
 sg13g2_a22oi_1 _7452_ (.Y(_0083_),
    .B1(_3204_),
    .B2(_3205_),
    .A2(_3538_),
    .A1(net1571));
 sg13g2_o21ai_1 _7453_ (.B1(net1212),
    .Y(_3206_),
    .A1(net1628),
    .A2(net1201));
 sg13g2_a21oi_1 _7454_ (.A1(net1621),
    .A2(net1206),
    .Y(_3207_),
    .B1(_3206_));
 sg13g2_inv_1 _7455_ (.Y(_3208_),
    .A(_3207_));
 sg13g2_o21ai_1 _7456_ (.B1(_3208_),
    .Y(_3209_),
    .A1(net1212),
    .A2(_3097_));
 sg13g2_or2_1 _7457_ (.X(_3210_),
    .B(net1206),
    .A(net504));
 sg13g2_o21ai_1 _7458_ (.B1(net1195),
    .Y(_3211_),
    .A1(net504),
    .A2(net1215));
 sg13g2_o21ai_1 _7459_ (.B1(_3211_),
    .Y(_3212_),
    .A1(net1201),
    .A2(_3206_));
 sg13g2_a21oi_1 _7460_ (.A1(_3207_),
    .A2(_3210_),
    .Y(_3213_),
    .B1(_3212_));
 sg13g2_o21ai_1 _7461_ (.B1(net1709),
    .Y(_3214_),
    .A1(net620),
    .A2(_3209_));
 sg13g2_nor2_1 _7462_ (.A(_3213_),
    .B(_3214_),
    .Y(_0084_));
 sg13g2_nor2_1 _7463_ (.A(net1572),
    .B(_3209_),
    .Y(_0085_));
 sg13g2_and2_1 _7464_ (.A(net1731),
    .B(net370),
    .X(_0086_));
 sg13g2_mux2_1 _7465_ (.A0(\s0.data_out[0][2] ),
    .A1(\s0.data_out[1][2] ),
    .S(net1217),
    .X(_3215_));
 sg13g2_mux2_1 _7466_ (.A0(\s0.data_out[1][2] ),
    .A1(\s0.data_out[0][2] ),
    .S(net1207),
    .X(_3216_));
 sg13g2_nor2b_1 _7467_ (.A(net1203),
    .B_N(net1340),
    .Y(_3217_));
 sg13g2_a21oi_1 _7468_ (.A1(net1204),
    .A2(_3216_),
    .Y(_3218_),
    .B1(_3217_));
 sg13g2_nor2_1 _7469_ (.A(net1194),
    .B(_3218_),
    .Y(_3219_));
 sg13g2_a21oi_1 _7470_ (.A1(net1194),
    .A2(_3215_),
    .Y(_3220_),
    .B1(_3219_));
 sg13g2_nand2b_1 _7471_ (.Y(_3221_),
    .B(net431),
    .A_N(net1215));
 sg13g2_a21oi_1 _7472_ (.A1(_3112_),
    .A2(_3221_),
    .Y(_3222_),
    .B1(net1209));
 sg13g2_mux2_1 _7473_ (.A0(\s0.data_out[1][1] ),
    .A1(\s0.data_out[0][1] ),
    .S(net1206),
    .X(_3223_));
 sg13g2_nor2b_1 _7474_ (.A(net1200),
    .B_N(net1344),
    .Y(_3224_));
 sg13g2_a21o_1 _7475_ (.A2(_3223_),
    .A1(net1200),
    .B1(_3224_),
    .X(_3225_));
 sg13g2_a21oi_1 _7476_ (.A1(net1210),
    .A2(_3225_),
    .Y(_3226_),
    .B1(_3222_));
 sg13g2_mux2_1 _7477_ (.A0(\s0.data_out[0][0] ),
    .A1(\s0.data_out[1][0] ),
    .S(net1216),
    .X(_3227_));
 sg13g2_nand2_1 _7478_ (.Y(_3228_),
    .A(net1195),
    .B(_3227_));
 sg13g2_mux2_1 _7479_ (.A0(\s0.data_out[1][0] ),
    .A1(\s0.data_out[0][0] ),
    .S(net1206),
    .X(_3229_));
 sg13g2_nor2b_1 _7480_ (.A(net1200),
    .B_N(net1348),
    .Y(_3230_));
 sg13g2_a21oi_1 _7481_ (.A1(net1200),
    .A2(_3229_),
    .Y(_3231_),
    .B1(_3230_));
 sg13g2_nand2b_1 _7482_ (.Y(_3232_),
    .B(net1209),
    .A_N(_3231_));
 sg13g2_or2_1 _7483_ (.X(_3233_),
    .B(_3226_),
    .A(net1691));
 sg13g2_a221oi_1 _7484_ (.B2(_3232_),
    .C1(net1700),
    .B1(_3228_),
    .A1(net1691),
    .Y(_3234_),
    .A2(_3226_));
 sg13g2_o21ai_1 _7485_ (.B1(_3233_),
    .Y(_3235_),
    .A1(net1684),
    .A2(_3220_));
 sg13g2_o21ai_1 _7486_ (.B1(_3130_),
    .Y(_3236_),
    .A1(net1217),
    .A2(_3543_));
 sg13g2_mux2_1 _7487_ (.A0(\s0.data_out[1][3] ),
    .A1(\s0.data_out[0][3] ),
    .S(net1208),
    .X(_3237_));
 sg13g2_nor2b_1 _7488_ (.A(net1204),
    .B_N(net1339),
    .Y(_3238_));
 sg13g2_a21oi_1 _7489_ (.A1(net1204),
    .A2(_3237_),
    .Y(_3239_),
    .B1(_3238_));
 sg13g2_nor2_1 _7490_ (.A(net1193),
    .B(_3239_),
    .Y(_3240_));
 sg13g2_a21oi_1 _7491_ (.A1(net1193),
    .A2(_3236_),
    .Y(_3241_),
    .B1(_3240_));
 sg13g2_a22oi_1 _7492_ (.Y(_3242_),
    .B1(_3241_),
    .B2(net1674),
    .A2(_3220_),
    .A1(net1684));
 sg13g2_o21ai_1 _7493_ (.B1(_3242_),
    .Y(_3243_),
    .A1(_3234_),
    .A2(_3235_));
 sg13g2_mux2_1 _7494_ (.A0(\s0.data_out[0][7] ),
    .A1(\s0.data_out[1][7] ),
    .S(net1216),
    .X(_3244_));
 sg13g2_mux2_1 _7495_ (.A0(\s0.data_out[1][7] ),
    .A1(\s0.data_out[0][7] ),
    .S(net1206),
    .X(_3245_));
 sg13g2_nor2b_1 _7496_ (.A(net1202),
    .B_N(net1321),
    .Y(_3246_));
 sg13g2_a21oi_1 _7497_ (.A1(net1202),
    .A2(_3245_),
    .Y(_3247_),
    .B1(_3246_));
 sg13g2_nor2_1 _7498_ (.A(net1212),
    .B(_3244_),
    .Y(_3248_));
 sg13g2_a21o_1 _7499_ (.A2(_3247_),
    .A1(net1214),
    .B1(_3248_),
    .X(_3249_));
 sg13g2_mux2_1 _7500_ (.A0(\s0.data_out[0][6] ),
    .A1(\s0.data_out[1][6] ),
    .S(net1216),
    .X(_3250_));
 sg13g2_mux2_1 _7501_ (.A0(\s0.data_out[1][6] ),
    .A1(\s0.data_out[0][6] ),
    .S(net1207),
    .X(_3251_));
 sg13g2_nor2b_1 _7502_ (.A(net1201),
    .B_N(net1326),
    .Y(_3252_));
 sg13g2_a21oi_1 _7503_ (.A1(net1201),
    .A2(_3251_),
    .Y(_3253_),
    .B1(_3252_));
 sg13g2_nor2_1 _7504_ (.A(net1212),
    .B(_3250_),
    .Y(_3254_));
 sg13g2_a21o_1 _7505_ (.A2(_3253_),
    .A1(net1212),
    .B1(_3254_),
    .X(_3255_));
 sg13g2_a22oi_1 _7506_ (.Y(_3256_),
    .B1(_3255_),
    .B2(net1647),
    .A2(_3249_),
    .A1(net1635));
 sg13g2_or2_1 _7507_ (.X(_3257_),
    .B(_3249_),
    .A(net1635));
 sg13g2_or2_1 _7508_ (.X(_3258_),
    .B(_3255_),
    .A(net1647));
 sg13g2_nand3_1 _7509_ (.B(_3257_),
    .C(_3258_),
    .A(_3256_),
    .Y(_3259_));
 sg13g2_mux2_1 _7510_ (.A0(\s0.data_out[0][5] ),
    .A1(\s0.data_out[1][5] ),
    .S(net1218),
    .X(_3260_));
 sg13g2_nand2_1 _7511_ (.Y(_3261_),
    .A(net1194),
    .B(_3260_));
 sg13g2_mux2_1 _7512_ (.A0(\s0.data_out[1][5] ),
    .A1(\s0.data_out[0][5] ),
    .S(net1207),
    .X(_3262_));
 sg13g2_nor2b_1 _7513_ (.A(net1205),
    .B_N(net1330),
    .Y(_3263_));
 sg13g2_a21oi_1 _7514_ (.A1(net1205),
    .A2(_3262_),
    .Y(_3264_),
    .B1(_3263_));
 sg13g2_nand2b_1 _7515_ (.Y(_3265_),
    .B(net1214),
    .A_N(_3264_));
 sg13g2_nand3_1 _7516_ (.B(_3261_),
    .C(_3265_),
    .A(net1656),
    .Y(_3266_));
 sg13g2_inv_1 _7517_ (.Y(_3267_),
    .A(_3266_));
 sg13g2_mux2_1 _7518_ (.A0(\s0.data_out[0][4] ),
    .A1(\s0.data_out[1][4] ),
    .S(net1217),
    .X(_3268_));
 sg13g2_nand2_1 _7519_ (.Y(_3269_),
    .A(net1193),
    .B(_3268_));
 sg13g2_mux2_1 _7520_ (.A0(\s0.data_out[1][4] ),
    .A1(\s0.data_out[0][4] ),
    .S(net1207),
    .X(_3270_));
 sg13g2_nor2b_1 _7521_ (.A(net1204),
    .B_N(net1335),
    .Y(_3271_));
 sg13g2_a21oi_1 _7522_ (.A1(net1204),
    .A2(_3270_),
    .Y(_3272_),
    .B1(_3271_));
 sg13g2_nand2b_1 _7523_ (.Y(_3273_),
    .B(net1214),
    .A_N(_3272_));
 sg13g2_a21oi_1 _7524_ (.A1(_3269_),
    .A2(_3273_),
    .Y(_3274_),
    .B1(net1665));
 sg13g2_nand3_1 _7525_ (.B(_3269_),
    .C(_3273_),
    .A(net1665),
    .Y(_3275_));
 sg13g2_o21ai_1 _7526_ (.B1(_3275_),
    .Y(_3276_),
    .A1(net1674),
    .A2(_3241_));
 sg13g2_a21oi_1 _7527_ (.A1(_3261_),
    .A2(_3265_),
    .Y(_3277_),
    .B1(net1656));
 sg13g2_nor4_1 _7528_ (.A(_3267_),
    .B(_3274_),
    .C(_3276_),
    .D(_3277_),
    .Y(_3278_));
 sg13g2_nand3b_1 _7529_ (.B(_3278_),
    .C(_3243_),
    .Y(_3279_),
    .A_N(_3259_));
 sg13g2_o21ai_1 _7530_ (.B1(_3266_),
    .Y(_3280_),
    .A1(_3275_),
    .A2(_3277_));
 sg13g2_nor2b_1 _7531_ (.A(_3259_),
    .B_N(_3280_),
    .Y(_3281_));
 sg13g2_nor2b_1 _7532_ (.A(_3256_),
    .B_N(_3257_),
    .Y(_3282_));
 sg13g2_nor3_1 _7533_ (.A(_3209_),
    .B(_3281_),
    .C(_3282_),
    .Y(_3283_));
 sg13g2_or2_1 _7534_ (.X(_3284_),
    .B(net1555),
    .A(net395));
 sg13g2_a21oi_1 _7535_ (.A1(_3279_),
    .A2(_3283_),
    .Y(_0087_),
    .B1(_3284_));
 sg13g2_and2_1 _7536_ (.A(net1200),
    .B(\s0.data_out[0][0] ),
    .X(_3285_));
 sg13g2_o21ai_1 _7537_ (.B1(net1212),
    .Y(_3286_),
    .A1(_3230_),
    .A2(_3285_));
 sg13g2_nand3_1 _7538_ (.B(_3228_),
    .C(_3286_),
    .A(net1709),
    .Y(_3287_));
 sg13g2_o21ai_1 _7539_ (.B1(_3287_),
    .Y(_3288_),
    .A1(net1709),
    .A2(net791));
 sg13g2_inv_1 _7540_ (.Y(_0088_),
    .A(net792));
 sg13g2_and2_1 _7541_ (.A(net1200),
    .B(net431),
    .X(_3289_));
 sg13g2_o21ai_1 _7542_ (.B1(net1209),
    .Y(_3290_),
    .A1(_3224_),
    .A2(_3289_));
 sg13g2_nor2_1 _7543_ (.A(net1572),
    .B(_3222_),
    .Y(_3291_));
 sg13g2_a22oi_1 _7544_ (.Y(_0089_),
    .B1(_3290_),
    .B2(_3291_),
    .A2(_3542_),
    .A1(net1572));
 sg13g2_a21oi_1 _7545_ (.A1(net1203),
    .A2(net469),
    .Y(_3292_),
    .B1(_3217_));
 sg13g2_a21oi_1 _7546_ (.A1(net1194),
    .A2(_3215_),
    .Y(_3293_),
    .B1(net1576));
 sg13g2_o21ai_1 _7547_ (.B1(_3293_),
    .Y(_3294_),
    .A1(net1195),
    .A2(_3292_));
 sg13g2_o21ai_1 _7548_ (.B1(_3294_),
    .Y(_3295_),
    .A1(net1710),
    .A2(net762));
 sg13g2_inv_1 _7549_ (.Y(_0090_),
    .A(net763));
 sg13g2_a21oi_1 _7550_ (.A1(net1204),
    .A2(net441),
    .Y(_3296_),
    .B1(_3238_));
 sg13g2_a21oi_1 _7551_ (.A1(net1193),
    .A2(_3236_),
    .Y(_3297_),
    .B1(net1575));
 sg13g2_o21ai_1 _7552_ (.B1(_3297_),
    .Y(_3298_),
    .A1(net1193),
    .A2(_3296_));
 sg13g2_o21ai_1 _7553_ (.B1(_3298_),
    .Y(_3299_),
    .A1(net1712),
    .A2(net602));
 sg13g2_inv_1 _7554_ (.Y(_0091_),
    .A(net603));
 sg13g2_a21oi_1 _7555_ (.A1(net1205),
    .A2(net443),
    .Y(_3300_),
    .B1(_3271_));
 sg13g2_a21oi_1 _7556_ (.A1(net1193),
    .A2(_3268_),
    .Y(_3301_),
    .B1(net1575));
 sg13g2_o21ai_1 _7557_ (.B1(_3301_),
    .Y(_3302_),
    .A1(net1193),
    .A2(_3300_));
 sg13g2_o21ai_1 _7558_ (.B1(_3302_),
    .Y(_3303_),
    .A1(net1712),
    .A2(net566));
 sg13g2_inv_1 _7559_ (.Y(_0092_),
    .A(_3303_));
 sg13g2_a21oi_1 _7560_ (.A1(net1205),
    .A2(net435),
    .Y(_3304_),
    .B1(_3263_));
 sg13g2_a21oi_1 _7561_ (.A1(net1193),
    .A2(_3260_),
    .Y(_3305_),
    .B1(net1575));
 sg13g2_o21ai_1 _7562_ (.B1(_3305_),
    .Y(_3306_),
    .A1(net1194),
    .A2(_3304_));
 sg13g2_o21ai_1 _7563_ (.B1(_3306_),
    .Y(_3307_),
    .A1(net1713),
    .A2(net745));
 sg13g2_inv_1 _7564_ (.Y(_0093_),
    .A(_3307_));
 sg13g2_a21oi_1 _7565_ (.A1(net1201),
    .A2(net494),
    .Y(_3308_),
    .B1(_3252_));
 sg13g2_a21oi_1 _7566_ (.A1(net1195),
    .A2(_3250_),
    .Y(_3309_),
    .B1(net1572));
 sg13g2_o21ai_1 _7567_ (.B1(_3309_),
    .Y(_3310_),
    .A1(net1195),
    .A2(_3308_));
 sg13g2_o21ai_1 _7568_ (.B1(_3310_),
    .Y(_3311_),
    .A1(net1710),
    .A2(net822));
 sg13g2_inv_1 _7569_ (.Y(_0094_),
    .A(_3311_));
 sg13g2_a21oi_1 _7570_ (.A1(net1202),
    .A2(net451),
    .Y(_3312_),
    .B1(_3246_));
 sg13g2_a21oi_1 _7571_ (.A1(net1195),
    .A2(_3244_),
    .Y(_3313_),
    .B1(net1576));
 sg13g2_o21ai_1 _7572_ (.B1(_3313_),
    .Y(_3314_),
    .A1(net1195),
    .A2(_3312_));
 sg13g2_o21ai_1 _7573_ (.B1(_3314_),
    .Y(_3315_),
    .A1(net1710),
    .A2(net801));
 sg13g2_inv_1 _7574_ (.Y(_0095_),
    .A(_3315_));
 sg13g2_a21oi_1 _7575_ (.A1(net504),
    .A2(_3393_),
    .Y(_3316_),
    .B1(net1627));
 sg13g2_o21ai_1 _7576_ (.B1(net1710),
    .Y(_3317_),
    .A1(net1206),
    .A2(net1201));
 sg13g2_nor2_1 _7577_ (.A(_3316_),
    .B(_3317_),
    .Y(_0096_));
 sg13g2_nor2_1 _7578_ (.A(net1627),
    .B(_3317_),
    .Y(_0097_));
 sg13g2_and2_1 _7579_ (.A(net1727),
    .B(net388),
    .X(_0098_));
 sg13g2_a21oi_1 _7580_ (.A1(net1207),
    .A2(net494),
    .Y(_3318_),
    .B1(net1201));
 sg13g2_a21oi_1 _7581_ (.A1(net1201),
    .A2(_3401_),
    .Y(_3319_),
    .B1(_3318_));
 sg13g2_a21o_1 _7582_ (.A2(net451),
    .A1(net1207),
    .B1(net1202),
    .X(_3320_));
 sg13g2_o21ai_1 _7583_ (.B1(_3320_),
    .Y(_3321_),
    .A1(_3393_),
    .A2(net1321));
 sg13g2_nor2_1 _7584_ (.A(net1635),
    .B(_3321_),
    .Y(_3322_));
 sg13g2_a21oi_1 _7585_ (.A1(_3402_),
    .A2(_3319_),
    .Y(_3323_),
    .B1(_3322_));
 sg13g2_nor2_1 _7586_ (.A(_3402_),
    .B(_3319_),
    .Y(_3324_));
 sg13g2_a21o_1 _7587_ (.A2(net435),
    .A1(net1207),
    .B1(net1205),
    .X(_3325_));
 sg13g2_o21ai_1 _7588_ (.B1(_3325_),
    .Y(_3326_),
    .A1(_3393_),
    .A2(net1330));
 sg13g2_nor2_1 _7589_ (.A(net1656),
    .B(_3326_),
    .Y(_3327_));
 sg13g2_a21o_1 _7590_ (.A2(net431),
    .A1(net1206),
    .B1(net1200),
    .X(_3328_));
 sg13g2_o21ai_1 _7591_ (.B1(_3328_),
    .Y(_3329_),
    .A1(_3393_),
    .A2(net1345));
 sg13g2_nand2_1 _7592_ (.Y(_3330_),
    .A(net1200),
    .B(net1348));
 sg13g2_nand3_1 _7593_ (.B(_3393_),
    .C(net604),
    .A(net1206),
    .Y(_3331_));
 sg13g2_a221oi_1 _7594_ (.B2(_3331_),
    .C1(net1700),
    .B1(_3330_),
    .A1(net1691),
    .Y(_3332_),
    .A2(_3329_));
 sg13g2_nor2_1 _7595_ (.A(net1691),
    .B(_3329_),
    .Y(_3333_));
 sg13g2_a21o_1 _7596_ (.A2(net469),
    .A1(net1208),
    .B1(net1203),
    .X(_3334_));
 sg13g2_o21ai_1 _7597_ (.B1(_3334_),
    .Y(_3335_),
    .A1(_3393_),
    .A2(net1341));
 sg13g2_nor2_1 _7598_ (.A(net1685),
    .B(_3335_),
    .Y(_3336_));
 sg13g2_or3_1 _7599_ (.A(_3332_),
    .B(_3333_),
    .C(_3336_),
    .X(_3337_));
 sg13g2_a21oi_1 _7600_ (.A1(net1208),
    .A2(net441),
    .Y(_3338_),
    .B1(net1204));
 sg13g2_a21oi_1 _7601_ (.A1(net1204),
    .A2(net1160),
    .Y(_3339_),
    .B1(_3338_));
 sg13g2_inv_1 _7602_ (.Y(_3340_),
    .A(_3339_));
 sg13g2_a22oi_1 _7603_ (.Y(_3341_),
    .B1(_3340_),
    .B2(net1674),
    .A2(_3335_),
    .A1(net1684));
 sg13g2_a21o_1 _7604_ (.A2(net443),
    .A1(net1208),
    .B1(net1205),
    .X(_3342_));
 sg13g2_o21ai_1 _7605_ (.B1(_3342_),
    .Y(_3343_),
    .A1(_3393_),
    .A2(net1335));
 sg13g2_nand2b_1 _7606_ (.Y(_3344_),
    .B(_3406_),
    .A_N(_3343_));
 sg13g2_o21ai_1 _7607_ (.B1(_3344_),
    .Y(_3345_),
    .A1(net1674),
    .A2(_3340_));
 sg13g2_a21o_1 _7608_ (.A2(_3341_),
    .A1(_3337_),
    .B1(_3345_),
    .X(_3346_));
 sg13g2_a22oi_1 _7609_ (.Y(_3347_),
    .B1(_3343_),
    .B2(net1666),
    .A2(_3326_),
    .A1(net1656));
 sg13g2_a21oi_1 _7610_ (.A1(_3346_),
    .A2(_3347_),
    .Y(_3348_),
    .B1(_3327_));
 sg13g2_o21ai_1 _7611_ (.B1(_3323_),
    .Y(_3349_),
    .A1(_3324_),
    .A2(_3348_));
 sg13g2_a21oi_1 _7612_ (.A1(net1635),
    .A2(_3321_),
    .Y(_3350_),
    .B1(net1628));
 sg13g2_or2_1 _7613_ (.X(_3351_),
    .B(net1555),
    .A(net384));
 sg13g2_a21oi_1 _7614_ (.A1(_3349_),
    .A2(_3350_),
    .Y(_0099_),
    .B1(_3351_));
 sg13g2_a21oi_1 _7615_ (.A1(_3330_),
    .A2(_3331_),
    .Y(_3352_),
    .B1(net1572));
 sg13g2_a21o_1 _7616_ (.A2(net604),
    .A1(net1572),
    .B1(_3352_),
    .X(_0100_));
 sg13g2_nor2_1 _7617_ (.A(net1709),
    .B(net431),
    .Y(_3353_));
 sg13g2_a21oi_1 _7618_ (.A1(net1709),
    .A2(_3329_),
    .Y(_0101_),
    .B1(_3353_));
 sg13g2_nor2_1 _7619_ (.A(net1710),
    .B(net469),
    .Y(_3354_));
 sg13g2_a21oi_1 _7620_ (.A1(net1710),
    .A2(_3335_),
    .Y(_0102_),
    .B1(_3354_));
 sg13g2_nor2_1 _7621_ (.A(net1712),
    .B(net441),
    .Y(_3355_));
 sg13g2_a21oi_1 _7622_ (.A1(net1712),
    .A2(_3340_),
    .Y(_0103_),
    .B1(_3355_));
 sg13g2_nor2_1 _7623_ (.A(net1712),
    .B(net443),
    .Y(_3356_));
 sg13g2_a21oi_1 _7624_ (.A1(net1712),
    .A2(_3343_),
    .Y(_0104_),
    .B1(_3356_));
 sg13g2_nor2_1 _7625_ (.A(net1712),
    .B(net435),
    .Y(_3357_));
 sg13g2_a21oi_1 _7626_ (.A1(net1712),
    .A2(_3326_),
    .Y(_0105_),
    .B1(_3357_));
 sg13g2_mux2_1 _7627_ (.A0(net494),
    .A1(_3319_),
    .S(net1709),
    .X(_0106_));
 sg13g2_nor2_1 _7628_ (.A(net1710),
    .B(net451),
    .Y(_3358_));
 sg13g2_a21oi_1 _7629_ (.A1(net1711),
    .A2(_3321_),
    .Y(_0107_),
    .B1(_3358_));
 sg13g2_dfrbpq_1 _7630_ (.RESET_B(net204),
    .D(_0108_),
    .Q(\s0.module0.bubble ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _7631_ (.RESET_B(net56),
    .D(net770),
    .Q(\s0.was_valid_out[27] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _7632_ (.RESET_B(net54),
    .D(_0110_),
    .Q(\s0.valid_out[27] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _7633_ (.RESET_B(net53),
    .D(_0111_),
    .Q(\s0.genblk1[26].modules.bubble ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _7634_ (.RESET_B(net52),
    .D(_0112_),
    .Q(\s0.shift_out[27] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _7635_ (.RESET_B(net51),
    .D(net525),
    .Q(\s0.data_out[27][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _7636_ (.RESET_B(net50),
    .D(net601),
    .Q(\s0.data_out[27][1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _7637_ (.RESET_B(net49),
    .D(net508),
    .Q(\s0.data_out[27][2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _7638_ (.RESET_B(net48),
    .D(net457),
    .Q(\s0.data_out[27][3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _7639_ (.RESET_B(net47),
    .D(net464),
    .Q(\s0.data_out[27][4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _7640_ (.RESET_B(net46),
    .D(net468),
    .Q(\s0.data_out[27][5] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _7641_ (.RESET_B(net45),
    .D(net487),
    .Q(\s0.data_out[27][6] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _7642_ (.RESET_B(net44),
    .D(net613),
    .Q(\s0.data_out[27][7] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _7643_ (.RESET_B(net43),
    .D(_0121_),
    .Q(\s0.was_valid_out[26] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _7644_ (.RESET_B(net41),
    .D(_0122_),
    .Q(\s0.valid_out[26] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _7645_ (.RESET_B(net40),
    .D(_0123_),
    .Q(\s0.genblk1[25].modules.bubble ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _7646_ (.RESET_B(net39),
    .D(_0124_),
    .Q(\s0.shift_out[26] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _7647_ (.RESET_B(net38),
    .D(_0125_),
    .Q(\s0.data_out[26][0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _7648_ (.RESET_B(net37),
    .D(net671),
    .Q(\s0.data_out[26][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _7649_ (.RESET_B(net36),
    .D(net478),
    .Q(\s0.data_out[26][2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _7650_ (.RESET_B(net35),
    .D(net825),
    .Q(\s0.data_out[26][3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _7651_ (.RESET_B(net34),
    .D(_0129_),
    .Q(\s0.data_out[26][4] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _7652_ (.RESET_B(net33),
    .D(net513),
    .Q(\s0.data_out[26][5] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _7653_ (.RESET_B(net32),
    .D(_0131_),
    .Q(\s0.data_out[26][6] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _7654_ (.RESET_B(net31),
    .D(net537),
    .Q(\s0.data_out[26][7] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _7655_ (.RESET_B(net30),
    .D(net419),
    .Q(\s0.was_valid_out[25] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _7656_ (.RESET_B(net28),
    .D(_0134_),
    .Q(\s0.valid_out[25] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _7657_ (.RESET_B(net27),
    .D(_0135_),
    .Q(\s0.genblk1[24].modules.bubble ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _7658_ (.RESET_B(net26),
    .D(_0136_),
    .Q(\s0.shift_out[25] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _7659_ (.RESET_B(net25),
    .D(net557),
    .Q(\s0.data_out[25][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _7660_ (.RESET_B(net24),
    .D(net768),
    .Q(\s0.data_out[25][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _7661_ (.RESET_B(net367),
    .D(_0139_),
    .Q(\s0.data_out[25][2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _7662_ (.RESET_B(net366),
    .D(net776),
    .Q(\s0.data_out[25][3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _7663_ (.RESET_B(net365),
    .D(_0141_),
    .Q(\s0.data_out[25][4] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _7664_ (.RESET_B(net364),
    .D(_0142_),
    .Q(\s0.data_out[25][5] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _7665_ (.RESET_B(net363),
    .D(_0143_),
    .Q(\s0.data_out[25][6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _7666_ (.RESET_B(net362),
    .D(_0144_),
    .Q(\s0.data_out[25][7] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _7667_ (.RESET_B(net361),
    .D(_0145_),
    .Q(\s0.was_valid_out[24] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _7668_ (.RESET_B(net359),
    .D(_0146_),
    .Q(\s0.valid_out[24] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _7669_ (.RESET_B(net358),
    .D(_0147_),
    .Q(\s0.genblk1[23].modules.bubble ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _7670_ (.RESET_B(net357),
    .D(_0148_),
    .Q(\s0.shift_out[24] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _7671_ (.RESET_B(net356),
    .D(_0149_),
    .Q(\s0.data_out[24][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _7672_ (.RESET_B(net355),
    .D(net510),
    .Q(\s0.data_out[24][1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _7673_ (.RESET_B(net354),
    .D(net632),
    .Q(\s0.data_out[24][2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _7674_ (.RESET_B(net353),
    .D(net503),
    .Q(\s0.data_out[24][3] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _7675_ (.RESET_B(net352),
    .D(net593),
    .Q(\s0.data_out[24][4] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _7676_ (.RESET_B(net351),
    .D(_0154_),
    .Q(\s0.data_out[24][5] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _7677_ (.RESET_B(net350),
    .D(net555),
    .Q(\s0.data_out[24][6] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _7678_ (.RESET_B(net349),
    .D(net541),
    .Q(\s0.data_out[24][7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _7679_ (.RESET_B(net348),
    .D(_0157_),
    .Q(\s0.was_valid_out[23] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _7680_ (.RESET_B(net346),
    .D(_0158_),
    .Q(\s0.valid_out[23] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _7681_ (.RESET_B(net345),
    .D(_0159_),
    .Q(\s0.genblk1[22].modules.bubble ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _7682_ (.RESET_B(net344),
    .D(_0160_),
    .Q(\s0.shift_out[23] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _7683_ (.RESET_B(net343),
    .D(_0161_),
    .Q(\s0.data_out[23][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _7684_ (.RESET_B(net342),
    .D(net818),
    .Q(\s0.data_out[23][1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _7685_ (.RESET_B(net341),
    .D(_0163_),
    .Q(\s0.data_out[23][2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _7686_ (.RESET_B(net340),
    .D(net803),
    .Q(\s0.data_out[23][3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _7687_ (.RESET_B(net339),
    .D(_0165_),
    .Q(\s0.data_out[23][4] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _7688_ (.RESET_B(net338),
    .D(_0166_),
    .Q(\s0.data_out[23][5] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _7689_ (.RESET_B(net337),
    .D(_0167_),
    .Q(\s0.data_out[23][6] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _7690_ (.RESET_B(net336),
    .D(_0168_),
    .Q(\s0.data_out[23][7] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _7691_ (.RESET_B(net335),
    .D(_0169_),
    .Q(\s0.was_valid_out[22] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _7692_ (.RESET_B(net333),
    .D(_0170_),
    .Q(\s0.valid_out[22] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _7693_ (.RESET_B(net332),
    .D(_0171_),
    .Q(\s0.genblk1[21].modules.bubble ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _7694_ (.RESET_B(net331),
    .D(_0172_),
    .Q(\s0.shift_out[22] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _7695_ (.RESET_B(net330),
    .D(_0173_),
    .Q(\s0.data_out[22][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _7696_ (.RESET_B(net329),
    .D(_0174_),
    .Q(\s0.data_out[22][1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _7697_ (.RESET_B(net328),
    .D(_0175_),
    .Q(\s0.data_out[22][2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _7698_ (.RESET_B(net327),
    .D(_0176_),
    .Q(\s0.data_out[22][3] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _7699_ (.RESET_B(net326),
    .D(_0177_),
    .Q(\s0.data_out[22][4] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _7700_ (.RESET_B(net325),
    .D(_0178_),
    .Q(\s0.data_out[22][5] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _7701_ (.RESET_B(net324),
    .D(net489),
    .Q(\s0.data_out[22][6] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _7702_ (.RESET_B(net323),
    .D(net527),
    .Q(\s0.data_out[22][7] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _7703_ (.RESET_B(net322),
    .D(net401),
    .Q(\s0.was_valid_out[21] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _7704_ (.RESET_B(net320),
    .D(_0182_),
    .Q(\s0.valid_out[21] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _7705_ (.RESET_B(net319),
    .D(_0183_),
    .Q(\s0.shift_out[21] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _7706_ (.RESET_B(net318),
    .D(_0184_),
    .Q(\s0.data_out[21][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _7707_ (.RESET_B(net317),
    .D(_0185_),
    .Q(\s0.data_out[21][1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _7708_ (.RESET_B(net316),
    .D(_0186_),
    .Q(\s0.data_out[21][2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _7709_ (.RESET_B(net315),
    .D(net500),
    .Q(\s0.data_out[21][3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _7710_ (.RESET_B(net314),
    .D(_0188_),
    .Q(\s0.data_out[21][4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _7711_ (.RESET_B(net313),
    .D(_0189_),
    .Q(\s0.data_out[21][5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _7712_ (.RESET_B(net312),
    .D(_0190_),
    .Q(\s0.data_out[21][6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _7713_ (.RESET_B(net311),
    .D(net545),
    .Q(\s0.data_out[21][7] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _7714_ (.RESET_B(net310),
    .D(_0192_),
    .Q(\s0.genblk1[20].modules.bubble ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _7715_ (.RESET_B(net309),
    .D(net619),
    .Q(\s0.was_valid_out[20] [0]),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _7716_ (.RESET_B(net307),
    .D(_0194_),
    .Q(\s0.valid_out[20] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _7717_ (.RESET_B(net306),
    .D(_0195_),
    .Q(\s0.genblk1[1].modules.bubble ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _7718_ (.RESET_B(net305),
    .D(_0196_),
    .Q(\s0.shift_out[20] [0]),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _7719_ (.RESET_B(net304),
    .D(_0197_),
    .Q(\s0.data_out[20][0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _7720_ (.RESET_B(net303),
    .D(net561),
    .Q(\s0.data_out[20][1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _7721_ (.RESET_B(net302),
    .D(_0199_),
    .Q(\s0.data_out[20][2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _7722_ (.RESET_B(net301),
    .D(net645),
    .Q(\s0.data_out[20][3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _7723_ (.RESET_B(net300),
    .D(net517),
    .Q(\s0.data_out[20][4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _7724_ (.RESET_B(net299),
    .D(net493),
    .Q(\s0.data_out[20][5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _7725_ (.RESET_B(net298),
    .D(_0203_),
    .Q(\s0.data_out[20][6] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _7726_ (.RESET_B(net297),
    .D(net695),
    .Q(\s0.data_out[20][7] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _7727_ (.RESET_B(net296),
    .D(net410),
    .Q(\s0.was_valid_out[19] [0]),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _7728_ (.RESET_B(net294),
    .D(_0206_),
    .Q(\s0.valid_out[19] [0]),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _7729_ (.RESET_B(net293),
    .D(_0207_),
    .Q(\s0.genblk1[18].modules.bubble ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _7730_ (.RESET_B(net292),
    .D(_0208_),
    .Q(\s0.shift_out[19] [0]),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _7731_ (.RESET_B(net291),
    .D(_0209_),
    .Q(\s0.data_out[19][0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _7732_ (.RESET_B(net290),
    .D(net726),
    .Q(\s0.data_out[19][1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _7733_ (.RESET_B(net289),
    .D(net663),
    .Q(\s0.data_out[19][2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _7734_ (.RESET_B(net288),
    .D(net657),
    .Q(\s0.data_out[19][3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _7735_ (.RESET_B(net287),
    .D(_0213_),
    .Q(\s0.data_out[19][4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _7736_ (.RESET_B(net286),
    .D(_0214_),
    .Q(\s0.data_out[19][5] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _7737_ (.RESET_B(net285),
    .D(net765),
    .Q(\s0.data_out[19][6] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _7738_ (.RESET_B(net284),
    .D(net756),
    .Q(\s0.data_out[19][7] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _7739_ (.RESET_B(net283),
    .D(net827),
    .Q(\s0.was_valid_out[18] [0]),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _7740_ (.RESET_B(net281),
    .D(_0218_),
    .Q(\s0.valid_out[18] [0]),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _7741_ (.RESET_B(net280),
    .D(_0219_),
    .Q(\s0.genblk1[17].modules.bubble ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _7742_ (.RESET_B(net279),
    .D(_0220_),
    .Q(\s0.shift_out[18] [0]),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _7743_ (.RESET_B(net278),
    .D(_0221_),
    .Q(\s0.data_out[18][0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _7744_ (.RESET_B(net277),
    .D(_0222_),
    .Q(\s0.data_out[18][1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _7745_ (.RESET_B(net276),
    .D(_0223_),
    .Q(\s0.data_out[18][2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _7746_ (.RESET_B(net275),
    .D(net483),
    .Q(\s0.data_out[18][3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _7747_ (.RESET_B(net274),
    .D(net599),
    .Q(\s0.data_out[18][4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _7748_ (.RESET_B(net273),
    .D(net575),
    .Q(\s0.data_out[18][5] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _7749_ (.RESET_B(net272),
    .D(_0227_),
    .Q(\s0.data_out[18][6] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _7750_ (.RESET_B(net271),
    .D(_0228_),
    .Q(\s0.data_out[18][7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _7751_ (.RESET_B(net270),
    .D(net421),
    .Q(\s0.was_valid_out[17] [0]),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _7752_ (.RESET_B(net268),
    .D(_0230_),
    .Q(\s0.valid_out[17] [0]),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _7753_ (.RESET_B(net267),
    .D(_0231_),
    .Q(\s0.genblk1[16].modules.bubble ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _7754_ (.RESET_B(net266),
    .D(_0232_),
    .Q(\s0.shift_out[17] [0]),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _7755_ (.RESET_B(net265),
    .D(_0233_),
    .Q(\s0.data_out[17][0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _7756_ (.RESET_B(net264),
    .D(_0234_),
    .Q(\s0.data_out[17][1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _7757_ (.RESET_B(net263),
    .D(_0235_),
    .Q(\s0.data_out[17][2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _7758_ (.RESET_B(net262),
    .D(_0236_),
    .Q(\s0.data_out[17][3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _7759_ (.RESET_B(net261),
    .D(_0237_),
    .Q(\s0.data_out[17][4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _7760_ (.RESET_B(net260),
    .D(_0238_),
    .Q(\s0.data_out[17][5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _7761_ (.RESET_B(net259),
    .D(_0239_),
    .Q(\s0.data_out[17][6] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _7762_ (.RESET_B(net258),
    .D(_0240_),
    .Q(\s0.data_out[17][7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _7763_ (.RESET_B(net257),
    .D(net617),
    .Q(\s0.was_valid_out[16] [0]),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _7764_ (.RESET_B(net255),
    .D(_0242_),
    .Q(\s0.valid_out[16] [0]),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _7765_ (.RESET_B(net254),
    .D(_0243_),
    .Q(\s0.genblk1[15].modules.bubble ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _7766_ (.RESET_B(net253),
    .D(_0244_),
    .Q(\s0.shift_out[16] [0]),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _7767_ (.RESET_B(net252),
    .D(_0245_),
    .Q(\s0.data_out[16][0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _7768_ (.RESET_B(net251),
    .D(net485),
    .Q(\s0.data_out[16][1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _7769_ (.RESET_B(net250),
    .D(net565),
    .Q(\s0.data_out[16][2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _7770_ (.RESET_B(net249),
    .D(net472),
    .Q(\s0.data_out[16][3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _7771_ (.RESET_B(net248),
    .D(net717),
    .Q(\s0.data_out[16][4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _7772_ (.RESET_B(net247),
    .D(_0250_),
    .Q(\s0.data_out[16][5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _7773_ (.RESET_B(net246),
    .D(_0251_),
    .Q(\s0.data_out[16][6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _7774_ (.RESET_B(net245),
    .D(net539),
    .Q(\s0.data_out[16][7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _7775_ (.RESET_B(net244),
    .D(net399),
    .Q(\s0.was_valid_out[15] [0]),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _7776_ (.RESET_B(net242),
    .D(_0254_),
    .Q(\s0.valid_out[15] [0]),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _7777_ (.RESET_B(net241),
    .D(_0255_),
    .Q(\s0.genblk1[14].modules.bubble ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _7778_ (.RESET_B(net240),
    .D(_0256_),
    .Q(\s0.shift_out[15] [0]),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _7779_ (.RESET_B(net239),
    .D(_0257_),
    .Q(\s0.data_out[15][0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _7780_ (.RESET_B(net238),
    .D(net815),
    .Q(\s0.data_out[15][1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _7781_ (.RESET_B(net237),
    .D(_0259_),
    .Q(\s0.data_out[15][2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _7782_ (.RESET_B(net236),
    .D(_0260_),
    .Q(\s0.data_out[15][3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _7783_ (.RESET_B(net235),
    .D(_0261_),
    .Q(\s0.data_out[15][4] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _7784_ (.RESET_B(net234),
    .D(_0262_),
    .Q(\s0.data_out[15][5] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _7785_ (.RESET_B(net233),
    .D(_0263_),
    .Q(\s0.data_out[15][6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _7786_ (.RESET_B(net232),
    .D(net579),
    .Q(\s0.data_out[15][7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _7787_ (.RESET_B(net231),
    .D(net674),
    .Q(\s0.was_valid_out[14] [0]),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _7788_ (.RESET_B(net229),
    .D(_0266_),
    .Q(\s0.valid_out[14] [0]),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _7789_ (.RESET_B(net228),
    .D(_0267_),
    .Q(\s0.genblk1[13].modules.bubble ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _7790_ (.RESET_B(net227),
    .D(_0268_),
    .Q(\s0.shift_out[14] [0]),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _7791_ (.RESET_B(net226),
    .D(_0269_),
    .Q(\s0.data_out[14][0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _7792_ (.RESET_B(net225),
    .D(_0270_),
    .Q(\s0.data_out[14][1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _7793_ (.RESET_B(net224),
    .D(net649),
    .Q(\s0.data_out[14][2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _7794_ (.RESET_B(net223),
    .D(_0272_),
    .Q(\s0.data_out[14][3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _7795_ (.RESET_B(net222),
    .D(_0273_),
    .Q(\s0.data_out[14][4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _7796_ (.RESET_B(net221),
    .D(_0274_),
    .Q(\s0.data_out[14][5] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _7797_ (.RESET_B(net220),
    .D(_0275_),
    .Q(\s0.data_out[14][6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _7798_ (.RESET_B(net219),
    .D(_0276_),
    .Q(\s0.data_out[14][7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _7799_ (.RESET_B(net218),
    .D(net440),
    .Q(\s0.was_valid_out[13] [0]),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _7800_ (.RESET_B(net216),
    .D(_0278_),
    .Q(\s0.valid_out[13] [0]),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _7801_ (.RESET_B(net215),
    .D(_0279_),
    .Q(\s0.genblk1[12].modules.bubble ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _7802_ (.RESET_B(net214),
    .D(_0280_),
    .Q(\s0.shift_out[13] [0]),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _7803_ (.RESET_B(net213),
    .D(_0281_),
    .Q(\s0.data_out[13][0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _7804_ (.RESET_B(net212),
    .D(_0282_),
    .Q(\s0.data_out[13][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _7805_ (.RESET_B(net211),
    .D(_0283_),
    .Q(\s0.data_out[13][2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _7806_ (.RESET_B(net210),
    .D(net693),
    .Q(\s0.data_out[13][3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _7807_ (.RESET_B(net209),
    .D(net519),
    .Q(\s0.data_out[13][4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _7808_ (.RESET_B(net208),
    .D(net584),
    .Q(\s0.data_out[13][5] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _7809_ (.RESET_B(net207),
    .D(_0287_),
    .Q(\s0.data_out[13][6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _7810_ (.RESET_B(net206),
    .D(net609),
    .Q(\s0.data_out[13][7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _7811_ (.RESET_B(net205),
    .D(_0289_),
    .Q(\s0.was_valid_out[12] [0]),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _7812_ (.RESET_B(net203),
    .D(_0290_),
    .Q(\s0.valid_out[12] [0]),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _7813_ (.RESET_B(net202),
    .D(_0291_),
    .Q(\s0.genblk1[11].modules.bubble ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _7814_ (.RESET_B(net201),
    .D(_0292_),
    .Q(\s0.shift_out[12] [0]),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _7815_ (.RESET_B(net200),
    .D(_0293_),
    .Q(\s0.data_out[12][0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _7816_ (.RESET_B(net199),
    .D(net821),
    .Q(\s0.data_out[12][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _7817_ (.RESET_B(net198),
    .D(net750),
    .Q(\s0.data_out[12][2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _7818_ (.RESET_B(net197),
    .D(net581),
    .Q(\s0.data_out[12][3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _7819_ (.RESET_B(net196),
    .D(_0297_),
    .Q(\s0.data_out[12][4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _7820_ (.RESET_B(net195),
    .D(net661),
    .Q(\s0.data_out[12][5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _7821_ (.RESET_B(net194),
    .D(_0299_),
    .Q(\s0.data_out[12][6] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _7822_ (.RESET_B(net193),
    .D(net523),
    .Q(\s0.data_out[12][7] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _7823_ (.RESET_B(net192),
    .D(net446),
    .Q(\s0.was_valid_out[11] [0]),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _7824_ (.RESET_B(net190),
    .D(_0302_),
    .Q(\s0.valid_out[11] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _7825_ (.RESET_B(net189),
    .D(_0303_),
    .Q(\s0.genblk1[10].modules.bubble ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7826_ (.RESET_B(net188),
    .D(_0304_),
    .Q(\s0.shift_out[11] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _7827_ (.RESET_B(net187),
    .D(_0305_),
    .Q(\s0.data_out[11][0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _7828_ (.RESET_B(net186),
    .D(_0306_),
    .Q(\s0.data_out[11][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _7829_ (.RESET_B(net185),
    .D(_0307_),
    .Q(\s0.data_out[11][2] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7830_ (.RESET_B(net184),
    .D(net747),
    .Q(\s0.data_out[11][3] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7831_ (.RESET_B(net183),
    .D(net789),
    .Q(\s0.data_out[11][4] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7832_ (.RESET_B(net182),
    .D(net606),
    .Q(\s0.data_out[11][5] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _7833_ (.RESET_B(net181),
    .D(_0311_),
    .Q(\s0.data_out[11][6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _7834_ (.RESET_B(net180),
    .D(net569),
    .Q(\s0.data_out[11][7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _7835_ (.RESET_B(net179),
    .D(_0313_),
    .Q(\s0.was_valid_out[10] [0]),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _7836_ (.RESET_B(net177),
    .D(_0314_),
    .Q(\s0.valid_out[10] [0]),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _7837_ (.RESET_B(net176),
    .D(_0315_),
    .Q(\s0.data_new_delayed[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _7838_ (.RESET_B(net175),
    .D(_0316_),
    .Q(\s0.data_new_delayed[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _7839_ (.RESET_B(net174),
    .D(_0317_),
    .Q(\s0.data_new_delayed[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _7840_ (.RESET_B(net173),
    .D(_0318_),
    .Q(\s0.data_new_delayed[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _7841_ (.RESET_B(net172),
    .D(_0319_),
    .Q(\s0.data_new_delayed[4] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _7842_ (.RESET_B(net171),
    .D(_0320_),
    .Q(\s0.data_new_delayed[5] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _7843_ (.RESET_B(net170),
    .D(_0321_),
    .Q(\s0.data_new_delayed[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _7844_ (.RESET_B(net169),
    .D(_0322_),
    .Q(\s0.data_new_delayed[7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _7845_ (.RESET_B(net168),
    .D(_0323_),
    .Q(\s0.shift_out[10] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _7846_ (.RESET_B(net167),
    .D(_0324_),
    .Q(\s0.data_out[10][0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _7847_ (.RESET_B(net166),
    .D(_0325_),
    .Q(\s0.data_out[10][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _7848_ (.RESET_B(net165),
    .D(net480),
    .Q(\s0.data_out[10][2] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7849_ (.RESET_B(net164),
    .D(net667),
    .Q(\s0.data_out[10][3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7850_ (.RESET_B(net163),
    .D(_0328_),
    .Q(\s0.data_out[10][4] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7851_ (.RESET_B(net162),
    .D(net498),
    .Q(\s0.data_out[10][5] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _7852_ (.RESET_B(net161),
    .D(_0330_),
    .Q(\s0.data_out[10][6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _7853_ (.RESET_B(net160),
    .D(net515),
    .Q(\s0.data_out[10][7] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _7854_ (.RESET_B(net159),
    .D(net448),
    .Q(\s0.was_valid_out[9] [0]),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _7855_ (.RESET_B(net157),
    .D(_0333_),
    .Q(\s0.valid_out[9] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _7856_ (.RESET_B(net156),
    .D(_0334_),
    .Q(\s0.genblk1[8].modules.bubble ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _7857_ (.RESET_B(net155),
    .D(_0335_),
    .Q(\s0.shift_out[9] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _7858_ (.RESET_B(net154),
    .D(_0336_),
    .Q(\s0.data_out[9][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _7859_ (.RESET_B(net153),
    .D(net476),
    .Q(\s0.data_out[9][1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _7860_ (.RESET_B(net152),
    .D(net491),
    .Q(\s0.data_out[9][2] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7861_ (.RESET_B(net151),
    .D(_0339_),
    .Q(\s0.data_out[9][3] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7862_ (.RESET_B(net150),
    .D(_0340_),
    .Q(\s0.data_out[9][4] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7863_ (.RESET_B(net149),
    .D(_0341_),
    .Q(\s0.data_out[9][5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _7864_ (.RESET_B(net148),
    .D(_0342_),
    .Q(\s0.data_out[9][6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _7865_ (.RESET_B(net147),
    .D(net535),
    .Q(\s0.data_out[9][7] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _7866_ (.RESET_B(net146),
    .D(_0000_),
    .Q(\s0.was_valid_out[8] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _7867_ (.RESET_B(net144),
    .D(_0001_),
    .Q(\s0.valid_out[8] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _7868_ (.RESET_B(net143),
    .D(_0002_),
    .Q(\s0.genblk1[7].modules.bubble ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _7869_ (.RESET_B(net142),
    .D(_0003_),
    .Q(\s0.shift_out[8] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _7870_ (.RESET_B(net141),
    .D(_0004_),
    .Q(\s0.data_out[8][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _7871_ (.RESET_B(net140),
    .D(net595),
    .Q(\s0.data_out[8][1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _7872_ (.RESET_B(net139),
    .D(net563),
    .Q(\s0.data_out[8][2] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7873_ (.RESET_B(net138),
    .D(_0007_),
    .Q(\s0.data_out[8][3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7874_ (.RESET_B(net137),
    .D(_0008_),
    .Q(\s0.data_out[8][4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _7875_ (.RESET_B(net136),
    .D(_0009_),
    .Q(\s0.data_out[8][5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _7876_ (.RESET_B(net135),
    .D(net641),
    .Q(\s0.data_out[8][6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _7877_ (.RESET_B(net134),
    .D(_0011_),
    .Q(\s0.data_out[8][7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _7878_ (.RESET_B(net133),
    .D(_0012_),
    .Q(\s0.was_valid_out[7] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _7879_ (.RESET_B(net131),
    .D(_0013_),
    .Q(\s0.valid_out[7] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _7880_ (.RESET_B(net130),
    .D(_0014_),
    .Q(\s0.genblk1[6].modules.bubble ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _7881_ (.RESET_B(net129),
    .D(_0015_),
    .Q(\s0.shift_out[7] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _7882_ (.RESET_B(net128),
    .D(_0016_),
    .Q(\s0.data_out[7][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _7883_ (.RESET_B(net127),
    .D(net797),
    .Q(\s0.data_out[7][1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _7884_ (.RESET_B(net126),
    .D(net591),
    .Q(\s0.data_out[7][2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _7885_ (.RESET_B(net125),
    .D(net577),
    .Q(\s0.data_out[7][3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7886_ (.RESET_B(net124),
    .D(_0020_),
    .Q(\s0.data_out[7][4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _7887_ (.RESET_B(net123),
    .D(_0021_),
    .Q(\s0.data_out[7][5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _7888_ (.RESET_B(net122),
    .D(_0022_),
    .Q(\s0.data_out[7][6] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _7889_ (.RESET_B(net121),
    .D(_0023_),
    .Q(\s0.data_out[7][7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _7890_ (.RESET_B(net120),
    .D(net423),
    .Q(\s0.was_valid_out[6] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _7891_ (.RESET_B(net118),
    .D(_0025_),
    .Q(\s0.valid_out[6] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _7892_ (.RESET_B(net117),
    .D(_0026_),
    .Q(\s0.genblk1[5].modules.bubble ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _7893_ (.RESET_B(net116),
    .D(_0027_),
    .Q(\s0.shift_out[6] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _7894_ (.RESET_B(net115),
    .D(_0028_),
    .Q(\s0.data_out[6][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _7895_ (.RESET_B(net114),
    .D(_0029_),
    .Q(\s0.data_out[6][1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _7896_ (.RESET_B(net113),
    .D(_0030_),
    .Q(\s0.data_out[6][2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _7897_ (.RESET_B(net112),
    .D(net428),
    .Q(\s0.data_out[6][3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _7898_ (.RESET_B(net111),
    .D(_0032_),
    .Q(\s0.data_out[6][4] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _7899_ (.RESET_B(net110),
    .D(_0033_),
    .Q(\s0.data_out[6][5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _7900_ (.RESET_B(net109),
    .D(_0034_),
    .Q(\s0.data_out[6][6] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _7901_ (.RESET_B(net108),
    .D(_0035_),
    .Q(\s0.data_out[6][7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _7902_ (.RESET_B(net107),
    .D(_0036_),
    .Q(\s0.was_valid_out[5] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _7903_ (.RESET_B(net105),
    .D(_0037_),
    .Q(\s0.valid_out[5] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _7904_ (.RESET_B(net104),
    .D(_0038_),
    .Q(\s0.genblk1[4].modules.bubble ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _7905_ (.RESET_B(net103),
    .D(_0039_),
    .Q(\s0.shift_out[5] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _7906_ (.RESET_B(net102),
    .D(_0040_),
    .Q(\s0.data_out[5][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _7907_ (.RESET_B(net101),
    .D(net547),
    .Q(\s0.data_out[5][1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _7908_ (.RESET_B(net100),
    .D(net647),
    .Q(\s0.data_out[5][2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _7909_ (.RESET_B(net99),
    .D(net573),
    .Q(\s0.data_out[5][3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _7910_ (.RESET_B(net98),
    .D(_0044_),
    .Q(\s0.data_out[5][4] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _7911_ (.RESET_B(net97),
    .D(net652),
    .Q(\s0.data_out[5][5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _7912_ (.RESET_B(net96),
    .D(net597),
    .Q(\s0.data_out[5][6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _7913_ (.RESET_B(net95),
    .D(net529),
    .Q(\s0.data_out[5][7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _7914_ (.RESET_B(net94),
    .D(net417),
    .Q(\s0.was_valid_out[4] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _7915_ (.RESET_B(net92),
    .D(_0049_),
    .Q(\s0.valid_out[4] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _7916_ (.RESET_B(net91),
    .D(_0050_),
    .Q(\s0.genblk1[3].modules.bubble ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _7917_ (.RESET_B(net90),
    .D(_0051_),
    .Q(\s0.shift_out[4] [0]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _7918_ (.RESET_B(net89),
    .D(_0052_),
    .Q(\s0.data_out[4][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _7919_ (.RESET_B(net88),
    .D(_0053_),
    .Q(\s0.data_out[4][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _7920_ (.RESET_B(net87),
    .D(_0054_),
    .Q(\s0.data_out[4][2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _7921_ (.RESET_B(net86),
    .D(_0055_),
    .Q(\s0.data_out[4][3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _7922_ (.RESET_B(net85),
    .D(_0056_),
    .Q(\s0.data_out[4][4] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _7923_ (.RESET_B(net84),
    .D(_0057_),
    .Q(\s0.data_out[4][5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _7924_ (.RESET_B(net83),
    .D(net559),
    .Q(\s0.data_out[4][6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _7925_ (.RESET_B(net82),
    .D(net625),
    .Q(\s0.data_out[4][7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _7926_ (.RESET_B(net81),
    .D(net407),
    .Q(\s0.was_valid_out[3] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _7927_ (.RESET_B(net79),
    .D(_0061_),
    .Q(\s0.valid_out[3] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _7928_ (.RESET_B(net78),
    .D(_0062_),
    .Q(\s0.genblk1[2].modules.bubble ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _7929_ (.RESET_B(net77),
    .D(_0063_),
    .Q(\s0.shift_out[3] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _7930_ (.RESET_B(net76),
    .D(_0064_),
    .Q(\s0.data_out[3][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _7931_ (.RESET_B(net75),
    .D(_0065_),
    .Q(\s0.data_out[3][1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _7932_ (.RESET_B(net74),
    .D(_0066_),
    .Q(\s0.data_out[3][2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _7933_ (.RESET_B(net73),
    .D(_0067_),
    .Q(\s0.data_out[3][3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _7934_ (.RESET_B(net72),
    .D(net701),
    .Q(\s0.data_out[3][4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _7935_ (.RESET_B(net71),
    .D(_0069_),
    .Q(\s0.data_out[3][5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _7936_ (.RESET_B(net70),
    .D(_0070_),
    .Q(\s0.data_out[3][6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _7937_ (.RESET_B(net69),
    .D(net635),
    .Q(\s0.data_out[3][7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _7938_ (.RESET_B(net68),
    .D(net433),
    .Q(\s0.was_valid_out[2] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _7939_ (.RESET_B(net66),
    .D(_0073_),
    .Q(\s0.valid_out[2] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _7940_ (.RESET_B(net65),
    .D(_0074_),
    .Q(\s0.genblk1[27].modules.bubble ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _7941_ (.RESET_B(net64),
    .D(_0075_),
    .Q(\s0.shift_out[2] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _7942_ (.RESET_B(net63),
    .D(_0076_),
    .Q(\s0.data_out[2][0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _7943_ (.RESET_B(net62),
    .D(_0077_),
    .Q(\s0.data_out[2][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _7944_ (.RESET_B(net61),
    .D(_0078_),
    .Q(\s0.data_out[2][2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _7945_ (.RESET_B(net60),
    .D(net785),
    .Q(\s0.data_out[2][3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _7946_ (.RESET_B(net59),
    .D(_0080_),
    .Q(\s0.data_out[2][4] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _7947_ (.RESET_B(net58),
    .D(_0081_),
    .Q(\s0.data_out[2][5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _7948_ (.RESET_B(net57),
    .D(_0082_),
    .Q(\s0.data_out[2][6] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _7949_ (.RESET_B(net55),
    .D(net543),
    .Q(\s0.data_out[2][7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _7950_ (.RESET_B(net42),
    .D(_0084_),
    .Q(\s0.was_valid_out[1] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _7951_ (.RESET_B(net360),
    .D(_0085_),
    .Q(\s0.valid_out[1] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _7952_ (.RESET_B(net347),
    .D(_0086_),
    .Q(\s0.genblk1[19].modules.bubble ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _7953_ (.RESET_B(net334),
    .D(_0087_),
    .Q(\s0.shift_out[1] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _7954_ (.RESET_B(net321),
    .D(_0088_),
    .Q(\s0.data_out[1][0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _7955_ (.RESET_B(net308),
    .D(_0089_),
    .Q(\s0.data_out[1][1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _7956_ (.RESET_B(net295),
    .D(_0090_),
    .Q(\s0.data_out[1][2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _7957_ (.RESET_B(net282),
    .D(_0091_),
    .Q(\s0.data_out[1][3] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _7958_ (.RESET_B(net269),
    .D(_0092_),
    .Q(\s0.data_out[1][4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _7959_ (.RESET_B(net256),
    .D(_0093_),
    .Q(\s0.data_out[1][5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _7960_ (.RESET_B(net243),
    .D(_0094_),
    .Q(\s0.data_out[1][6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _7961_ (.RESET_B(net230),
    .D(_0095_),
    .Q(\s0.data_out[1][7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _7962_ (.RESET_B(net217),
    .D(_0096_),
    .Q(\s0.was_valid_out[0] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _7963_ (.RESET_B(net191),
    .D(_0097_),
    .Q(\s0.valid_out[0] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _7964_ (.RESET_B(net178),
    .D(_0098_),
    .Q(\s0.genblk1[9].modules.bubble ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _7965_ (.RESET_B(net158),
    .D(_0099_),
    .Q(\s0.shift_out[0] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _7966_ (.RESET_B(net145),
    .D(_0100_),
    .Q(\s0.data_out[0][0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _7967_ (.RESET_B(net132),
    .D(_0101_),
    .Q(\s0.data_out[0][1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _7968_ (.RESET_B(net119),
    .D(_0102_),
    .Q(\s0.data_out[0][2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _7969_ (.RESET_B(net106),
    .D(net442),
    .Q(\s0.data_out[0][3] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _7970_ (.RESET_B(net93),
    .D(_0104_),
    .Q(\s0.data_out[0][4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _7971_ (.RESET_B(net80),
    .D(_0105_),
    .Q(\s0.data_out[0][5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _7972_ (.RESET_B(net67),
    .D(_0106_),
    .Q(\s0.data_out[0][6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _7973_ (.RESET_B(net29),
    .D(_0107_),
    .Q(\s0.data_out[0][7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_tiehi _7659__25 (.L_HI(net25));
 sg13g2_tiehi _7658__26 (.L_HI(net26));
 sg13g2_tiehi _7657__27 (.L_HI(net27));
 sg13g2_tiehi _7656__28 (.L_HI(net28));
 sg13g2_tiehi _7973__29 (.L_HI(net29));
 sg13g2_tiehi _7655__30 (.L_HI(net30));
 sg13g2_tiehi _7654__31 (.L_HI(net31));
 sg13g2_tiehi _7653__32 (.L_HI(net32));
 sg13g2_tiehi _7652__33 (.L_HI(net33));
 sg13g2_tiehi _7651__34 (.L_HI(net34));
 sg13g2_tiehi _7650__35 (.L_HI(net35));
 sg13g2_tiehi _7649__36 (.L_HI(net36));
 sg13g2_tiehi _7648__37 (.L_HI(net37));
 sg13g2_tiehi _7647__38 (.L_HI(net38));
 sg13g2_tiehi _7646__39 (.L_HI(net39));
 sg13g2_tiehi _7645__40 (.L_HI(net40));
 sg13g2_tiehi _7644__41 (.L_HI(net41));
 sg13g2_tiehi _7950__42 (.L_HI(net42));
 sg13g2_tiehi _7643__43 (.L_HI(net43));
 sg13g2_tiehi _7642__44 (.L_HI(net44));
 sg13g2_tiehi _7641__45 (.L_HI(net45));
 sg13g2_tiehi _7640__46 (.L_HI(net46));
 sg13g2_tiehi _7639__47 (.L_HI(net47));
 sg13g2_tiehi _7638__48 (.L_HI(net48));
 sg13g2_tiehi _7637__49 (.L_HI(net49));
 sg13g2_tiehi _7636__50 (.L_HI(net50));
 sg13g2_tiehi _7635__51 (.L_HI(net51));
 sg13g2_tiehi _7634__52 (.L_HI(net52));
 sg13g2_tiehi _7633__53 (.L_HI(net53));
 sg13g2_tiehi _7632__54 (.L_HI(net54));
 sg13g2_tiehi _7949__55 (.L_HI(net55));
 sg13g2_tiehi _7631__56 (.L_HI(net56));
 sg13g2_tiehi _7948__57 (.L_HI(net57));
 sg13g2_tiehi _7947__58 (.L_HI(net58));
 sg13g2_tiehi _7946__59 (.L_HI(net59));
 sg13g2_tiehi _7945__60 (.L_HI(net60));
 sg13g2_tiehi _7944__61 (.L_HI(net61));
 sg13g2_tiehi _7943__62 (.L_HI(net62));
 sg13g2_tiehi _7942__63 (.L_HI(net63));
 sg13g2_tiehi _7941__64 (.L_HI(net64));
 sg13g2_tiehi _7940__65 (.L_HI(net65));
 sg13g2_tiehi _7939__66 (.L_HI(net66));
 sg13g2_tiehi _7972__67 (.L_HI(net67));
 sg13g2_tiehi _7938__68 (.L_HI(net68));
 sg13g2_tiehi _7937__69 (.L_HI(net69));
 sg13g2_tiehi _7936__70 (.L_HI(net70));
 sg13g2_tiehi _7935__71 (.L_HI(net71));
 sg13g2_tiehi _7934__72 (.L_HI(net72));
 sg13g2_tiehi _7933__73 (.L_HI(net73));
 sg13g2_tiehi _7932__74 (.L_HI(net74));
 sg13g2_tiehi _7931__75 (.L_HI(net75));
 sg13g2_tiehi _7930__76 (.L_HI(net76));
 sg13g2_tiehi _7929__77 (.L_HI(net77));
 sg13g2_tiehi _7928__78 (.L_HI(net78));
 sg13g2_tiehi _7927__79 (.L_HI(net79));
 sg13g2_tiehi _7971__80 (.L_HI(net80));
 sg13g2_tiehi _7926__81 (.L_HI(net81));
 sg13g2_tiehi _7925__82 (.L_HI(net82));
 sg13g2_tiehi _7924__83 (.L_HI(net83));
 sg13g2_tiehi _7923__84 (.L_HI(net84));
 sg13g2_tiehi _7922__85 (.L_HI(net85));
 sg13g2_tiehi _7921__86 (.L_HI(net86));
 sg13g2_tiehi _7920__87 (.L_HI(net87));
 sg13g2_tiehi _7919__88 (.L_HI(net88));
 sg13g2_tiehi _7918__89 (.L_HI(net89));
 sg13g2_tiehi _7917__90 (.L_HI(net90));
 sg13g2_tiehi _7916__91 (.L_HI(net91));
 sg13g2_tiehi _7915__92 (.L_HI(net92));
 sg13g2_tiehi _7970__93 (.L_HI(net93));
 sg13g2_tiehi _7914__94 (.L_HI(net94));
 sg13g2_tiehi _7913__95 (.L_HI(net95));
 sg13g2_tiehi _7912__96 (.L_HI(net96));
 sg13g2_tiehi _7911__97 (.L_HI(net97));
 sg13g2_tiehi _7910__98 (.L_HI(net98));
 sg13g2_tiehi _7909__99 (.L_HI(net99));
 sg13g2_tiehi _7908__100 (.L_HI(net100));
 sg13g2_tiehi _7907__101 (.L_HI(net101));
 sg13g2_tiehi _7906__102 (.L_HI(net102));
 sg13g2_tiehi _7905__103 (.L_HI(net103));
 sg13g2_tiehi _7904__104 (.L_HI(net104));
 sg13g2_tiehi _7903__105 (.L_HI(net105));
 sg13g2_tiehi _7969__106 (.L_HI(net106));
 sg13g2_tiehi _7902__107 (.L_HI(net107));
 sg13g2_tiehi _7901__108 (.L_HI(net108));
 sg13g2_tiehi _7900__109 (.L_HI(net109));
 sg13g2_tiehi _7899__110 (.L_HI(net110));
 sg13g2_tiehi _7898__111 (.L_HI(net111));
 sg13g2_tiehi _7897__112 (.L_HI(net112));
 sg13g2_tiehi _7896__113 (.L_HI(net113));
 sg13g2_tiehi _7895__114 (.L_HI(net114));
 sg13g2_tiehi _7894__115 (.L_HI(net115));
 sg13g2_tiehi _7893__116 (.L_HI(net116));
 sg13g2_tiehi _7892__117 (.L_HI(net117));
 sg13g2_tiehi _7891__118 (.L_HI(net118));
 sg13g2_tiehi _7968__119 (.L_HI(net119));
 sg13g2_tiehi _7890__120 (.L_HI(net120));
 sg13g2_tiehi _7889__121 (.L_HI(net121));
 sg13g2_tiehi _7888__122 (.L_HI(net122));
 sg13g2_tiehi _7887__123 (.L_HI(net123));
 sg13g2_tiehi _7886__124 (.L_HI(net124));
 sg13g2_tiehi _7885__125 (.L_HI(net125));
 sg13g2_tiehi _7884__126 (.L_HI(net126));
 sg13g2_tiehi _7883__127 (.L_HI(net127));
 sg13g2_tiehi _7882__128 (.L_HI(net128));
 sg13g2_tiehi _7881__129 (.L_HI(net129));
 sg13g2_tiehi _7880__130 (.L_HI(net130));
 sg13g2_tiehi _7879__131 (.L_HI(net131));
 sg13g2_tiehi _7967__132 (.L_HI(net132));
 sg13g2_tiehi _7878__133 (.L_HI(net133));
 sg13g2_tiehi _7877__134 (.L_HI(net134));
 sg13g2_tiehi _7876__135 (.L_HI(net135));
 sg13g2_tiehi _7875__136 (.L_HI(net136));
 sg13g2_tiehi _7874__137 (.L_HI(net137));
 sg13g2_tiehi _7873__138 (.L_HI(net138));
 sg13g2_tiehi _7872__139 (.L_HI(net139));
 sg13g2_tiehi _7871__140 (.L_HI(net140));
 sg13g2_tiehi _7870__141 (.L_HI(net141));
 sg13g2_tiehi _7869__142 (.L_HI(net142));
 sg13g2_tiehi _7868__143 (.L_HI(net143));
 sg13g2_tiehi _7867__144 (.L_HI(net144));
 sg13g2_tiehi _7966__145 (.L_HI(net145));
 sg13g2_tiehi _7866__146 (.L_HI(net146));
 sg13g2_tiehi _7865__147 (.L_HI(net147));
 sg13g2_tiehi _7864__148 (.L_HI(net148));
 sg13g2_tiehi _7863__149 (.L_HI(net149));
 sg13g2_tiehi _7862__150 (.L_HI(net150));
 sg13g2_tiehi _7861__151 (.L_HI(net151));
 sg13g2_tiehi _7860__152 (.L_HI(net152));
 sg13g2_tiehi _7859__153 (.L_HI(net153));
 sg13g2_tiehi _7858__154 (.L_HI(net154));
 sg13g2_tiehi _7857__155 (.L_HI(net155));
 sg13g2_tiehi _7856__156 (.L_HI(net156));
 sg13g2_tiehi _7855__157 (.L_HI(net157));
 sg13g2_tiehi _7965__158 (.L_HI(net158));
 sg13g2_tiehi _7854__159 (.L_HI(net159));
 sg13g2_tiehi _7853__160 (.L_HI(net160));
 sg13g2_tiehi _7852__161 (.L_HI(net161));
 sg13g2_tiehi _7851__162 (.L_HI(net162));
 sg13g2_tiehi _7850__163 (.L_HI(net163));
 sg13g2_tiehi _7849__164 (.L_HI(net164));
 sg13g2_tiehi _7848__165 (.L_HI(net165));
 sg13g2_tiehi _7847__166 (.L_HI(net166));
 sg13g2_tiehi _7846__167 (.L_HI(net167));
 sg13g2_tiehi _7845__168 (.L_HI(net168));
 sg13g2_tiehi _7844__169 (.L_HI(net169));
 sg13g2_tiehi _7843__170 (.L_HI(net170));
 sg13g2_tiehi _7842__171 (.L_HI(net171));
 sg13g2_tiehi _7841__172 (.L_HI(net172));
 sg13g2_tiehi _7840__173 (.L_HI(net173));
 sg13g2_tiehi _7839__174 (.L_HI(net174));
 sg13g2_tiehi _7838__175 (.L_HI(net175));
 sg13g2_tiehi _7837__176 (.L_HI(net176));
 sg13g2_tiehi _7836__177 (.L_HI(net177));
 sg13g2_tiehi _7964__178 (.L_HI(net178));
 sg13g2_tiehi _7835__179 (.L_HI(net179));
 sg13g2_tiehi _7834__180 (.L_HI(net180));
 sg13g2_tiehi _7833__181 (.L_HI(net181));
 sg13g2_tiehi _7832__182 (.L_HI(net182));
 sg13g2_tiehi _7831__183 (.L_HI(net183));
 sg13g2_tiehi _7830__184 (.L_HI(net184));
 sg13g2_tiehi _7829__185 (.L_HI(net185));
 sg13g2_tiehi _7828__186 (.L_HI(net186));
 sg13g2_tiehi _7827__187 (.L_HI(net187));
 sg13g2_tiehi _7826__188 (.L_HI(net188));
 sg13g2_tiehi _7825__189 (.L_HI(net189));
 sg13g2_tiehi _7824__190 (.L_HI(net190));
 sg13g2_tiehi _7963__191 (.L_HI(net191));
 sg13g2_tiehi _7823__192 (.L_HI(net192));
 sg13g2_tiehi _7822__193 (.L_HI(net193));
 sg13g2_tiehi _7821__194 (.L_HI(net194));
 sg13g2_tiehi _7820__195 (.L_HI(net195));
 sg13g2_tiehi _7819__196 (.L_HI(net196));
 sg13g2_tiehi _7818__197 (.L_HI(net197));
 sg13g2_tiehi _7817__198 (.L_HI(net198));
 sg13g2_tiehi _7816__199 (.L_HI(net199));
 sg13g2_tiehi _7815__200 (.L_HI(net200));
 sg13g2_tiehi _7814__201 (.L_HI(net201));
 sg13g2_tiehi _7813__202 (.L_HI(net202));
 sg13g2_tiehi _7812__203 (.L_HI(net203));
 sg13g2_tiehi _7630__204 (.L_HI(net204));
 sg13g2_tiehi _7811__205 (.L_HI(net205));
 sg13g2_tiehi _7810__206 (.L_HI(net206));
 sg13g2_tiehi _7809__207 (.L_HI(net207));
 sg13g2_tiehi _7808__208 (.L_HI(net208));
 sg13g2_tiehi _7807__209 (.L_HI(net209));
 sg13g2_tiehi _7806__210 (.L_HI(net210));
 sg13g2_tiehi _7805__211 (.L_HI(net211));
 sg13g2_tiehi _7804__212 (.L_HI(net212));
 sg13g2_tiehi _7803__213 (.L_HI(net213));
 sg13g2_tiehi _7802__214 (.L_HI(net214));
 sg13g2_tiehi _7801__215 (.L_HI(net215));
 sg13g2_tiehi _7800__216 (.L_HI(net216));
 sg13g2_tiehi _7962__217 (.L_HI(net217));
 sg13g2_tiehi _7799__218 (.L_HI(net218));
 sg13g2_tiehi _7798__219 (.L_HI(net219));
 sg13g2_tiehi _7797__220 (.L_HI(net220));
 sg13g2_tiehi _7796__221 (.L_HI(net221));
 sg13g2_tiehi _7795__222 (.L_HI(net222));
 sg13g2_tiehi _7794__223 (.L_HI(net223));
 sg13g2_tiehi _7793__224 (.L_HI(net224));
 sg13g2_tiehi _7792__225 (.L_HI(net225));
 sg13g2_tiehi _7791__226 (.L_HI(net226));
 sg13g2_tiehi _7790__227 (.L_HI(net227));
 sg13g2_tiehi _7789__228 (.L_HI(net228));
 sg13g2_tiehi _7788__229 (.L_HI(net229));
 sg13g2_tiehi _7961__230 (.L_HI(net230));
 sg13g2_tiehi _7787__231 (.L_HI(net231));
 sg13g2_tiehi _7786__232 (.L_HI(net232));
 sg13g2_tiehi _7785__233 (.L_HI(net233));
 sg13g2_tiehi _7784__234 (.L_HI(net234));
 sg13g2_tiehi _7783__235 (.L_HI(net235));
 sg13g2_tiehi _7782__236 (.L_HI(net236));
 sg13g2_tiehi _7781__237 (.L_HI(net237));
 sg13g2_tiehi _7780__238 (.L_HI(net238));
 sg13g2_tiehi _7779__239 (.L_HI(net239));
 sg13g2_tiehi _7778__240 (.L_HI(net240));
 sg13g2_tiehi _7777__241 (.L_HI(net241));
 sg13g2_tiehi _7776__242 (.L_HI(net242));
 sg13g2_tiehi _7960__243 (.L_HI(net243));
 sg13g2_tiehi _7775__244 (.L_HI(net244));
 sg13g2_tiehi _7774__245 (.L_HI(net245));
 sg13g2_tiehi _7773__246 (.L_HI(net246));
 sg13g2_tiehi _7772__247 (.L_HI(net247));
 sg13g2_tiehi _7771__248 (.L_HI(net248));
 sg13g2_tiehi _7770__249 (.L_HI(net249));
 sg13g2_tiehi _7769__250 (.L_HI(net250));
 sg13g2_tiehi _7768__251 (.L_HI(net251));
 sg13g2_tiehi _7767__252 (.L_HI(net252));
 sg13g2_tiehi _7766__253 (.L_HI(net253));
 sg13g2_tiehi _7765__254 (.L_HI(net254));
 sg13g2_tiehi _7764__255 (.L_HI(net255));
 sg13g2_tiehi _7959__256 (.L_HI(net256));
 sg13g2_tiehi _7763__257 (.L_HI(net257));
 sg13g2_tiehi _7762__258 (.L_HI(net258));
 sg13g2_tiehi _7761__259 (.L_HI(net259));
 sg13g2_tiehi _7760__260 (.L_HI(net260));
 sg13g2_tiehi _7759__261 (.L_HI(net261));
 sg13g2_tiehi _7758__262 (.L_HI(net262));
 sg13g2_tiehi _7757__263 (.L_HI(net263));
 sg13g2_tiehi _7756__264 (.L_HI(net264));
 sg13g2_tiehi _7755__265 (.L_HI(net265));
 sg13g2_tiehi _7754__266 (.L_HI(net266));
 sg13g2_tiehi _7753__267 (.L_HI(net267));
 sg13g2_tiehi _7752__268 (.L_HI(net268));
 sg13g2_tiehi _7958__269 (.L_HI(net269));
 sg13g2_tiehi _7751__270 (.L_HI(net270));
 sg13g2_tiehi _7750__271 (.L_HI(net271));
 sg13g2_tiehi _7749__272 (.L_HI(net272));
 sg13g2_tiehi _7748__273 (.L_HI(net273));
 sg13g2_tiehi _7747__274 (.L_HI(net274));
 sg13g2_tiehi _7746__275 (.L_HI(net275));
 sg13g2_tiehi _7745__276 (.L_HI(net276));
 sg13g2_tiehi _7744__277 (.L_HI(net277));
 sg13g2_tiehi _7743__278 (.L_HI(net278));
 sg13g2_tiehi _7742__279 (.L_HI(net279));
 sg13g2_tiehi _7741__280 (.L_HI(net280));
 sg13g2_tiehi _7740__281 (.L_HI(net281));
 sg13g2_tiehi _7957__282 (.L_HI(net282));
 sg13g2_tiehi _7739__283 (.L_HI(net283));
 sg13g2_tiehi _7738__284 (.L_HI(net284));
 sg13g2_tiehi _7737__285 (.L_HI(net285));
 sg13g2_tiehi _7736__286 (.L_HI(net286));
 sg13g2_tiehi _7735__287 (.L_HI(net287));
 sg13g2_tiehi _7734__288 (.L_HI(net288));
 sg13g2_tiehi _7733__289 (.L_HI(net289));
 sg13g2_tiehi _7732__290 (.L_HI(net290));
 sg13g2_tiehi _7731__291 (.L_HI(net291));
 sg13g2_tiehi _7730__292 (.L_HI(net292));
 sg13g2_tiehi _7729__293 (.L_HI(net293));
 sg13g2_tiehi _7728__294 (.L_HI(net294));
 sg13g2_tiehi _7956__295 (.L_HI(net295));
 sg13g2_tiehi _7727__296 (.L_HI(net296));
 sg13g2_tiehi _7726__297 (.L_HI(net297));
 sg13g2_tiehi _7725__298 (.L_HI(net298));
 sg13g2_tiehi _7724__299 (.L_HI(net299));
 sg13g2_tiehi _7723__300 (.L_HI(net300));
 sg13g2_tiehi _7722__301 (.L_HI(net301));
 sg13g2_tiehi _7721__302 (.L_HI(net302));
 sg13g2_tiehi _7720__303 (.L_HI(net303));
 sg13g2_tiehi _7719__304 (.L_HI(net304));
 sg13g2_tiehi _7718__305 (.L_HI(net305));
 sg13g2_tiehi _7717__306 (.L_HI(net306));
 sg13g2_tiehi _7716__307 (.L_HI(net307));
 sg13g2_tiehi _7955__308 (.L_HI(net308));
 sg13g2_tiehi _7715__309 (.L_HI(net309));
 sg13g2_tiehi _7714__310 (.L_HI(net310));
 sg13g2_tiehi _7713__311 (.L_HI(net311));
 sg13g2_tiehi _7712__312 (.L_HI(net312));
 sg13g2_tiehi _7711__313 (.L_HI(net313));
 sg13g2_tiehi _7710__314 (.L_HI(net314));
 sg13g2_tiehi _7709__315 (.L_HI(net315));
 sg13g2_tiehi _7708__316 (.L_HI(net316));
 sg13g2_tiehi _7707__317 (.L_HI(net317));
 sg13g2_tiehi _7706__318 (.L_HI(net318));
 sg13g2_tiehi _7705__319 (.L_HI(net319));
 sg13g2_tiehi _7704__320 (.L_HI(net320));
 sg13g2_tiehi _7954__321 (.L_HI(net321));
 sg13g2_tiehi _7703__322 (.L_HI(net322));
 sg13g2_tiehi _7702__323 (.L_HI(net323));
 sg13g2_tiehi _7701__324 (.L_HI(net324));
 sg13g2_tiehi _7700__325 (.L_HI(net325));
 sg13g2_tiehi _7699__326 (.L_HI(net326));
 sg13g2_tiehi _7698__327 (.L_HI(net327));
 sg13g2_tiehi _7697__328 (.L_HI(net328));
 sg13g2_tiehi _7696__329 (.L_HI(net329));
 sg13g2_tiehi _7695__330 (.L_HI(net330));
 sg13g2_tiehi _7694__331 (.L_HI(net331));
 sg13g2_tiehi _7693__332 (.L_HI(net332));
 sg13g2_tiehi _7692__333 (.L_HI(net333));
 sg13g2_tiehi _7953__334 (.L_HI(net334));
 sg13g2_tiehi _7691__335 (.L_HI(net335));
 sg13g2_tiehi _7690__336 (.L_HI(net336));
 sg13g2_tiehi _7689__337 (.L_HI(net337));
 sg13g2_tiehi _7688__338 (.L_HI(net338));
 sg13g2_tiehi _7687__339 (.L_HI(net339));
 sg13g2_tiehi _7686__340 (.L_HI(net340));
 sg13g2_tiehi _7685__341 (.L_HI(net341));
 sg13g2_tiehi _7684__342 (.L_HI(net342));
 sg13g2_tiehi _7683__343 (.L_HI(net343));
 sg13g2_tiehi _7682__344 (.L_HI(net344));
 sg13g2_tiehi _7681__345 (.L_HI(net345));
 sg13g2_tiehi _7680__346 (.L_HI(net346));
 sg13g2_tiehi _7952__347 (.L_HI(net347));
 sg13g2_tiehi _7679__348 (.L_HI(net348));
 sg13g2_tiehi _7678__349 (.L_HI(net349));
 sg13g2_tiehi _7677__350 (.L_HI(net350));
 sg13g2_tiehi _7676__351 (.L_HI(net351));
 sg13g2_tiehi _7675__352 (.L_HI(net352));
 sg13g2_tiehi _7674__353 (.L_HI(net353));
 sg13g2_tiehi _7673__354 (.L_HI(net354));
 sg13g2_tiehi _7672__355 (.L_HI(net355));
 sg13g2_tiehi _7671__356 (.L_HI(net356));
 sg13g2_tiehi _7670__357 (.L_HI(net357));
 sg13g2_tiehi _7669__358 (.L_HI(net358));
 sg13g2_tiehi _7668__359 (.L_HI(net359));
 sg13g2_tiehi _7951__360 (.L_HI(net360));
 sg13g2_tiehi _7667__361 (.L_HI(net361));
 sg13g2_tiehi _7666__362 (.L_HI(net362));
 sg13g2_tiehi _7665__363 (.L_HI(net363));
 sg13g2_tiehi _7664__364 (.L_HI(net364));
 sg13g2_tiehi _7663__365 (.L_HI(net365));
 sg13g2_tiehi _7662__366 (.L_HI(net366));
 sg13g2_tiehi _7661__367 (.L_HI(net367));
 sg13g2_tiehi heichips25_top_sorter_368 (.L_HI(net368));
 sg13g2_tiehi heichips25_top_sorter_369 (.L_HI(net369));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo heichips25_top_sorter_12 (.L_LO(net12));
 sg13g2_tielo heichips25_top_sorter_13 (.L_LO(net13));
 sg13g2_tielo heichips25_top_sorter_14 (.L_LO(net14));
 sg13g2_tielo heichips25_top_sorter_15 (.L_LO(net15));
 sg13g2_tielo heichips25_top_sorter_16 (.L_LO(net16));
 sg13g2_tielo heichips25_top_sorter_17 (.L_LO(net17));
 sg13g2_tielo heichips25_top_sorter_18 (.L_LO(net18));
 sg13g2_tielo heichips25_top_sorter_19 (.L_LO(net19));
 sg13g2_tielo heichips25_top_sorter_20 (.L_LO(net20));
 sg13g2_tielo heichips25_top_sorter_21 (.L_LO(net21));
 sg13g2_tielo heichips25_top_sorter_22 (.L_LO(net22));
 sg13g2_tielo heichips25_top_sorter_23 (.L_LO(net23));
 sg13g2_tiehi _7660__24 (.L_HI(net24));
 sg13g2_buf_1 _8333_ (.A(\s0.was_valid_out[27] [0]),
    .X(net2));
 sg13g2_buf_8 fanout1158 (.A(net1159),
    .X(net1158));
 sg13g2_buf_8 fanout1159 (.A(_3544_),
    .X(net1159));
 sg13g2_buf_8 fanout1160 (.A(net1162),
    .X(net1160));
 sg13g2_buf_8 fanout1161 (.A(net1162),
    .X(net1161));
 sg13g2_buf_8 fanout1162 (.A(_3411_),
    .X(net1162));
 sg13g2_buf_8 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(net1166),
    .X(net1164));
 sg13g2_buf_8 fanout1165 (.A(net1166),
    .X(net1165));
 sg13g2_buf_1 fanout1166 (.A(_3397_),
    .X(net1166));
 sg13g2_buf_8 fanout1167 (.A(_3396_),
    .X(net1167));
 sg13g2_buf_8 fanout1168 (.A(_3396_),
    .X(net1168));
 sg13g2_buf_8 fanout1169 (.A(net1170),
    .X(net1169));
 sg13g2_buf_8 fanout1170 (.A(_3395_),
    .X(net1170));
 sg13g2_buf_8 fanout1171 (.A(net1172),
    .X(net1171));
 sg13g2_buf_8 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_8 fanout1173 (.A(_3391_),
    .X(net1173));
 sg13g2_buf_8 fanout1174 (.A(net1176),
    .X(net1174));
 sg13g2_buf_8 fanout1175 (.A(net1176),
    .X(net1175));
 sg13g2_buf_8 fanout1176 (.A(_3390_),
    .X(net1176));
 sg13g2_buf_8 fanout1177 (.A(net1179),
    .X(net1177));
 sg13g2_buf_1 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_buf_8 fanout1179 (.A(_3388_),
    .X(net1179));
 sg13g2_buf_8 fanout1180 (.A(net1182),
    .X(net1180));
 sg13g2_buf_8 fanout1181 (.A(net1182),
    .X(net1181));
 sg13g2_buf_8 fanout1182 (.A(_3387_),
    .X(net1182));
 sg13g2_buf_8 fanout1183 (.A(net1184),
    .X(net1183));
 sg13g2_buf_8 fanout1184 (.A(_3384_),
    .X(net1184));
 sg13g2_buf_8 fanout1185 (.A(net1186),
    .X(net1185));
 sg13g2_buf_2 fanout1186 (.A(net1187),
    .X(net1186));
 sg13g2_buf_2 fanout1187 (.A(_3382_),
    .X(net1187));
 sg13g2_buf_8 fanout1188 (.A(_3381_),
    .X(net1188));
 sg13g2_buf_8 fanout1189 (.A(_3380_),
    .X(net1189));
 sg13g2_buf_8 fanout1190 (.A(_3380_),
    .X(net1190));
 sg13g2_buf_8 fanout1191 (.A(net1192),
    .X(net1191));
 sg13g2_buf_8 fanout1192 (.A(_3379_),
    .X(net1192));
 sg13g2_buf_8 fanout1193 (.A(net1194),
    .X(net1193));
 sg13g2_buf_8 fanout1194 (.A(net1195),
    .X(net1194));
 sg13g2_buf_8 fanout1195 (.A(_3378_),
    .X(net1195));
 sg13g2_buf_8 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_buf_8 fanout1197 (.A(_3377_),
    .X(net1197));
 sg13g2_buf_8 fanout1198 (.A(net1199),
    .X(net1198));
 sg13g2_buf_8 fanout1199 (.A(_3375_),
    .X(net1199));
 sg13g2_buf_2 fanout1200 (.A(net1203),
    .X(net1200));
 sg13g2_buf_8 fanout1201 (.A(net1203),
    .X(net1201));
 sg13g2_buf_2 fanout1202 (.A(net1203),
    .X(net1202));
 sg13g2_buf_8 fanout1203 (.A(\s0.shift_out[0] [0]),
    .X(net1203));
 sg13g2_buf_8 fanout1204 (.A(\s0.shift_out[0] [0]),
    .X(net1204));
 sg13g2_buf_1 fanout1205 (.A(\s0.shift_out[0] [0]),
    .X(net1205));
 sg13g2_buf_8 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_8 fanout1207 (.A(\s0.valid_out[0] [0]),
    .X(net1207));
 sg13g2_buf_1 fanout1208 (.A(\s0.valid_out[0] [0]),
    .X(net1208));
 sg13g2_buf_8 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_8 fanout1210 (.A(net1211),
    .X(net1210));
 sg13g2_buf_1 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_8 fanout1212 (.A(net474),
    .X(net1212));
 sg13g2_buf_2 fanout1213 (.A(net1214),
    .X(net1213));
 sg13g2_buf_8 fanout1214 (.A(net474),
    .X(net1214));
 sg13g2_buf_8 fanout1215 (.A(net1218),
    .X(net1215));
 sg13g2_buf_1 fanout1216 (.A(net1218),
    .X(net1216));
 sg13g2_buf_8 fanout1217 (.A(net1218),
    .X(net1217));
 sg13g2_buf_2 fanout1218 (.A(\s0.valid_out[1] [0]),
    .X(net1218));
 sg13g2_buf_2 fanout1219 (.A(net1220),
    .X(net1219));
 sg13g2_buf_1 fanout1220 (.A(net1221),
    .X(net1220));
 sg13g2_buf_1 fanout1221 (.A(\s0.shift_out[2] [0]),
    .X(net1221));
 sg13g2_buf_8 fanout1222 (.A(net1225),
    .X(net1222));
 sg13g2_buf_2 fanout1223 (.A(net1225),
    .X(net1223));
 sg13g2_buf_1 fanout1224 (.A(net1225),
    .X(net1224));
 sg13g2_buf_2 fanout1225 (.A(net831),
    .X(net1225));
 sg13g2_buf_8 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_buf_8 fanout1227 (.A(net1229),
    .X(net1227));
 sg13g2_buf_8 fanout1228 (.A(net1229),
    .X(net1228));
 sg13g2_buf_8 fanout1229 (.A(\s0.valid_out[2] [0]),
    .X(net1229));
 sg13g2_buf_8 fanout1230 (.A(net1234),
    .X(net1230));
 sg13g2_buf_8 fanout1231 (.A(net1234),
    .X(net1231));
 sg13g2_buf_8 fanout1232 (.A(net1234),
    .X(net1232));
 sg13g2_buf_8 fanout1233 (.A(net1234),
    .X(net1233));
 sg13g2_buf_8 fanout1234 (.A(net806),
    .X(net1234));
 sg13g2_buf_8 fanout1235 (.A(net806),
    .X(net1235));
 sg13g2_buf_8 fanout1236 (.A(net1237),
    .X(net1236));
 sg13g2_buf_8 fanout1237 (.A(net828),
    .X(net1237));
 sg13g2_buf_8 fanout1238 (.A(net838),
    .X(net1238));
 sg13g2_buf_8 fanout1239 (.A(net458),
    .X(net1239));
 sg13g2_buf_1 fanout1240 (.A(net458),
    .X(net1240));
 sg13g2_buf_2 fanout1241 (.A(net1242),
    .X(net1241));
 sg13g2_buf_1 fanout1242 (.A(net1244),
    .X(net1242));
 sg13g2_buf_8 fanout1243 (.A(net1244),
    .X(net1243));
 sg13g2_buf_1 fanout1244 (.A(\s0.shift_out[4] [0]),
    .X(net1244));
 sg13g2_buf_8 fanout1245 (.A(net1249),
    .X(net1245));
 sg13g2_buf_1 fanout1246 (.A(net1249),
    .X(net1246));
 sg13g2_buf_8 fanout1247 (.A(net1249),
    .X(net1247));
 sg13g2_buf_1 fanout1248 (.A(net1249),
    .X(net1248));
 sg13g2_buf_2 fanout1249 (.A(\s0.valid_out[4] [0]),
    .X(net1249));
 sg13g2_buf_8 fanout1250 (.A(net1259),
    .X(net1250));
 sg13g2_buf_1 fanout1251 (.A(net1259),
    .X(net1251));
 sg13g2_buf_8 fanout1252 (.A(net1254),
    .X(net1252));
 sg13g2_buf_2 fanout1253 (.A(net1254),
    .X(net1253));
 sg13g2_buf_1 fanout1254 (.A(net1255),
    .X(net1254));
 sg13g2_buf_1 fanout1255 (.A(net1259),
    .X(net1255));
 sg13g2_buf_2 fanout1256 (.A(net1258),
    .X(net1256));
 sg13g2_buf_2 fanout1257 (.A(net1258),
    .X(net1257));
 sg13g2_buf_1 fanout1258 (.A(net1259),
    .X(net1258));
 sg13g2_buf_1 fanout1259 (.A(net829),
    .X(net1259));
 sg13g2_buf_8 fanout1260 (.A(net1262),
    .X(net1260));
 sg13g2_buf_1 fanout1261 (.A(net1262),
    .X(net1261));
 sg13g2_buf_8 fanout1262 (.A(net1264),
    .X(net1262));
 sg13g2_buf_8 fanout1263 (.A(net1264),
    .X(net1263));
 sg13g2_buf_8 fanout1264 (.A(\s0.valid_out[5] [0]),
    .X(net1264));
 sg13g2_buf_8 fanout1265 (.A(net1267),
    .X(net1265));
 sg13g2_buf_1 fanout1266 (.A(net1267),
    .X(net1266));
 sg13g2_buf_2 fanout1267 (.A(net426),
    .X(net1267));
 sg13g2_buf_8 fanout1268 (.A(net1269),
    .X(net1268));
 sg13g2_buf_1 fanout1269 (.A(net1271),
    .X(net1269));
 sg13g2_buf_8 fanout1270 (.A(net1271),
    .X(net1270));
 sg13g2_buf_1 fanout1271 (.A(\s0.shift_out[6] [0]),
    .X(net1271));
 sg13g2_buf_8 fanout1272 (.A(net1273),
    .X(net1272));
 sg13g2_buf_1 fanout1273 (.A(\s0.valid_out[6] [0]),
    .X(net1273));
 sg13g2_buf_8 fanout1274 (.A(net1275),
    .X(net1274));
 sg13g2_buf_8 fanout1275 (.A(\s0.valid_out[6] [0]),
    .X(net1275));
 sg13g2_buf_8 fanout1276 (.A(net1277),
    .X(net1276));
 sg13g2_buf_2 fanout1277 (.A(\s0.shift_out[7] [0]),
    .X(net1277));
 sg13g2_buf_8 fanout1278 (.A(\s0.shift_out[7] [0]),
    .X(net1278));
 sg13g2_buf_8 fanout1279 (.A(net1282),
    .X(net1279));
 sg13g2_buf_2 fanout1280 (.A(net1282),
    .X(net1280));
 sg13g2_buf_1 fanout1281 (.A(net1282),
    .X(net1281));
 sg13g2_buf_1 fanout1282 (.A(\s0.shift_out[7] [0]),
    .X(net1282));
 sg13g2_buf_8 fanout1283 (.A(net1286),
    .X(net1283));
 sg13g2_buf_8 fanout1284 (.A(net1286),
    .X(net1284));
 sg13g2_buf_2 fanout1285 (.A(net1286),
    .X(net1285));
 sg13g2_buf_8 fanout1286 (.A(\s0.valid_out[7] [0]),
    .X(net1286));
 sg13g2_buf_2 fanout1287 (.A(net1288),
    .X(net1287));
 sg13g2_buf_8 fanout1288 (.A(net1289),
    .X(net1288));
 sg13g2_buf_8 fanout1289 (.A(net470),
    .X(net1289));
 sg13g2_buf_8 fanout1290 (.A(net1293),
    .X(net1290));
 sg13g2_buf_8 fanout1291 (.A(net1293),
    .X(net1291));
 sg13g2_buf_1 fanout1292 (.A(net1293),
    .X(net1292));
 sg13g2_buf_2 fanout1293 (.A(net470),
    .X(net1293));
 sg13g2_buf_8 fanout1294 (.A(\s0.valid_out[8] [0]),
    .X(net1294));
 sg13g2_buf_1 fanout1295 (.A(\s0.valid_out[8] [0]),
    .X(net1295));
 sg13g2_buf_8 fanout1296 (.A(net1297),
    .X(net1296));
 sg13g2_buf_8 fanout1297 (.A(\s0.valid_out[8] [0]),
    .X(net1297));
 sg13g2_buf_2 fanout1298 (.A(net1299),
    .X(net1298));
 sg13g2_buf_8 fanout1299 (.A(net473),
    .X(net1299));
 sg13g2_buf_2 fanout1300 (.A(net1301),
    .X(net1300));
 sg13g2_buf_2 fanout1301 (.A(\s0.shift_out[9] [0]),
    .X(net1301));
 sg13g2_buf_8 fanout1302 (.A(net1305),
    .X(net1302));
 sg13g2_buf_8 fanout1303 (.A(net1304),
    .X(net1303));
 sg13g2_buf_1 fanout1304 (.A(net1305),
    .X(net1304));
 sg13g2_buf_2 fanout1305 (.A(net473),
    .X(net1305));
 sg13g2_buf_8 fanout1306 (.A(net1310),
    .X(net1306));
 sg13g2_buf_8 fanout1307 (.A(net1310),
    .X(net1307));
 sg13g2_buf_8 fanout1308 (.A(net1310),
    .X(net1308));
 sg13g2_buf_1 fanout1309 (.A(net1310),
    .X(net1309));
 sg13g2_buf_8 fanout1310 (.A(\s0.valid_out[9] [0]),
    .X(net1310));
 sg13g2_buf_2 fanout1311 (.A(net1312),
    .X(net1311));
 sg13g2_buf_8 fanout1312 (.A(net1319),
    .X(net1312));
 sg13g2_buf_2 fanout1313 (.A(net1314),
    .X(net1313));
 sg13g2_buf_1 fanout1314 (.A(net1319),
    .X(net1314));
 sg13g2_buf_8 fanout1315 (.A(net1316),
    .X(net1315));
 sg13g2_buf_1 fanout1316 (.A(net1319),
    .X(net1316));
 sg13g2_buf_2 fanout1317 (.A(net1319),
    .X(net1317));
 sg13g2_buf_1 fanout1318 (.A(net1319),
    .X(net1318));
 sg13g2_buf_2 fanout1319 (.A(\s0.shift_out[10] [0]),
    .X(net1319));
 sg13g2_buf_8 fanout1320 (.A(net1321),
    .X(net1320));
 sg13g2_buf_8 fanout1321 (.A(net1324),
    .X(net1321));
 sg13g2_buf_8 fanout1322 (.A(net1324),
    .X(net1322));
 sg13g2_buf_8 fanout1323 (.A(net1324),
    .X(net1323));
 sg13g2_buf_8 fanout1324 (.A(\s0.data_new_delayed[7] ),
    .X(net1324));
 sg13g2_buf_8 fanout1325 (.A(net1326),
    .X(net1325));
 sg13g2_buf_8 fanout1326 (.A(net1329),
    .X(net1326));
 sg13g2_buf_8 fanout1327 (.A(net1329),
    .X(net1327));
 sg13g2_buf_8 fanout1328 (.A(net1329),
    .X(net1328));
 sg13g2_buf_8 fanout1329 (.A(\s0.data_new_delayed[6] ),
    .X(net1329));
 sg13g2_buf_8 fanout1330 (.A(net1331),
    .X(net1330));
 sg13g2_buf_8 fanout1331 (.A(net1334),
    .X(net1331));
 sg13g2_buf_8 fanout1332 (.A(net1334),
    .X(net1332));
 sg13g2_buf_8 fanout1333 (.A(net1334),
    .X(net1333));
 sg13g2_buf_8 fanout1334 (.A(\s0.data_new_delayed[5] ),
    .X(net1334));
 sg13g2_buf_8 fanout1335 (.A(net1336),
    .X(net1335));
 sg13g2_buf_8 fanout1336 (.A(net832),
    .X(net1336));
 sg13g2_buf_8 fanout1337 (.A(net1338),
    .X(net1337));
 sg13g2_buf_8 fanout1338 (.A(\s0.data_new_delayed[4] ),
    .X(net1338));
 sg13g2_buf_8 fanout1339 (.A(\s0.data_new_delayed[3] ),
    .X(net1339));
 sg13g2_buf_8 fanout1340 (.A(net1341),
    .X(net1340));
 sg13g2_buf_8 fanout1341 (.A(net830),
    .X(net1341));
 sg13g2_buf_8 fanout1342 (.A(net1343),
    .X(net1342));
 sg13g2_buf_8 fanout1343 (.A(\s0.data_new_delayed[2] ),
    .X(net1343));
 sg13g2_buf_8 fanout1344 (.A(net1345),
    .X(net1344));
 sg13g2_buf_8 fanout1345 (.A(\s0.data_new_delayed[1] ),
    .X(net1345));
 sg13g2_buf_8 fanout1346 (.A(net1347),
    .X(net1346));
 sg13g2_buf_8 fanout1347 (.A(\s0.data_new_delayed[1] ),
    .X(net1347));
 sg13g2_buf_8 fanout1348 (.A(net1349),
    .X(net1348));
 sg13g2_buf_8 fanout1349 (.A(net834),
    .X(net1349));
 sg13g2_buf_8 fanout1350 (.A(net1351),
    .X(net1350));
 sg13g2_buf_8 fanout1351 (.A(\s0.data_new_delayed[0] ),
    .X(net1351));
 sg13g2_buf_8 fanout1352 (.A(net1356),
    .X(net1352));
 sg13g2_buf_2 fanout1353 (.A(net1356),
    .X(net1353));
 sg13g2_buf_8 fanout1354 (.A(net1356),
    .X(net1354));
 sg13g2_buf_1 fanout1355 (.A(net1356),
    .X(net1355));
 sg13g2_buf_8 fanout1356 (.A(\s0.valid_out[10] [0]),
    .X(net1356));
 sg13g2_buf_8 fanout1357 (.A(net1358),
    .X(net1357));
 sg13g2_buf_8 fanout1358 (.A(net1359),
    .X(net1358));
 sg13g2_buf_8 fanout1359 (.A(\s0.shift_out[11] [0]),
    .X(net1359));
 sg13g2_buf_8 fanout1360 (.A(net1363),
    .X(net1360));
 sg13g2_buf_1 fanout1361 (.A(net1363),
    .X(net1361));
 sg13g2_buf_8 fanout1362 (.A(net1363),
    .X(net1362));
 sg13g2_buf_8 fanout1363 (.A(\s0.shift_out[11] [0]),
    .X(net1363));
 sg13g2_buf_8 fanout1364 (.A(net1365),
    .X(net1364));
 sg13g2_buf_8 fanout1365 (.A(\s0.valid_out[11] [0]),
    .X(net1365));
 sg13g2_buf_8 fanout1366 (.A(\s0.valid_out[11] [0]),
    .X(net1366));
 sg13g2_buf_8 fanout1367 (.A(\s0.valid_out[11] [0]),
    .X(net1367));
 sg13g2_buf_8 fanout1368 (.A(net1370),
    .X(net1368));
 sg13g2_buf_8 fanout1369 (.A(net1370),
    .X(net1369));
 sg13g2_buf_2 fanout1370 (.A(net1371),
    .X(net1370));
 sg13g2_buf_1 fanout1371 (.A(net1372),
    .X(net1371));
 sg13g2_buf_1 fanout1372 (.A(net1377),
    .X(net1372));
 sg13g2_buf_8 fanout1373 (.A(net1377),
    .X(net1373));
 sg13g2_buf_1 fanout1374 (.A(net1377),
    .X(net1374));
 sg13g2_buf_8 fanout1375 (.A(net1376),
    .X(net1375));
 sg13g2_buf_8 fanout1376 (.A(net1377),
    .X(net1376));
 sg13g2_buf_2 fanout1377 (.A(\s0.shift_out[12] [0]),
    .X(net1377));
 sg13g2_buf_8 fanout1378 (.A(net1379),
    .X(net1378));
 sg13g2_buf_1 fanout1379 (.A(\s0.valid_out[12] [0]),
    .X(net1379));
 sg13g2_buf_8 fanout1380 (.A(\s0.valid_out[12] [0]),
    .X(net1380));
 sg13g2_buf_8 fanout1381 (.A(\s0.valid_out[12] [0]),
    .X(net1381));
 sg13g2_buf_8 fanout1382 (.A(net1383),
    .X(net1382));
 sg13g2_buf_8 fanout1383 (.A(net1386),
    .X(net1383));
 sg13g2_buf_8 fanout1384 (.A(net1386),
    .X(net1384));
 sg13g2_buf_1 fanout1385 (.A(net1386),
    .X(net1385));
 sg13g2_buf_2 fanout1386 (.A(\s0.shift_out[13] [0]),
    .X(net1386));
 sg13g2_buf_8 fanout1387 (.A(net1388),
    .X(net1387));
 sg13g2_buf_2 fanout1388 (.A(\s0.shift_out[13] [0]),
    .X(net1388));
 sg13g2_buf_8 fanout1389 (.A(net1390),
    .X(net1389));
 sg13g2_buf_8 fanout1390 (.A(net1392),
    .X(net1390));
 sg13g2_buf_8 fanout1391 (.A(net1392),
    .X(net1391));
 sg13g2_buf_8 fanout1392 (.A(net833),
    .X(net1392));
 sg13g2_buf_8 fanout1393 (.A(net1394),
    .X(net1393));
 sg13g2_buf_8 fanout1394 (.A(net1395),
    .X(net1394));
 sg13g2_buf_8 fanout1395 (.A(net444),
    .X(net1395));
 sg13g2_buf_8 fanout1396 (.A(net1399),
    .X(net1396));
 sg13g2_buf_8 fanout1397 (.A(net1398),
    .X(net1397));
 sg13g2_buf_8 fanout1398 (.A(net1399),
    .X(net1398));
 sg13g2_buf_8 fanout1399 (.A(net444),
    .X(net1399));
 sg13g2_buf_8 fanout1400 (.A(net1401),
    .X(net1400));
 sg13g2_buf_8 fanout1401 (.A(\s0.valid_out[14] [0]),
    .X(net1401));
 sg13g2_buf_8 fanout1402 (.A(net1403),
    .X(net1402));
 sg13g2_buf_8 fanout1403 (.A(\s0.valid_out[14] [0]),
    .X(net1403));
 sg13g2_buf_8 fanout1404 (.A(net1405),
    .X(net1404));
 sg13g2_buf_8 fanout1405 (.A(net1406),
    .X(net1405));
 sg13g2_buf_1 fanout1406 (.A(net1410),
    .X(net1406));
 sg13g2_buf_2 fanout1407 (.A(net1408),
    .X(net1407));
 sg13g2_buf_8 fanout1408 (.A(net1410),
    .X(net1408));
 sg13g2_buf_8 fanout1409 (.A(net1410),
    .X(net1409));
 sg13g2_buf_8 fanout1410 (.A(net505),
    .X(net1410));
 sg13g2_buf_8 fanout1411 (.A(net1412),
    .X(net1411));
 sg13g2_buf_2 fanout1412 (.A(\s0.valid_out[15] [0]),
    .X(net1412));
 sg13g2_buf_8 fanout1413 (.A(net1414),
    .X(net1413));
 sg13g2_buf_8 fanout1414 (.A(\s0.valid_out[15] [0]),
    .X(net1414));
 sg13g2_buf_8 fanout1415 (.A(net1418),
    .X(net1415));
 sg13g2_buf_1 fanout1416 (.A(net1418),
    .X(net1416));
 sg13g2_buf_8 fanout1417 (.A(net1418),
    .X(net1417));
 sg13g2_buf_8 fanout1418 (.A(net1423),
    .X(net1418));
 sg13g2_buf_8 fanout1419 (.A(net1423),
    .X(net1419));
 sg13g2_buf_1 fanout1420 (.A(net1423),
    .X(net1420));
 sg13g2_buf_8 fanout1421 (.A(net1422),
    .X(net1421));
 sg13g2_buf_8 fanout1422 (.A(net1423),
    .X(net1422));
 sg13g2_buf_8 fanout1423 (.A(\s0.shift_out[16] [0]),
    .X(net1423));
 sg13g2_buf_8 fanout1424 (.A(net1427),
    .X(net1424));
 sg13g2_buf_8 fanout1425 (.A(net1426),
    .X(net1425));
 sg13g2_buf_8 fanout1426 (.A(net1427),
    .X(net1426));
 sg13g2_buf_8 fanout1427 (.A(\s0.valid_out[16] [0]),
    .X(net1427));
 sg13g2_buf_8 fanout1428 (.A(net1429),
    .X(net1428));
 sg13g2_buf_1 fanout1429 (.A(net1430),
    .X(net1429));
 sg13g2_buf_2 fanout1430 (.A(net481),
    .X(net1430));
 sg13g2_buf_8 fanout1431 (.A(net1434),
    .X(net1431));
 sg13g2_buf_8 fanout1432 (.A(net1434),
    .X(net1432));
 sg13g2_buf_1 fanout1433 (.A(net1434),
    .X(net1433));
 sg13g2_buf_8 fanout1434 (.A(net481),
    .X(net1434));
 sg13g2_buf_8 fanout1435 (.A(net1439),
    .X(net1435));
 sg13g2_buf_8 fanout1436 (.A(net1438),
    .X(net1436));
 sg13g2_buf_1 fanout1437 (.A(net1438),
    .X(net1437));
 sg13g2_buf_8 fanout1438 (.A(net1439),
    .X(net1438));
 sg13g2_buf_8 fanout1439 (.A(\s0.valid_out[17] [0]),
    .X(net1439));
 sg13g2_buf_8 fanout1440 (.A(net1441),
    .X(net1440));
 sg13g2_buf_8 fanout1441 (.A(net1443),
    .X(net1441));
 sg13g2_buf_8 fanout1442 (.A(net1443),
    .X(net1442));
 sg13g2_buf_8 fanout1443 (.A(net1446),
    .X(net1443));
 sg13g2_buf_8 fanout1444 (.A(net1445),
    .X(net1444));
 sg13g2_buf_8 fanout1445 (.A(net1446),
    .X(net1445));
 sg13g2_buf_8 fanout1446 (.A(net403),
    .X(net1446));
 sg13g2_buf_8 fanout1447 (.A(net1450),
    .X(net1447));
 sg13g2_buf_8 fanout1448 (.A(net1450),
    .X(net1448));
 sg13g2_buf_8 fanout1449 (.A(net1450),
    .X(net1449));
 sg13g2_buf_8 fanout1450 (.A(\s0.valid_out[18] [0]),
    .X(net1450));
 sg13g2_buf_8 fanout1451 (.A(\s0.shift_out[19] [0]),
    .X(net1451));
 sg13g2_buf_1 fanout1452 (.A(net1453),
    .X(net1452));
 sg13g2_buf_8 fanout1453 (.A(\s0.shift_out[19] [0]),
    .X(net1453));
 sg13g2_buf_8 fanout1454 (.A(net1455),
    .X(net1454));
 sg13g2_buf_8 fanout1455 (.A(net1456),
    .X(net1455));
 sg13g2_buf_8 fanout1456 (.A(\s0.shift_out[19] [0]),
    .X(net1456));
 sg13g2_buf_8 fanout1457 (.A(\s0.valid_out[19] [0]),
    .X(net1457));
 sg13g2_buf_1 fanout1458 (.A(\s0.valid_out[19] [0]),
    .X(net1458));
 sg13g2_buf_8 fanout1459 (.A(net1460),
    .X(net1459));
 sg13g2_buf_8 fanout1460 (.A(\s0.valid_out[19] [0]),
    .X(net1460));
 sg13g2_buf_8 fanout1461 (.A(net1462),
    .X(net1461));
 sg13g2_buf_8 fanout1462 (.A(net1469),
    .X(net1462));
 sg13g2_buf_2 fanout1463 (.A(net1464),
    .X(net1463));
 sg13g2_buf_1 fanout1464 (.A(net1465),
    .X(net1464));
 sg13g2_buf_2 fanout1465 (.A(net1469),
    .X(net1465));
 sg13g2_buf_8 fanout1466 (.A(net1468),
    .X(net1466));
 sg13g2_buf_1 fanout1467 (.A(net1468),
    .X(net1467));
 sg13g2_buf_8 fanout1468 (.A(net1469),
    .X(net1468));
 sg13g2_buf_8 fanout1469 (.A(net408),
    .X(net1469));
 sg13g2_buf_8 fanout1470 (.A(net1473),
    .X(net1470));
 sg13g2_buf_8 fanout1471 (.A(net1473),
    .X(net1471));
 sg13g2_buf_8 fanout1472 (.A(net1473),
    .X(net1472));
 sg13g2_buf_8 fanout1473 (.A(\s0.valid_out[20] [0]),
    .X(net1473));
 sg13g2_buf_2 fanout1474 (.A(net1477),
    .X(net1474));
 sg13g2_buf_8 fanout1475 (.A(net1477),
    .X(net1475));
 sg13g2_buf_1 fanout1476 (.A(net1477),
    .X(net1476));
 sg13g2_buf_2 fanout1477 (.A(net734),
    .X(net1477));
 sg13g2_buf_2 fanout1478 (.A(net1479),
    .X(net1478));
 sg13g2_buf_1 fanout1479 (.A(net1480),
    .X(net1479));
 sg13g2_buf_1 fanout1480 (.A(net1481),
    .X(net1480));
 sg13g2_buf_1 fanout1481 (.A(\s0.shift_out[21] [0]),
    .X(net1481));
 sg13g2_buf_8 fanout1482 (.A(net1483),
    .X(net1482));
 sg13g2_buf_8 fanout1483 (.A(net1485),
    .X(net1483));
 sg13g2_buf_8 fanout1484 (.A(net1485),
    .X(net1484));
 sg13g2_buf_8 fanout1485 (.A(\s0.valid_out[21] [0]),
    .X(net1485));
 sg13g2_buf_8 fanout1486 (.A(net1494),
    .X(net1486));
 sg13g2_buf_1 fanout1487 (.A(net1494),
    .X(net1487));
 sg13g2_buf_2 fanout1488 (.A(net1489),
    .X(net1488));
 sg13g2_buf_1 fanout1489 (.A(net1494),
    .X(net1489));
 sg13g2_buf_8 fanout1490 (.A(net1491),
    .X(net1490));
 sg13g2_buf_8 fanout1491 (.A(net1494),
    .X(net1491));
 sg13g2_buf_8 fanout1492 (.A(net1493),
    .X(net1492));
 sg13g2_buf_2 fanout1493 (.A(net1494),
    .X(net1493));
 sg13g2_buf_8 fanout1494 (.A(net413),
    .X(net1494));
 sg13g2_buf_8 fanout1495 (.A(\s0.valid_out[22] [0]),
    .X(net1495));
 sg13g2_buf_2 fanout1496 (.A(\s0.valid_out[22] [0]),
    .X(net1496));
 sg13g2_buf_8 fanout1497 (.A(net1498),
    .X(net1497));
 sg13g2_buf_8 fanout1498 (.A(\s0.valid_out[22] [0]),
    .X(net1498));
 sg13g2_buf_8 fanout1499 (.A(net1502),
    .X(net1499));
 sg13g2_buf_1 fanout1500 (.A(net1502),
    .X(net1500));
 sg13g2_buf_8 fanout1501 (.A(net1502),
    .X(net1501));
 sg13g2_buf_2 fanout1502 (.A(net1505),
    .X(net1502));
 sg13g2_buf_8 fanout1503 (.A(net1504),
    .X(net1503));
 sg13g2_buf_8 fanout1504 (.A(net1505),
    .X(net1504));
 sg13g2_buf_1 fanout1505 (.A(\s0.shift_out[23] [0]),
    .X(net1505));
 sg13g2_buf_8 fanout1506 (.A(net1507),
    .X(net1506));
 sg13g2_buf_8 fanout1507 (.A(\s0.valid_out[23] [0]),
    .X(net1507));
 sg13g2_buf_8 fanout1508 (.A(\s0.valid_out[23] [0]),
    .X(net1508));
 sg13g2_buf_2 fanout1509 (.A(net1517),
    .X(net1509));
 sg13g2_buf_1 fanout1510 (.A(net1517),
    .X(net1510));
 sg13g2_buf_2 fanout1511 (.A(net1512),
    .X(net1511));
 sg13g2_buf_1 fanout1512 (.A(net1517),
    .X(net1512));
 sg13g2_buf_8 fanout1513 (.A(net1514),
    .X(net1513));
 sg13g2_buf_8 fanout1514 (.A(net1517),
    .X(net1514));
 sg13g2_buf_8 fanout1515 (.A(net1517),
    .X(net1515));
 sg13g2_buf_1 fanout1516 (.A(net1517),
    .X(net1516));
 sg13g2_buf_8 fanout1517 (.A(\s0.shift_out[24] [0]),
    .X(net1517));
 sg13g2_buf_8 fanout1518 (.A(net1522),
    .X(net1518));
 sg13g2_buf_1 fanout1519 (.A(net1522),
    .X(net1519));
 sg13g2_buf_2 fanout1520 (.A(net1522),
    .X(net1520));
 sg13g2_buf_1 fanout1521 (.A(net1522),
    .X(net1521));
 sg13g2_buf_1 fanout1522 (.A(\s0.valid_out[24] [0]),
    .X(net1522));
 sg13g2_buf_2 fanout1523 (.A(net1526),
    .X(net1523));
 sg13g2_buf_1 fanout1524 (.A(net1526),
    .X(net1524));
 sg13g2_buf_8 fanout1525 (.A(net1526),
    .X(net1525));
 sg13g2_buf_2 fanout1526 (.A(net1529),
    .X(net1526));
 sg13g2_buf_8 fanout1527 (.A(net1528),
    .X(net1527));
 sg13g2_buf_8 fanout1528 (.A(net1529),
    .X(net1528));
 sg13g2_buf_1 fanout1529 (.A(\s0.shift_out[25] [0]),
    .X(net1529));
 sg13g2_buf_8 fanout1530 (.A(net1534),
    .X(net1530));
 sg13g2_buf_8 fanout1531 (.A(net1534),
    .X(net1531));
 sg13g2_buf_8 fanout1532 (.A(net1534),
    .X(net1532));
 sg13g2_buf_1 fanout1533 (.A(net1534),
    .X(net1533));
 sg13g2_buf_8 fanout1534 (.A(\s0.valid_out[25] [0]),
    .X(net1534));
 sg13g2_buf_8 fanout1535 (.A(net1539),
    .X(net1535));
 sg13g2_buf_1 fanout1536 (.A(net1539),
    .X(net1536));
 sg13g2_buf_8 fanout1537 (.A(net1539),
    .X(net1537));
 sg13g2_buf_1 fanout1538 (.A(net1539),
    .X(net1538));
 sg13g2_buf_2 fanout1539 (.A(\s0.shift_out[26] [0]),
    .X(net1539));
 sg13g2_buf_8 fanout1540 (.A(net1544),
    .X(net1540));
 sg13g2_buf_1 fanout1541 (.A(net1544),
    .X(net1541));
 sg13g2_buf_8 fanout1542 (.A(net1544),
    .X(net1542));
 sg13g2_buf_1 fanout1543 (.A(net1544),
    .X(net1543));
 sg13g2_buf_2 fanout1544 (.A(\s0.shift_out[26] [0]),
    .X(net1544));
 sg13g2_buf_8 fanout1545 (.A(\s0.valid_out[26] [0]),
    .X(net1545));
 sg13g2_buf_1 fanout1546 (.A(\s0.valid_out[26] [0]),
    .X(net1546));
 sg13g2_buf_8 fanout1547 (.A(net1548),
    .X(net1547));
 sg13g2_buf_8 fanout1548 (.A(\s0.valid_out[26] [0]),
    .X(net1548));
 sg13g2_buf_8 fanout1549 (.A(net1550),
    .X(net1549));
 sg13g2_buf_8 fanout1550 (.A(net1552),
    .X(net1550));
 sg13g2_buf_8 fanout1551 (.A(net1552),
    .X(net1551));
 sg13g2_buf_8 fanout1552 (.A(\s0.shift_out[27] [0]),
    .X(net1552));
 sg13g2_buf_8 fanout1553 (.A(net1554),
    .X(net1553));
 sg13g2_buf_8 fanout1554 (.A(net454),
    .X(net1554));
 sg13g2_buf_8 fanout1555 (.A(_0349_),
    .X(net1555));
 sg13g2_buf_8 fanout1556 (.A(_0349_),
    .X(net1556));
 sg13g2_buf_8 fanout1557 (.A(net1558),
    .X(net1557));
 sg13g2_buf_8 fanout1558 (.A(_0349_),
    .X(net1558));
 sg13g2_buf_8 fanout1559 (.A(_3418_),
    .X(net1559));
 sg13g2_buf_8 fanout1560 (.A(net1563),
    .X(net1560));
 sg13g2_buf_2 fanout1561 (.A(net1563),
    .X(net1561));
 sg13g2_buf_8 fanout1562 (.A(net1563),
    .X(net1562));
 sg13g2_buf_8 fanout1563 (.A(_3414_),
    .X(net1563));
 sg13g2_buf_8 fanout1564 (.A(net1565),
    .X(net1564));
 sg13g2_buf_8 fanout1565 (.A(net1567),
    .X(net1565));
 sg13g2_buf_8 fanout1566 (.A(net1567),
    .X(net1566));
 sg13g2_buf_2 fanout1567 (.A(net1577),
    .X(net1567));
 sg13g2_buf_8 fanout1568 (.A(net1570),
    .X(net1568));
 sg13g2_buf_1 fanout1569 (.A(net1570),
    .X(net1569));
 sg13g2_buf_8 fanout1570 (.A(net1577),
    .X(net1570));
 sg13g2_buf_8 fanout1571 (.A(net1572),
    .X(net1571));
 sg13g2_buf_8 fanout1572 (.A(net1576),
    .X(net1572));
 sg13g2_buf_8 fanout1573 (.A(net1574),
    .X(net1573));
 sg13g2_buf_8 fanout1574 (.A(net1575),
    .X(net1574));
 sg13g2_buf_8 fanout1575 (.A(net1576),
    .X(net1575));
 sg13g2_buf_8 fanout1576 (.A(net1577),
    .X(net1576));
 sg13g2_buf_8 fanout1577 (.A(net1620),
    .X(net1577));
 sg13g2_buf_8 fanout1578 (.A(net1579),
    .X(net1578));
 sg13g2_buf_8 fanout1579 (.A(net1583),
    .X(net1579));
 sg13g2_buf_8 fanout1580 (.A(net1582),
    .X(net1580));
 sg13g2_buf_1 fanout1581 (.A(net1582),
    .X(net1581));
 sg13g2_buf_8 fanout1582 (.A(net1583),
    .X(net1582));
 sg13g2_buf_8 fanout1583 (.A(net1620),
    .X(net1583));
 sg13g2_buf_8 fanout1584 (.A(net1586),
    .X(net1584));
 sg13g2_buf_8 fanout1585 (.A(net1586),
    .X(net1585));
 sg13g2_buf_8 fanout1586 (.A(net1591),
    .X(net1586));
 sg13g2_buf_8 fanout1587 (.A(net1591),
    .X(net1587));
 sg13g2_buf_1 fanout1588 (.A(net1591),
    .X(net1588));
 sg13g2_buf_8 fanout1589 (.A(net1590),
    .X(net1589));
 sg13g2_buf_8 fanout1590 (.A(net1591),
    .X(net1590));
 sg13g2_buf_8 fanout1591 (.A(net1620),
    .X(net1591));
 sg13g2_buf_8 fanout1592 (.A(net1593),
    .X(net1592));
 sg13g2_buf_8 fanout1593 (.A(net1604),
    .X(net1593));
 sg13g2_buf_8 fanout1594 (.A(net1604),
    .X(net1594));
 sg13g2_buf_1 fanout1595 (.A(net1604),
    .X(net1595));
 sg13g2_buf_8 fanout1596 (.A(net1598),
    .X(net1596));
 sg13g2_buf_1 fanout1597 (.A(net1598),
    .X(net1597));
 sg13g2_buf_8 fanout1598 (.A(net1603),
    .X(net1598));
 sg13g2_buf_8 fanout1599 (.A(net1602),
    .X(net1599));
 sg13g2_buf_1 fanout1600 (.A(net1602),
    .X(net1600));
 sg13g2_buf_8 fanout1601 (.A(net1602),
    .X(net1601));
 sg13g2_buf_8 fanout1602 (.A(net1603),
    .X(net1602));
 sg13g2_buf_8 fanout1603 (.A(net1604),
    .X(net1603));
 sg13g2_buf_8 fanout1604 (.A(net1620),
    .X(net1604));
 sg13g2_buf_8 fanout1605 (.A(net1612),
    .X(net1605));
 sg13g2_buf_2 fanout1606 (.A(net1612),
    .X(net1606));
 sg13g2_buf_8 fanout1607 (.A(net1608),
    .X(net1607));
 sg13g2_buf_8 fanout1608 (.A(net1612),
    .X(net1608));
 sg13g2_buf_8 fanout1609 (.A(net1611),
    .X(net1609));
 sg13g2_buf_8 fanout1610 (.A(net1611),
    .X(net1610));
 sg13g2_buf_8 fanout1611 (.A(net1612),
    .X(net1611));
 sg13g2_buf_8 fanout1612 (.A(net1620),
    .X(net1612));
 sg13g2_buf_8 fanout1613 (.A(net1614),
    .X(net1613));
 sg13g2_buf_8 fanout1614 (.A(net1616),
    .X(net1614));
 sg13g2_buf_8 fanout1615 (.A(net1616),
    .X(net1615));
 sg13g2_buf_8 fanout1616 (.A(net1619),
    .X(net1616));
 sg13g2_buf_8 fanout1617 (.A(net1618),
    .X(net1617));
 sg13g2_buf_8 fanout1618 (.A(net1619),
    .X(net1618));
 sg13g2_buf_8 fanout1619 (.A(net1620),
    .X(net1619));
 sg13g2_buf_8 fanout1620 (.A(_3374_),
    .X(net1620));
 sg13g2_buf_8 fanout1621 (.A(net1624),
    .X(net1621));
 sg13g2_buf_8 fanout1622 (.A(net1624),
    .X(net1622));
 sg13g2_buf_8 fanout1623 (.A(net1624),
    .X(net1623));
 sg13g2_buf_8 fanout1624 (.A(_3373_),
    .X(net1624));
 sg13g2_buf_8 fanout1625 (.A(net1626),
    .X(net1625));
 sg13g2_buf_8 fanout1626 (.A(net1),
    .X(net1626));
 sg13g2_buf_8 fanout1627 (.A(net1629),
    .X(net1627));
 sg13g2_buf_8 fanout1628 (.A(net1629),
    .X(net1628));
 sg13g2_buf_8 fanout1629 (.A(net1634),
    .X(net1629));
 sg13g2_buf_8 fanout1630 (.A(net1633),
    .X(net1630));
 sg13g2_buf_1 fanout1631 (.A(net1633),
    .X(net1631));
 sg13g2_buf_8 fanout1632 (.A(net1633),
    .X(net1632));
 sg13g2_buf_8 fanout1633 (.A(net1634),
    .X(net1633));
 sg13g2_buf_8 fanout1634 (.A(uio_in[0]),
    .X(net1634));
 sg13g2_buf_8 fanout1635 (.A(net1636),
    .X(net1635));
 sg13g2_buf_8 fanout1636 (.A(net1640),
    .X(net1636));
 sg13g2_buf_8 fanout1637 (.A(net1640),
    .X(net1637));
 sg13g2_buf_8 fanout1638 (.A(net1640),
    .X(net1638));
 sg13g2_buf_1 fanout1639 (.A(net1640),
    .X(net1639));
 sg13g2_buf_8 fanout1640 (.A(ui_in[7]),
    .X(net1640));
 sg13g2_buf_8 fanout1641 (.A(net1645),
    .X(net1641));
 sg13g2_buf_8 fanout1642 (.A(net1644),
    .X(net1642));
 sg13g2_buf_8 fanout1643 (.A(net1645),
    .X(net1643));
 sg13g2_buf_1 fanout1644 (.A(net1645),
    .X(net1644));
 sg13g2_buf_8 fanout1645 (.A(ui_in[7]),
    .X(net1645));
 sg13g2_buf_8 fanout1646 (.A(net1650),
    .X(net1646));
 sg13g2_buf_8 fanout1647 (.A(net1650),
    .X(net1647));
 sg13g2_buf_8 fanout1648 (.A(net1650),
    .X(net1648));
 sg13g2_buf_1 fanout1649 (.A(net1650),
    .X(net1649));
 sg13g2_buf_8 fanout1650 (.A(ui_in[6]),
    .X(net1650));
 sg13g2_buf_8 fanout1651 (.A(net1654),
    .X(net1651));
 sg13g2_buf_8 fanout1652 (.A(net1654),
    .X(net1652));
 sg13g2_buf_8 fanout1653 (.A(net1654),
    .X(net1653));
 sg13g2_buf_8 fanout1654 (.A(ui_in[6]),
    .X(net1654));
 sg13g2_buf_8 fanout1655 (.A(net1659),
    .X(net1655));
 sg13g2_buf_1 fanout1656 (.A(net1659),
    .X(net1656));
 sg13g2_buf_8 fanout1657 (.A(net1659),
    .X(net1657));
 sg13g2_buf_8 fanout1658 (.A(net1659),
    .X(net1658));
 sg13g2_buf_8 fanout1659 (.A(ui_in[5]),
    .X(net1659));
 sg13g2_buf_8 fanout1660 (.A(net1664),
    .X(net1660));
 sg13g2_buf_8 fanout1661 (.A(net1663),
    .X(net1661));
 sg13g2_buf_8 fanout1662 (.A(net1663),
    .X(net1662));
 sg13g2_buf_8 fanout1663 (.A(net1664),
    .X(net1663));
 sg13g2_buf_8 fanout1664 (.A(ui_in[5]),
    .X(net1664));
 sg13g2_buf_8 fanout1665 (.A(net1669),
    .X(net1665));
 sg13g2_buf_1 fanout1666 (.A(net1669),
    .X(net1666));
 sg13g2_buf_8 fanout1667 (.A(net1669),
    .X(net1667));
 sg13g2_buf_2 fanout1668 (.A(net1669),
    .X(net1668));
 sg13g2_buf_8 fanout1669 (.A(ui_in[4]),
    .X(net1669));
 sg13g2_buf_8 fanout1670 (.A(net1673),
    .X(net1670));
 sg13g2_buf_8 fanout1671 (.A(net1672),
    .X(net1671));
 sg13g2_buf_8 fanout1672 (.A(net1673),
    .X(net1672));
 sg13g2_buf_8 fanout1673 (.A(ui_in[4]),
    .X(net1673));
 sg13g2_buf_8 fanout1674 (.A(net1675),
    .X(net1674));
 sg13g2_buf_8 fanout1675 (.A(net1677),
    .X(net1675));
 sg13g2_buf_8 fanout1676 (.A(net1677),
    .X(net1676));
 sg13g2_buf_8 fanout1677 (.A(net1683),
    .X(net1677));
 sg13g2_buf_8 fanout1678 (.A(net1683),
    .X(net1678));
 sg13g2_buf_2 fanout1679 (.A(net1683),
    .X(net1679));
 sg13g2_buf_8 fanout1680 (.A(net1682),
    .X(net1680));
 sg13g2_buf_8 fanout1681 (.A(net1682),
    .X(net1681));
 sg13g2_buf_8 fanout1682 (.A(net1683),
    .X(net1682));
 sg13g2_buf_8 fanout1683 (.A(ui_in[3]),
    .X(net1683));
 sg13g2_buf_8 fanout1684 (.A(net1685),
    .X(net1684));
 sg13g2_buf_8 fanout1685 (.A(net1689),
    .X(net1685));
 sg13g2_buf_8 fanout1686 (.A(net1689),
    .X(net1686));
 sg13g2_buf_1 fanout1687 (.A(net1689),
    .X(net1687));
 sg13g2_buf_8 fanout1688 (.A(net1689),
    .X(net1688));
 sg13g2_buf_8 fanout1689 (.A(ui_in[2]),
    .X(net1689));
 sg13g2_buf_8 fanout1690 (.A(net1693),
    .X(net1690));
 sg13g2_buf_1 fanout1691 (.A(net1693),
    .X(net1691));
 sg13g2_buf_8 fanout1692 (.A(net1693),
    .X(net1692));
 sg13g2_buf_8 fanout1693 (.A(ui_in[1]),
    .X(net1693));
 sg13g2_buf_8 fanout1694 (.A(net1699),
    .X(net1694));
 sg13g2_buf_8 fanout1695 (.A(net1698),
    .X(net1695));
 sg13g2_buf_1 fanout1696 (.A(net1698),
    .X(net1696));
 sg13g2_buf_8 fanout1697 (.A(net1698),
    .X(net1697));
 sg13g2_buf_8 fanout1698 (.A(net1699),
    .X(net1698));
 sg13g2_buf_8 fanout1699 (.A(ui_in[1]),
    .X(net1699));
 sg13g2_buf_8 fanout1700 (.A(net1703),
    .X(net1700));
 sg13g2_buf_8 fanout1701 (.A(net1703),
    .X(net1701));
 sg13g2_buf_8 fanout1702 (.A(net1703),
    .X(net1702));
 sg13g2_buf_8 fanout1703 (.A(ui_in[0]),
    .X(net1703));
 sg13g2_buf_8 fanout1704 (.A(net1707),
    .X(net1704));
 sg13g2_buf_8 fanout1705 (.A(net1707),
    .X(net1705));
 sg13g2_buf_8 fanout1706 (.A(net1707),
    .X(net1706));
 sg13g2_buf_8 fanout1707 (.A(net1721),
    .X(net1707));
 sg13g2_buf_8 fanout1708 (.A(net1711),
    .X(net1708));
 sg13g2_buf_8 fanout1709 (.A(net1710),
    .X(net1709));
 sg13g2_buf_8 fanout1710 (.A(net1711),
    .X(net1710));
 sg13g2_buf_8 fanout1711 (.A(net1721),
    .X(net1711));
 sg13g2_buf_8 fanout1712 (.A(net1713),
    .X(net1712));
 sg13g2_buf_8 fanout1713 (.A(net1721),
    .X(net1713));
 sg13g2_buf_8 fanout1714 (.A(net1717),
    .X(net1714));
 sg13g2_buf_8 fanout1715 (.A(net1717),
    .X(net1715));
 sg13g2_buf_8 fanout1716 (.A(net1717),
    .X(net1716));
 sg13g2_buf_8 fanout1717 (.A(net1721),
    .X(net1717));
 sg13g2_buf_8 fanout1718 (.A(net1720),
    .X(net1718));
 sg13g2_buf_8 fanout1719 (.A(net1720),
    .X(net1719));
 sg13g2_buf_8 fanout1720 (.A(net1721),
    .X(net1720));
 sg13g2_buf_8 fanout1721 (.A(net1740),
    .X(net1721));
 sg13g2_buf_8 fanout1722 (.A(net1725),
    .X(net1722));
 sg13g2_buf_2 fanout1723 (.A(net1725),
    .X(net1723));
 sg13g2_buf_8 fanout1724 (.A(net1725),
    .X(net1724));
 sg13g2_buf_8 fanout1725 (.A(net1740),
    .X(net1725));
 sg13g2_buf_8 fanout1726 (.A(net1730),
    .X(net1726));
 sg13g2_buf_1 fanout1727 (.A(net1730),
    .X(net1727));
 sg13g2_buf_8 fanout1728 (.A(net1729),
    .X(net1728));
 sg13g2_buf_8 fanout1729 (.A(net1730),
    .X(net1729));
 sg13g2_buf_8 fanout1730 (.A(net1740),
    .X(net1730));
 sg13g2_buf_8 fanout1731 (.A(net1735),
    .X(net1731));
 sg13g2_buf_2 fanout1732 (.A(net1735),
    .X(net1732));
 sg13g2_buf_8 fanout1733 (.A(net1735),
    .X(net1733));
 sg13g2_buf_1 fanout1734 (.A(net1735),
    .X(net1734));
 sg13g2_buf_2 fanout1735 (.A(net1739),
    .X(net1735));
 sg13g2_buf_8 fanout1736 (.A(net1739),
    .X(net1736));
 sg13g2_buf_2 fanout1737 (.A(net1739),
    .X(net1737));
 sg13g2_buf_8 fanout1738 (.A(net1739),
    .X(net1738));
 sg13g2_buf_8 fanout1739 (.A(net1740),
    .X(net1739));
 sg13g2_buf_8 fanout1740 (.A(rst_n),
    .X(net1740));
 sg13g2_buf_1 input1 (.A(uio_in[1]),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uio_out[2]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[7]));
 sg13g2_tielo heichips25_top_sorter_11 (.L_LO(net11));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_46_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_2_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_36_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_38_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_30_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_leaf_32_clk));
 sg13g2_inv_8 clkload9 (.A(clknet_leaf_15_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_leaf_18_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_leaf_27_clk));
 sg13g2_inv_8 clkload12 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_26_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\s0.genblk1[19].modules.bubble ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold2 (.A(\s0.genblk1[26].modules.bubble ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold3 (.A(\s0.genblk1[2].modules.bubble ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold4 (.A(\s0.genblk1[10].modules.bubble ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold5 (.A(\s0.genblk1[22].modules.bubble ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold6 (.A(\s0.genblk1[13].modules.bubble ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold7 (.A(\s0.genblk1[20].modules.bubble ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold8 (.A(\s0.genblk1[3].modules.bubble ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold9 (.A(\s0.genblk1[23].modules.bubble ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold10 (.A(\s0.genblk1[25].modules.bubble ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold11 (.A(\s0.genblk1[4].modules.bubble ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold12 (.A(\s0.genblk1[18].modules.bubble ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold13 (.A(\s0.genblk1[24].modules.bubble ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold14 (.A(\s0.genblk1[27].modules.bubble ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold15 (.A(\s0.module0.bubble ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold16 (.A(\s0.genblk1[11].modules.bubble ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold17 (.A(\s0.genblk1[12].modules.bubble ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold18 (.A(\s0.genblk1[21].modules.bubble ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold19 (.A(\s0.genblk1[9].modules.bubble ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold20 (.A(\s0.genblk1[16].modules.bubble ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold21 (.A(\s0.genblk1[17].modules.bubble ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold22 (.A(\s0.genblk1[8].modules.bubble ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold23 (.A(\s0.genblk1[14].modules.bubble ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold24 (.A(\s0.genblk1[7].modules.bubble ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold25 (.A(\s0.genblk1[15].modules.bubble ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold26 (.A(\s0.genblk1[1].modules.bubble ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold27 (.A(\s0.genblk1[5].modules.bubble ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold28 (.A(\s0.genblk1[6].modules.bubble ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold29 (.A(\s0.was_valid_out[15] [0]),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0253_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold31 (.A(\s0.was_valid_out[21] [0]),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0181_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold33 (.A(\s0.data_out[10][4] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold34 (.A(\s0.shift_out[18] [0]),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold35 (.A(_1279_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold36 (.A(_1359_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold37 (.A(\s0.was_valid_out[3] [0]),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0060_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold39 (.A(\s0.shift_out[20] [0]),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold40 (.A(\s0.was_valid_out[19] [0]),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0205_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold42 (.A(\s0.was_valid_out[22] [0]),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold43 (.A(\s0.was_valid_out[23] [0]),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold44 (.A(\s0.shift_out[22] [0]),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0863_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold46 (.A(\s0.data_out[22][4] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold47 (.A(\s0.was_valid_out[4] [0]),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0048_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold49 (.A(\s0.was_valid_out[25] [0]),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0133_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold51 (.A(\s0.was_valid_out[17] [0]),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0229_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold53 (.A(\s0.was_valid_out[6] [0]),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0024_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold55 (.A(\s0.data_out[2][4] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold56 (.A(_3057_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold57 (.A(\s0.shift_out[6] [0]),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold58 (.A(_2745_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0031_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold60 (.A(\s0.data_out[24][5] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0672_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold62 (.A(\s0.data_out[0][1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold63 (.A(\s0.was_valid_out[2] [0]),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0072_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold65 (.A(\s0.was_valid_out[5] [0]),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold66 (.A(\s0.data_out[0][5] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold67 (.A(\s0.data_out[10][3] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold68 (.A(_2115_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold69 (.A(\s0.data_out[25][4] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold70 (.A(\s0.was_valid_out[13] [0]),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0277_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold72 (.A(\s0.data_out[0][3] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0103_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold74 (.A(\s0.data_out[0][4] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold75 (.A(\s0.shift_out[14] [0]),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold76 (.A(\s0.was_valid_out[11] [0]),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0301_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold78 (.A(\s0.was_valid_out[9] [0]),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0332_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold80 (.A(\s0.data_out[21][5] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold81 (.A(_1007_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold82 (.A(\s0.data_out[0][7] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold83 (.A(\s0.was_valid_out[10] [0]),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold84 (.A(\s0.data_out[12][4] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold85 (.A(\s0.valid_out[27] [0]),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold86 (.A(_3571_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold87 (.A(\s0.data_out[27][3] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0116_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold89 (.A(\s0.shift_out[4] [0]),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold90 (.A(\s0.was_valid_out[7] [0]),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold91 (.A(\s0.data_out[7][7] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold92 (.A(_2580_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold93 (.A(\s0.was_valid_out[12] [0]),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold94 (.A(\s0.data_out[27][4] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0117_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold96 (.A(\s0.data_out[16][5] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold97 (.A(_1580_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold98 (.A(\s0.data_out[27][5] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0118_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold100 (.A(\s0.data_out[0][2] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold101 (.A(\s0.shift_out[8] [0]),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold102 (.A(\s0.data_out[16][3] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0248_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold104 (.A(\s0.shift_out[9] [0]),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold105 (.A(\s0.shift_out[1] [0]),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold106 (.A(\s0.data_out[9][1] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0337_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold108 (.A(\s0.data_out[26][2] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0127_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold110 (.A(\s0.data_out[10][2] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0326_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold112 (.A(\s0.shift_out[17] [0]),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold113 (.A(\s0.data_out[18][3] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0224_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold115 (.A(\s0.data_out[16][1] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0246_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold117 (.A(\s0.data_out[27][6] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0119_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold119 (.A(\s0.data_out[22][6] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0179_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold121 (.A(\s0.data_out[9][2] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0338_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold123 (.A(\s0.data_out[20][5] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0202_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold125 (.A(\s0.data_out[0][6] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold126 (.A(\s0.data_out[4][3] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold127 (.A(_2798_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold128 (.A(\s0.data_out[10][5] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0329_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold130 (.A(\s0.data_out[21][3] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0187_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold132 (.A(\s0.data_out[3][3] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold133 (.A(\s0.data_out[24][3] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0152_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold135 (.A(\s0.was_valid_out[0] [0]),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold136 (.A(\s0.shift_out[15] [0]),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold137 (.A(\s0.was_valid_out[26] [0]),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold138 (.A(\s0.data_out[27][2] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0115_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold140 (.A(\s0.data_out[24][1] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0150_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold142 (.A(\s0.data_out[26][4] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold143 (.A(\s0.data_out[26][5] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0130_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold145 (.A(\s0.data_out[10][7] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0331_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold147 (.A(\s0.data_out[20][4] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0201_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold149 (.A(\s0.data_out[13][4] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0285_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold151 (.A(\s0.data_out[21][2] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold152 (.A(_1040_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold153 (.A(\s0.data_out[12][7] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0300_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold155 (.A(\s0.data_out[27][0] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0113_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold157 (.A(\s0.data_out[22][7] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0180_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold159 (.A(\s0.data_out[5][7] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0047_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold161 (.A(\s0.data_out[17][2] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold162 (.A(_1489_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold163 (.A(\s0.data_out[14][4] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold164 (.A(_1837_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold165 (.A(\s0.data_out[9][7] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0343_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold167 (.A(\s0.data_out[26][7] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0132_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold169 (.A(\s0.data_out[16][7] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0252_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold171 (.A(\s0.data_out[24][7] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0156_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold173 (.A(\s0.data_out[2][7] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0083_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold175 (.A(\s0.data_out[21][7] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0191_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold177 (.A(\s0.data_out[5][1] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0041_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold179 (.A(\s0.data_out[25][7] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold180 (.A(\s0.data_out[6][2] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold181 (.A(_2743_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold182 (.A(\s0.data_out[21][1] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold183 (.A(_1036_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold184 (.A(\s0.data_out[8][7] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold185 (.A(\s0.data_out[24][6] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0155_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold187 (.A(\s0.data_out[25][0] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0137_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold189 (.A(\s0.data_out[4][6] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0058_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold191 (.A(\s0.data_out[20][1] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0198_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold193 (.A(\s0.data_out[8][2] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0006_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold195 (.A(\s0.data_out[16][2] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0247_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold197 (.A(\s0.data_out[1][4] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold198 (.A(_3193_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold199 (.A(\s0.data_out[11][7] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0312_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold201 (.A(\s0.data_out[23][6] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold202 (.A(\s0.data_out[11][2] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold203 (.A(\s0.data_out[5][3] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0043_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold205 (.A(\s0.data_out[18][5] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0226_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold207 (.A(\s0.data_out[7][3] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0019_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold209 (.A(\s0.data_out[15][7] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0264_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold211 (.A(\s0.data_out[12][3] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0296_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold213 (.A(\s0.data_out[17][7] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold214 (.A(\s0.data_out[13][5] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0286_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold216 (.A(\s0.data_out[15][2] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold217 (.A(_1718_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold218 (.A(\s0.data_out[13][1] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold219 (.A(_1942_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold220 (.A(\s0.data_out[15][5] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold221 (.A(\s0.data_out[7][2] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0018_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold223 (.A(\s0.data_out[24][4] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0153_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold225 (.A(\s0.data_out[8][1] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0005_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold227 (.A(\s0.data_out[5][6] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0046_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold229 (.A(\s0.data_out[18][4] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0225_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold231 (.A(\s0.data_out[27][1] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0114_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold233 (.A(\s0.data_out[1][3] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold234 (.A(_3299_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold235 (.A(\s0.data_out[0][0] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold236 (.A(\s0.data_out[11][5] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0310_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold238 (.A(\s0.data_out[9][0] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold239 (.A(\s0.data_out[13][7] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0288_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold241 (.A(\s0.data_out[8][3] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold242 (.A(\s0.data_out[22][3] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold243 (.A(\s0.data_out[27][7] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0120_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold245 (.A(\s0.data_out[23][5] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0702_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold247 (.A(\s0.was_valid_out[16] [0]),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0241_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold249 (.A(\s0.was_valid_out[20] [0]),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0193_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold251 (.A(\s0.was_valid_out[1] [0]),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold252 (.A(\s0.data_out[15][0] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold253 (.A(\s0.data_out[2][5] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold254 (.A(_3198_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold255 (.A(\s0.data_out[4][7] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0059_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold257 (.A(\s0.data_out[10][6] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold258 (.A(\s0.data_out[18][2] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold259 (.A(_1372_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold260 (.A(\s0.data_out[7][0] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold261 (.A(_2621_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold262 (.A(\s0.data_out[24][2] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0151_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold264 (.A(\s0.data_out[9][5] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold265 (.A(\s0.data_out[3][7] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0071_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold267 (.A(\s0.data_out[14][0] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold268 (.A(_1824_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold269 (.A(\s0.data_out[17][6] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1504_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold271 (.A(\s0.data_out[8][6] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0010_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold273 (.A(\s0.data_out[4][4] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold274 (.A(_2972_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold275 (.A(\s0.data_out[20][3] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0200_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold277 (.A(\s0.data_out[5][2] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0042_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold279 (.A(\s0.data_out[14][2] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0271_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold281 (.A(\s0.data_out[11][0] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold282 (.A(\s0.data_out[5][5] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0045_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold284 (.A(\s0.data_out[16][0] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold285 (.A(\s0.data_out[6][4] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold286 (.A(_2750_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold287 (.A(\s0.data_out[19][3] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0212_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold289 (.A(\s0.data_out[22][1] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold290 (.A(\s0.data_out[10][1] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold291 (.A(\s0.data_out[12][5] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0298_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold293 (.A(\s0.data_out[19][2] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0211_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold295 (.A(\s0.data_out[9][3] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold296 (.A(_2291_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold297 (.A(_2292_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0327_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold299 (.A(\s0.data_out[6][7] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold300 (.A(_2644_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold301 (.A(\s0.data_out[26][1] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0126_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold303 (.A(\s0.data_out[9][4] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold304 (.A(\s0.was_valid_out[14] [0]),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0265_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold306 (.A(\s0.data_out[4][5] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold307 (.A(_2976_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold308 (.A(\s0.data_out[24][0] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold309 (.A(\s0.data_out[23][2] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0806_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold311 (.A(\s0.data_out[26][6] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold312 (.A(\s0.data_out[17][4] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold313 (.A(_1496_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold314 (.A(\s0.data_out[19][0] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold315 (.A(_1254_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold316 (.A(\s0.data_out[13][0] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold317 (.A(_1938_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold318 (.A(\s0.data_out[13][2] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold319 (.A(_1946_),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold320 (.A(\s0.was_valid_out[8] [0]),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold321 (.A(\s0.data_out[22][2] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold322 (.A(\s0.data_out[20][2] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold323 (.A(\s0.data_out[13][3] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0284_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold325 (.A(\s0.data_out[20][7] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0204_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold327 (.A(\s0.data_out[6][0] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold328 (.A(\s0.was_valid_out[24] [0]),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold329 (.A(\s0.data_out[2][1] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold330 (.A(_3184_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold331 (.A(\s0.data_out[3][4] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0068_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold333 (.A(\s0.data_out[21][4] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold334 (.A(\s0.data_out[3][2] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold335 (.A(_3079_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold336 (.A(\s0.data_out[10][0] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold337 (.A(\s0.data_out[2][0] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold338 (.A(_3180_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold339 (.A(\s0.data_out[17][5] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold340 (.A(\s0.data_out[12][6] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold341 (.A(\s0.data_out[4][0] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold342 (.A(_2957_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold343 (.A(\s0.data_out[14][7] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold344 (.A(\s0.data_out[21][0] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold345 (.A(_1032_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold346 (.A(\s0.data_out[21][6] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold347 (.A(\s0.data_out[16][4] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0249_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold349 (.A(\s0.data_out[11][6] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold350 (.A(_2183_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold351 (.A(\s0.data_out[22][5] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold352 (.A(\s0.data_out[14][6] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold353 (.A(_1844_),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold354 (.A(\s0.data_out[4][1] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold355 (.A(_2961_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold356 (.A(\s0.data_out[19][1] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0210_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold358 (.A(\s0.data_out[23][7] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold359 (.A(\s0.data_out[12][0] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold360 (.A(\s0.data_out[14][1] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold361 (.A(\s0.data_out[14][3] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold362 (.A(\s0.data_out[25][2] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0584_),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold364 (.A(\s0.data_out[20][0] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold365 (.A(\s0.shift_out[21] [0]),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold366 (.A(\s0.data_out[9][6] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold367 (.A(\s0.data_out[1][1] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold368 (.A(\s0.data_out[6][1] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold369 (.A(\s0.data_out[23][0] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0799_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold371 (.A(\s0.data_out[7][4] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold372 (.A(_2634_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold373 (.A(\s0.data_out[8][0] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold374 (.A(\s0.data_out[23][4] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold375 (.A(\s0.data_out[26][0] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold376 (.A(\s0.data_out[1][5] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold377 (.A(\s0.data_out[11][3] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0308_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold379 (.A(\s0.data_out[4][2] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold380 (.A(\s0.data_out[12][2] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0295_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold382 (.A(\s0.data_out[5][4] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold383 (.A(\s0.data_out[16][6] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold384 (.A(\s0.data_out[11][1] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold385 (.A(\s0.data_out[22][0] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold386 (.A(\s0.data_out[19][7] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0216_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold388 (.A(\s0.data_out[5][0] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold389 (.A(\s0.data_out[7][5] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold390 (.A(_2638_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold391 (.A(\s0.data_out[13][6] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold392 (.A(_1959_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold393 (.A(\s0.data_out[1][2] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold394 (.A(_3295_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold395 (.A(\s0.data_out[19][6] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0215_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold397 (.A(\s0.data_out[25][5] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold398 (.A(\s0.data_out[25][1] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0138_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold400 (.A(\s0.was_valid_out[27] [0]),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0109_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold402 (.A(\s0.data_out[3][1] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold403 (.A(_3075_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold404 (.A(\s0.data_out[8][4] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold405 (.A(\s0.data_out[2][2] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold406 (.A(\s0.data_out[25][3] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0140_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold408 (.A(\s0.data_out[25][6] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0599_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold410 (.A(\s0.data_out[6][6] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold411 (.A(\s0.data_out[17][0] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold412 (.A(\s0.data_out[20][6] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold413 (.A(\s0.data_out[3][0] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold414 (.A(\s0.data_out[14][5] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold415 (.A(\s0.data_out[2][3] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0079_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold417 (.A(\s0.data_out[15][3] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold418 (.A(\s0.data_out[18][0] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold419 (.A(\s0.data_out[11][4] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0309_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold421 (.A(\s0.data_out[19][4] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold422 (.A(\s0.data_out[1][0] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold423 (.A(_3288_),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold424 (.A(\s0.data_out[2][6] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold425 (.A(_3202_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold426 (.A(\s0.data_out[15][6] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold427 (.A(\s0.data_out[7][1] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0017_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold429 (.A(\s0.data_out[18][1] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold430 (.A(_1368_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold431 (.A(\s0.data_out[6][5] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold432 (.A(\s0.data_out[1][7] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold433 (.A(\s0.data_out[23][3] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0164_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold435 (.A(\s0.data_out[19][5] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold436 (.A(\s0.data_out[18][7] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold437 (.A(\s0.shift_out[3] [0]),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold438 (.A(\s0.data_out[15][4] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold439 (.A(\s0.data_out[18][6] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold440 (.A(_1385_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold441 (.A(\s0.data_out[7][6] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold442 (.A(_2642_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold443 (.A(\s0.data_out[3][5] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold444 (.A(\s0.data_out[8][5] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold445 (.A(\s0.data_out[15][1] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0258_),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold447 (.A(\s0.data_out[3][6] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold448 (.A(\s0.data_out[23][1] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0162_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold450 (.A(\s0.data_out[17][3] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold451 (.A(\s0.data_out[12][1] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0294_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold453 (.A(\s0.data_out[1][6] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold454 (.A(\s0.data_out[17][1] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold455 (.A(\s0.data_out[26][3] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0128_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold457 (.A(\s0.was_valid_out[18] [0]),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0217_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold459 (.A(\s0.valid_out[3] [0]),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold460 (.A(\s0.shift_out[5] [0]),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold461 (.A(\s0.data_new_delayed[2] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold462 (.A(\s0.shift_out[2] [0]),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold463 (.A(\s0.data_new_delayed[4] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold464 (.A(\s0.valid_out[13] [0]),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold465 (.A(\s0.data_new_delayed[0] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold466 (.A(\s0.data_out[20][6] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold467 (.A(_1053_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold468 (.A(\s0.data_out[9][6] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold469 (.A(\s0.valid_out[3] [0]),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold470 (.A(\s0.data_out[5][0] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold471 (.A(\s0.data_out[10][0] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold472 (.A(\s0.data_out[15][6] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold473 (.A(\s0.data_out[15][6] ),
    .X(net842));
 sg13g2_fill_1 FILLER_0_4 ();
 sg13g2_fill_2 FILLER_0_41 ();
 sg13g2_fill_1 FILLER_0_43 ();
 sg13g2_fill_1 FILLER_0_87 ();
 sg13g2_fill_1 FILLER_0_92 ();
 sg13g2_fill_1 FILLER_0_134 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_decap_4 FILLER_0_171 ();
 sg13g2_fill_1 FILLER_0_213 ();
 sg13g2_decap_4 FILLER_0_223 ();
 sg13g2_fill_2 FILLER_0_227 ();
 sg13g2_fill_2 FILLER_0_233 ();
 sg13g2_fill_1 FILLER_0_240 ();
 sg13g2_fill_2 FILLER_0_248 ();
 sg13g2_fill_2 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_4 FILLER_0_384 ();
 sg13g2_fill_2 FILLER_0_388 ();
 sg13g2_decap_4 FILLER_0_394 ();
 sg13g2_fill_1 FILLER_0_398 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_fill_1 FILLER_0_409 ();
 sg13g2_fill_2 FILLER_0_418 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_4 FILLER_0_441 ();
 sg13g2_fill_2 FILLER_0_445 ();
 sg13g2_fill_2 FILLER_0_479 ();
 sg13g2_decap_8 FILLER_0_526 ();
 sg13g2_fill_1 FILLER_0_533 ();
 sg13g2_fill_1 FILLER_0_538 ();
 sg13g2_decap_8 FILLER_0_543 ();
 sg13g2_fill_2 FILLER_0_550 ();
 sg13g2_fill_1 FILLER_0_552 ();
 sg13g2_fill_1 FILLER_0_566 ();
 sg13g2_fill_1 FILLER_0_604 ();
 sg13g2_decap_8 FILLER_0_617 ();
 sg13g2_decap_8 FILLER_0_624 ();
 sg13g2_decap_8 FILLER_0_631 ();
 sg13g2_decap_8 FILLER_0_638 ();
 sg13g2_decap_8 FILLER_0_645 ();
 sg13g2_decap_8 FILLER_0_652 ();
 sg13g2_decap_8 FILLER_0_659 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_8 FILLER_0_673 ();
 sg13g2_decap_8 FILLER_0_680 ();
 sg13g2_decap_4 FILLER_0_687 ();
 sg13g2_fill_1 FILLER_0_691 ();
 sg13g2_decap_8 FILLER_0_696 ();
 sg13g2_decap_8 FILLER_0_703 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_773 ();
 sg13g2_decap_8 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_787 ();
 sg13g2_decap_8 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_843 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_0_878 ();
 sg13g2_decap_8 FILLER_0_885 ();
 sg13g2_decap_8 FILLER_0_892 ();
 sg13g2_decap_8 FILLER_0_899 ();
 sg13g2_decap_8 FILLER_0_906 ();
 sg13g2_decap_8 FILLER_0_913 ();
 sg13g2_decap_8 FILLER_0_920 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_4 FILLER_0_1025 ();
 sg13g2_fill_2 FILLER_1_54 ();
 sg13g2_fill_2 FILLER_1_83 ();
 sg13g2_fill_1 FILLER_1_132 ();
 sg13g2_fill_1 FILLER_1_167 ();
 sg13g2_fill_1 FILLER_1_223 ();
 sg13g2_fill_1 FILLER_1_251 ();
 sg13g2_fill_1 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_446 ();
 sg13g2_decap_4 FILLER_1_453 ();
 sg13g2_fill_1 FILLER_1_457 ();
 sg13g2_fill_1 FILLER_1_528 ();
 sg13g2_decap_4 FILLER_1_616 ();
 sg13g2_fill_2 FILLER_1_620 ();
 sg13g2_decap_8 FILLER_1_649 ();
 sg13g2_fill_1 FILLER_1_656 ();
 sg13g2_decap_8 FILLER_1_666 ();
 sg13g2_fill_2 FILLER_1_673 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_fill_1 FILLER_1_686 ();
 sg13g2_decap_4 FILLER_1_715 ();
 sg13g2_fill_2 FILLER_1_719 ();
 sg13g2_decap_8 FILLER_1_725 ();
 sg13g2_decap_8 FILLER_1_732 ();
 sg13g2_decap_8 FILLER_1_739 ();
 sg13g2_decap_8 FILLER_1_746 ();
 sg13g2_decap_8 FILLER_1_753 ();
 sg13g2_decap_8 FILLER_1_760 ();
 sg13g2_decap_8 FILLER_1_767 ();
 sg13g2_decap_8 FILLER_1_774 ();
 sg13g2_decap_8 FILLER_1_781 ();
 sg13g2_decap_8 FILLER_1_788 ();
 sg13g2_decap_8 FILLER_1_795 ();
 sg13g2_decap_8 FILLER_1_802 ();
 sg13g2_decap_8 FILLER_1_809 ();
 sg13g2_decap_8 FILLER_1_816 ();
 sg13g2_decap_8 FILLER_1_823 ();
 sg13g2_decap_8 FILLER_1_830 ();
 sg13g2_decap_8 FILLER_1_837 ();
 sg13g2_decap_8 FILLER_1_844 ();
 sg13g2_decap_8 FILLER_1_851 ();
 sg13g2_decap_8 FILLER_1_858 ();
 sg13g2_decap_8 FILLER_1_865 ();
 sg13g2_decap_8 FILLER_1_872 ();
 sg13g2_decap_8 FILLER_1_879 ();
 sg13g2_decap_8 FILLER_1_886 ();
 sg13g2_decap_8 FILLER_1_893 ();
 sg13g2_decap_8 FILLER_1_900 ();
 sg13g2_decap_8 FILLER_1_907 ();
 sg13g2_decap_8 FILLER_1_914 ();
 sg13g2_decap_8 FILLER_1_921 ();
 sg13g2_decap_8 FILLER_1_928 ();
 sg13g2_decap_8 FILLER_1_935 ();
 sg13g2_decap_8 FILLER_1_942 ();
 sg13g2_decap_8 FILLER_1_949 ();
 sg13g2_decap_8 FILLER_1_956 ();
 sg13g2_decap_8 FILLER_1_963 ();
 sg13g2_decap_8 FILLER_1_970 ();
 sg13g2_decap_8 FILLER_1_977 ();
 sg13g2_decap_8 FILLER_1_984 ();
 sg13g2_decap_8 FILLER_1_991 ();
 sg13g2_decap_8 FILLER_1_998 ();
 sg13g2_decap_8 FILLER_1_1005 ();
 sg13g2_decap_8 FILLER_1_1012 ();
 sg13g2_decap_8 FILLER_1_1019 ();
 sg13g2_fill_2 FILLER_1_1026 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_fill_2 FILLER_2_4 ();
 sg13g2_fill_1 FILLER_2_6 ();
 sg13g2_fill_1 FILLER_2_60 ();
 sg13g2_fill_2 FILLER_2_74 ();
 sg13g2_fill_1 FILLER_2_76 ();
 sg13g2_fill_1 FILLER_2_126 ();
 sg13g2_fill_2 FILLER_2_192 ();
 sg13g2_fill_2 FILLER_2_258 ();
 sg13g2_fill_1 FILLER_2_260 ();
 sg13g2_fill_1 FILLER_2_265 ();
 sg13g2_fill_2 FILLER_2_275 ();
 sg13g2_fill_1 FILLER_2_277 ();
 sg13g2_decap_4 FILLER_2_282 ();
 sg13g2_fill_2 FILLER_2_286 ();
 sg13g2_fill_2 FILLER_2_298 ();
 sg13g2_fill_2 FILLER_2_347 ();
 sg13g2_fill_2 FILLER_2_359 ();
 sg13g2_fill_2 FILLER_2_377 ();
 sg13g2_fill_1 FILLER_2_379 ();
 sg13g2_fill_1 FILLER_2_423 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_4 FILLER_2_452 ();
 sg13g2_fill_1 FILLER_2_522 ();
 sg13g2_fill_2 FILLER_2_542 ();
 sg13g2_fill_2 FILLER_2_553 ();
 sg13g2_fill_1 FILLER_2_555 ();
 sg13g2_fill_2 FILLER_2_576 ();
 sg13g2_fill_1 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_4 FILLER_2_623 ();
 sg13g2_fill_1 FILLER_2_631 ();
 sg13g2_fill_1 FILLER_2_637 ();
 sg13g2_fill_2 FILLER_2_651 ();
 sg13g2_fill_2 FILLER_2_674 ();
 sg13g2_decap_4 FILLER_2_709 ();
 sg13g2_fill_2 FILLER_2_713 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_fill_1 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_761 ();
 sg13g2_decap_8 FILLER_2_768 ();
 sg13g2_decap_8 FILLER_2_775 ();
 sg13g2_decap_8 FILLER_2_782 ();
 sg13g2_decap_8 FILLER_2_789 ();
 sg13g2_decap_8 FILLER_2_796 ();
 sg13g2_decap_8 FILLER_2_803 ();
 sg13g2_decap_8 FILLER_2_810 ();
 sg13g2_decap_8 FILLER_2_817 ();
 sg13g2_decap_8 FILLER_2_824 ();
 sg13g2_decap_8 FILLER_2_831 ();
 sg13g2_decap_8 FILLER_2_838 ();
 sg13g2_decap_8 FILLER_2_845 ();
 sg13g2_decap_8 FILLER_2_852 ();
 sg13g2_decap_8 FILLER_2_859 ();
 sg13g2_decap_8 FILLER_2_866 ();
 sg13g2_decap_8 FILLER_2_873 ();
 sg13g2_decap_8 FILLER_2_880 ();
 sg13g2_decap_8 FILLER_2_887 ();
 sg13g2_decap_8 FILLER_2_894 ();
 sg13g2_decap_8 FILLER_2_901 ();
 sg13g2_decap_8 FILLER_2_908 ();
 sg13g2_decap_8 FILLER_2_915 ();
 sg13g2_decap_8 FILLER_2_922 ();
 sg13g2_decap_8 FILLER_2_929 ();
 sg13g2_decap_8 FILLER_2_936 ();
 sg13g2_decap_8 FILLER_2_943 ();
 sg13g2_decap_8 FILLER_2_950 ();
 sg13g2_decap_8 FILLER_2_957 ();
 sg13g2_decap_8 FILLER_2_964 ();
 sg13g2_decap_8 FILLER_2_971 ();
 sg13g2_decap_8 FILLER_2_978 ();
 sg13g2_decap_8 FILLER_2_985 ();
 sg13g2_decap_8 FILLER_2_992 ();
 sg13g2_decap_8 FILLER_2_999 ();
 sg13g2_decap_8 FILLER_2_1006 ();
 sg13g2_decap_8 FILLER_2_1013 ();
 sg13g2_decap_8 FILLER_2_1020 ();
 sg13g2_fill_2 FILLER_2_1027 ();
 sg13g2_fill_2 FILLER_3_37 ();
 sg13g2_fill_2 FILLER_3_73 ();
 sg13g2_fill_2 FILLER_3_88 ();
 sg13g2_fill_2 FILLER_3_94 ();
 sg13g2_fill_1 FILLER_3_96 ();
 sg13g2_fill_2 FILLER_3_110 ();
 sg13g2_fill_2 FILLER_3_157 ();
 sg13g2_fill_1 FILLER_3_200 ();
 sg13g2_fill_1 FILLER_3_233 ();
 sg13g2_fill_2 FILLER_3_244 ();
 sg13g2_fill_1 FILLER_3_246 ();
 sg13g2_fill_2 FILLER_3_252 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_1 FILLER_3_328 ();
 sg13g2_fill_2 FILLER_3_336 ();
 sg13g2_fill_1 FILLER_3_338 ();
 sg13g2_fill_2 FILLER_3_360 ();
 sg13g2_fill_2 FILLER_3_379 ();
 sg13g2_fill_2 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_438 ();
 sg13g2_fill_1 FILLER_3_471 ();
 sg13g2_fill_1 FILLER_3_482 ();
 sg13g2_fill_1 FILLER_3_504 ();
 sg13g2_fill_2 FILLER_3_514 ();
 sg13g2_fill_1 FILLER_3_516 ();
 sg13g2_fill_2 FILLER_3_522 ();
 sg13g2_fill_1 FILLER_3_524 ();
 sg13g2_fill_2 FILLER_3_558 ();
 sg13g2_fill_1 FILLER_3_560 ();
 sg13g2_fill_1 FILLER_3_567 ();
 sg13g2_fill_2 FILLER_3_621 ();
 sg13g2_decap_8 FILLER_3_627 ();
 sg13g2_fill_1 FILLER_3_634 ();
 sg13g2_fill_2 FILLER_3_676 ();
 sg13g2_fill_1 FILLER_3_678 ();
 sg13g2_fill_2 FILLER_3_702 ();
 sg13g2_fill_2 FILLER_3_718 ();
 sg13g2_fill_2 FILLER_3_725 ();
 sg13g2_fill_2 FILLER_3_732 ();
 sg13g2_fill_1 FILLER_3_734 ();
 sg13g2_fill_2 FILLER_3_748 ();
 sg13g2_fill_1 FILLER_3_750 ();
 sg13g2_decap_8 FILLER_3_779 ();
 sg13g2_decap_8 FILLER_3_786 ();
 sg13g2_decap_8 FILLER_3_793 ();
 sg13g2_decap_8 FILLER_3_800 ();
 sg13g2_decap_8 FILLER_3_807 ();
 sg13g2_decap_8 FILLER_3_814 ();
 sg13g2_decap_8 FILLER_3_821 ();
 sg13g2_decap_8 FILLER_3_828 ();
 sg13g2_fill_2 FILLER_3_835 ();
 sg13g2_fill_2 FILLER_3_841 ();
 sg13g2_fill_1 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_848 ();
 sg13g2_decap_8 FILLER_3_855 ();
 sg13g2_decap_4 FILLER_3_862 ();
 sg13g2_decap_8 FILLER_3_870 ();
 sg13g2_decap_8 FILLER_3_877 ();
 sg13g2_decap_8 FILLER_3_884 ();
 sg13g2_decap_8 FILLER_3_891 ();
 sg13g2_decap_8 FILLER_3_898 ();
 sg13g2_decap_8 FILLER_3_905 ();
 sg13g2_decap_8 FILLER_3_912 ();
 sg13g2_decap_8 FILLER_3_919 ();
 sg13g2_decap_8 FILLER_3_926 ();
 sg13g2_decap_8 FILLER_3_933 ();
 sg13g2_decap_8 FILLER_3_940 ();
 sg13g2_decap_8 FILLER_3_947 ();
 sg13g2_decap_8 FILLER_3_954 ();
 sg13g2_decap_8 FILLER_3_961 ();
 sg13g2_decap_8 FILLER_3_968 ();
 sg13g2_decap_8 FILLER_3_975 ();
 sg13g2_decap_8 FILLER_3_982 ();
 sg13g2_decap_8 FILLER_3_989 ();
 sg13g2_decap_8 FILLER_3_996 ();
 sg13g2_decap_8 FILLER_3_1003 ();
 sg13g2_decap_8 FILLER_3_1010 ();
 sg13g2_decap_8 FILLER_3_1017 ();
 sg13g2_decap_4 FILLER_3_1024 ();
 sg13g2_fill_1 FILLER_3_1028 ();
 sg13g2_fill_2 FILLER_4_36 ();
 sg13g2_fill_1 FILLER_4_130 ();
 sg13g2_fill_2 FILLER_4_149 ();
 sg13g2_fill_2 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_228 ();
 sg13g2_fill_1 FILLER_4_272 ();
 sg13g2_fill_2 FILLER_4_295 ();
 sg13g2_fill_1 FILLER_4_297 ();
 sg13g2_fill_1 FILLER_4_325 ();
 sg13g2_fill_1 FILLER_4_331 ();
 sg13g2_fill_1 FILLER_4_337 ();
 sg13g2_fill_1 FILLER_4_351 ();
 sg13g2_fill_2 FILLER_4_371 ();
 sg13g2_fill_1 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_482 ();
 sg13g2_fill_2 FILLER_4_545 ();
 sg13g2_fill_2 FILLER_4_552 ();
 sg13g2_fill_1 FILLER_4_580 ();
 sg13g2_fill_2 FILLER_4_586 ();
 sg13g2_fill_2 FILLER_4_615 ();
 sg13g2_fill_1 FILLER_4_617 ();
 sg13g2_decap_8 FILLER_4_787 ();
 sg13g2_decap_8 FILLER_4_794 ();
 sg13g2_fill_2 FILLER_4_801 ();
 sg13g2_decap_8 FILLER_4_822 ();
 sg13g2_fill_2 FILLER_4_871 ();
 sg13g2_fill_1 FILLER_4_873 ();
 sg13g2_decap_8 FILLER_4_906 ();
 sg13g2_fill_2 FILLER_4_913 ();
 sg13g2_decap_8 FILLER_4_919 ();
 sg13g2_decap_8 FILLER_4_926 ();
 sg13g2_decap_8 FILLER_4_933 ();
 sg13g2_decap_8 FILLER_4_940 ();
 sg13g2_decap_8 FILLER_4_947 ();
 sg13g2_decap_8 FILLER_4_954 ();
 sg13g2_decap_8 FILLER_4_961 ();
 sg13g2_decap_8 FILLER_4_968 ();
 sg13g2_decap_8 FILLER_4_975 ();
 sg13g2_decap_8 FILLER_4_982 ();
 sg13g2_decap_8 FILLER_4_989 ();
 sg13g2_decap_8 FILLER_4_996 ();
 sg13g2_decap_8 FILLER_4_1003 ();
 sg13g2_decap_8 FILLER_4_1010 ();
 sg13g2_decap_8 FILLER_4_1017 ();
 sg13g2_decap_4 FILLER_4_1024 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_fill_1 FILLER_5_4 ();
 sg13g2_fill_2 FILLER_5_32 ();
 sg13g2_fill_1 FILLER_5_54 ();
 sg13g2_fill_1 FILLER_5_60 ();
 sg13g2_fill_1 FILLER_5_66 ();
 sg13g2_fill_2 FILLER_5_72 ();
 sg13g2_fill_1 FILLER_5_93 ();
 sg13g2_fill_1 FILLER_5_101 ();
 sg13g2_fill_1 FILLER_5_121 ();
 sg13g2_fill_2 FILLER_5_135 ();
 sg13g2_fill_1 FILLER_5_226 ();
 sg13g2_fill_1 FILLER_5_259 ();
 sg13g2_fill_2 FILLER_5_265 ();
 sg13g2_fill_2 FILLER_5_337 ();
 sg13g2_fill_1 FILLER_5_339 ();
 sg13g2_fill_2 FILLER_5_345 ();
 sg13g2_fill_1 FILLER_5_347 ();
 sg13g2_decap_4 FILLER_5_384 ();
 sg13g2_fill_1 FILLER_5_398 ();
 sg13g2_fill_1 FILLER_5_447 ();
 sg13g2_fill_2 FILLER_5_507 ();
 sg13g2_fill_2 FILLER_5_514 ();
 sg13g2_fill_1 FILLER_5_516 ();
 sg13g2_fill_2 FILLER_5_527 ();
 sg13g2_fill_2 FILLER_5_547 ();
 sg13g2_fill_1 FILLER_5_562 ();
 sg13g2_fill_1 FILLER_5_568 ();
 sg13g2_fill_2 FILLER_5_586 ();
 sg13g2_fill_2 FILLER_5_598 ();
 sg13g2_fill_2 FILLER_5_657 ();
 sg13g2_decap_4 FILLER_5_720 ();
 sg13g2_fill_1 FILLER_5_724 ();
 sg13g2_fill_1 FILLER_5_734 ();
 sg13g2_fill_2 FILLER_5_775 ();
 sg13g2_fill_2 FILLER_5_914 ();
 sg13g2_decap_8 FILLER_5_926 ();
 sg13g2_decap_4 FILLER_5_933 ();
 sg13g2_fill_1 FILLER_5_937 ();
 sg13g2_decap_8 FILLER_5_942 ();
 sg13g2_decap_8 FILLER_5_949 ();
 sg13g2_decap_8 FILLER_5_956 ();
 sg13g2_decap_8 FILLER_5_963 ();
 sg13g2_decap_8 FILLER_5_970 ();
 sg13g2_decap_8 FILLER_5_977 ();
 sg13g2_decap_8 FILLER_5_984 ();
 sg13g2_decap_8 FILLER_5_991 ();
 sg13g2_decap_8 FILLER_5_998 ();
 sg13g2_decap_8 FILLER_5_1005 ();
 sg13g2_decap_8 FILLER_5_1012 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_fill_2 FILLER_5_1026 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_fill_1 FILLER_6_41 ();
 sg13g2_fill_2 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_64 ();
 sg13g2_fill_2 FILLER_6_108 ();
 sg13g2_fill_2 FILLER_6_115 ();
 sg13g2_fill_1 FILLER_6_117 ();
 sg13g2_fill_2 FILLER_6_136 ();
 sg13g2_fill_1 FILLER_6_138 ();
 sg13g2_fill_2 FILLER_6_143 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_fill_2 FILLER_6_168 ();
 sg13g2_fill_2 FILLER_6_186 ();
 sg13g2_decap_4 FILLER_6_196 ();
 sg13g2_fill_2 FILLER_6_200 ();
 sg13g2_fill_2 FILLER_6_217 ();
 sg13g2_fill_2 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_266 ();
 sg13g2_fill_1 FILLER_6_268 ();
 sg13g2_fill_1 FILLER_6_276 ();
 sg13g2_fill_2 FILLER_6_312 ();
 sg13g2_fill_1 FILLER_6_314 ();
 sg13g2_fill_1 FILLER_6_323 ();
 sg13g2_fill_2 FILLER_6_340 ();
 sg13g2_fill_2 FILLER_6_346 ();
 sg13g2_fill_1 FILLER_6_348 ();
 sg13g2_fill_2 FILLER_6_362 ();
 sg13g2_fill_2 FILLER_6_388 ();
 sg13g2_fill_2 FILLER_6_403 ();
 sg13g2_decap_4 FILLER_6_433 ();
 sg13g2_fill_2 FILLER_6_437 ();
 sg13g2_fill_2 FILLER_6_470 ();
 sg13g2_fill_1 FILLER_6_487 ();
 sg13g2_fill_1 FILLER_6_530 ();
 sg13g2_fill_1 FILLER_6_594 ();
 sg13g2_fill_2 FILLER_6_628 ();
 sg13g2_fill_2 FILLER_6_645 ();
 sg13g2_fill_1 FILLER_6_652 ();
 sg13g2_fill_1 FILLER_6_684 ();
 sg13g2_fill_1 FILLER_6_713 ();
 sg13g2_fill_2 FILLER_6_794 ();
 sg13g2_fill_2 FILLER_6_836 ();
 sg13g2_fill_1 FILLER_6_838 ();
 sg13g2_fill_2 FILLER_6_863 ();
 sg13g2_fill_1 FILLER_6_900 ();
 sg13g2_fill_1 FILLER_6_929 ();
 sg13g2_fill_1 FILLER_6_935 ();
 sg13g2_fill_1 FILLER_6_945 ();
 sg13g2_decap_8 FILLER_6_955 ();
 sg13g2_decap_8 FILLER_6_962 ();
 sg13g2_decap_8 FILLER_6_969 ();
 sg13g2_decap_8 FILLER_6_976 ();
 sg13g2_decap_8 FILLER_6_983 ();
 sg13g2_decap_8 FILLER_6_990 ();
 sg13g2_decap_8 FILLER_6_997 ();
 sg13g2_decap_8 FILLER_6_1004 ();
 sg13g2_decap_8 FILLER_6_1011 ();
 sg13g2_decap_8 FILLER_6_1018 ();
 sg13g2_decap_4 FILLER_6_1025 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_67 ();
 sg13g2_fill_1 FILLER_7_78 ();
 sg13g2_fill_1 FILLER_7_84 ();
 sg13g2_fill_2 FILLER_7_100 ();
 sg13g2_decap_4 FILLER_7_109 ();
 sg13g2_fill_1 FILLER_7_113 ();
 sg13g2_decap_4 FILLER_7_118 ();
 sg13g2_fill_1 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_178 ();
 sg13g2_decap_8 FILLER_7_183 ();
 sg13g2_decap_8 FILLER_7_190 ();
 sg13g2_decap_4 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_201 ();
 sg13g2_fill_1 FILLER_7_281 ();
 sg13g2_fill_2 FILLER_7_312 ();
 sg13g2_fill_1 FILLER_7_314 ();
 sg13g2_fill_2 FILLER_7_338 ();
 sg13g2_fill_1 FILLER_7_340 ();
 sg13g2_fill_1 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_415 ();
 sg13g2_fill_2 FILLER_7_426 ();
 sg13g2_decap_4 FILLER_7_441 ();
 sg13g2_fill_1 FILLER_7_478 ();
 sg13g2_decap_4 FILLER_7_505 ();
 sg13g2_fill_1 FILLER_7_514 ();
 sg13g2_decap_8 FILLER_7_520 ();
 sg13g2_fill_2 FILLER_7_527 ();
 sg13g2_fill_2 FILLER_7_554 ();
 sg13g2_fill_2 FILLER_7_591 ();
 sg13g2_fill_1 FILLER_7_593 ();
 sg13g2_fill_1 FILLER_7_604 ();
 sg13g2_fill_1 FILLER_7_613 ();
 sg13g2_fill_2 FILLER_7_623 ();
 sg13g2_fill_2 FILLER_7_668 ();
 sg13g2_fill_2 FILLER_7_679 ();
 sg13g2_fill_2 FILLER_7_697 ();
 sg13g2_fill_2 FILLER_7_723 ();
 sg13g2_fill_1 FILLER_7_758 ();
 sg13g2_fill_1 FILLER_7_766 ();
 sg13g2_fill_2 FILLER_7_841 ();
 sg13g2_fill_1 FILLER_7_884 ();
 sg13g2_fill_1 FILLER_7_916 ();
 sg13g2_fill_2 FILLER_7_922 ();
 sg13g2_fill_1 FILLER_7_924 ();
 sg13g2_fill_1 FILLER_7_932 ();
 sg13g2_decap_8 FILLER_7_961 ();
 sg13g2_decap_8 FILLER_7_968 ();
 sg13g2_decap_8 FILLER_7_975 ();
 sg13g2_decap_8 FILLER_7_982 ();
 sg13g2_decap_8 FILLER_7_989 ();
 sg13g2_decap_8 FILLER_7_996 ();
 sg13g2_decap_8 FILLER_7_1003 ();
 sg13g2_decap_8 FILLER_7_1010 ();
 sg13g2_decap_8 FILLER_7_1017 ();
 sg13g2_decap_4 FILLER_7_1024 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_41 ();
 sg13g2_fill_2 FILLER_8_83 ();
 sg13g2_fill_1 FILLER_8_148 ();
 sg13g2_decap_4 FILLER_8_201 ();
 sg13g2_fill_1 FILLER_8_205 ();
 sg13g2_decap_8 FILLER_8_226 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_fill_2 FILLER_8_245 ();
 sg13g2_fill_1 FILLER_8_247 ();
 sg13g2_decap_4 FILLER_8_262 ();
 sg13g2_fill_1 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_311 ();
 sg13g2_fill_1 FILLER_8_313 ();
 sg13g2_fill_1 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_1 FILLER_8_375 ();
 sg13g2_fill_2 FILLER_8_419 ();
 sg13g2_fill_1 FILLER_8_421 ();
 sg13g2_fill_2 FILLER_8_437 ();
 sg13g2_fill_1 FILLER_8_460 ();
 sg13g2_decap_4 FILLER_8_489 ();
 sg13g2_decap_8 FILLER_8_523 ();
 sg13g2_decap_8 FILLER_8_530 ();
 sg13g2_fill_2 FILLER_8_588 ();
 sg13g2_fill_2 FILLER_8_643 ();
 sg13g2_fill_1 FILLER_8_645 ();
 sg13g2_fill_1 FILLER_8_689 ();
 sg13g2_fill_1 FILLER_8_700 ();
 sg13g2_fill_2 FILLER_8_717 ();
 sg13g2_fill_1 FILLER_8_732 ();
 sg13g2_fill_2 FILLER_8_742 ();
 sg13g2_fill_1 FILLER_8_760 ();
 sg13g2_fill_1 FILLER_8_766 ();
 sg13g2_fill_1 FILLER_8_803 ();
 sg13g2_fill_1 FILLER_8_874 ();
 sg13g2_fill_1 FILLER_8_893 ();
 sg13g2_decap_8 FILLER_8_946 ();
 sg13g2_decap_8 FILLER_8_953 ();
 sg13g2_decap_8 FILLER_8_960 ();
 sg13g2_decap_8 FILLER_8_967 ();
 sg13g2_decap_8 FILLER_8_974 ();
 sg13g2_decap_8 FILLER_8_981 ();
 sg13g2_decap_8 FILLER_8_988 ();
 sg13g2_decap_8 FILLER_8_995 ();
 sg13g2_decap_8 FILLER_8_1002 ();
 sg13g2_decap_8 FILLER_8_1009 ();
 sg13g2_decap_8 FILLER_8_1016 ();
 sg13g2_decap_4 FILLER_8_1023 ();
 sg13g2_fill_2 FILLER_8_1027 ();
 sg13g2_fill_2 FILLER_9_65 ();
 sg13g2_fill_2 FILLER_9_85 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_142 ();
 sg13g2_fill_2 FILLER_9_171 ();
 sg13g2_fill_1 FILLER_9_221 ();
 sg13g2_fill_2 FILLER_9_226 ();
 sg13g2_fill_2 FILLER_9_238 ();
 sg13g2_fill_1 FILLER_9_240 ();
 sg13g2_fill_2 FILLER_9_250 ();
 sg13g2_fill_2 FILLER_9_269 ();
 sg13g2_fill_1 FILLER_9_271 ();
 sg13g2_decap_8 FILLER_9_276 ();
 sg13g2_decap_4 FILLER_9_283 ();
 sg13g2_fill_2 FILLER_9_344 ();
 sg13g2_fill_1 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_442 ();
 sg13g2_fill_1 FILLER_9_476 ();
 sg13g2_decap_4 FILLER_9_486 ();
 sg13g2_decap_4 FILLER_9_521 ();
 sg13g2_fill_2 FILLER_9_525 ();
 sg13g2_fill_1 FILLER_9_563 ();
 sg13g2_decap_8 FILLER_9_600 ();
 sg13g2_fill_2 FILLER_9_607 ();
 sg13g2_fill_2 FILLER_9_658 ();
 sg13g2_fill_1 FILLER_9_667 ();
 sg13g2_fill_2 FILLER_9_678 ();
 sg13g2_fill_1 FILLER_9_713 ();
 sg13g2_fill_2 FILLER_9_763 ();
 sg13g2_fill_1 FILLER_9_765 ();
 sg13g2_fill_2 FILLER_9_786 ();
 sg13g2_fill_1 FILLER_9_793 ();
 sg13g2_fill_2 FILLER_9_849 ();
 sg13g2_fill_1 FILLER_9_851 ();
 sg13g2_fill_2 FILLER_9_905 ();
 sg13g2_fill_2 FILLER_9_920 ();
 sg13g2_fill_1 FILLER_9_934 ();
 sg13g2_decap_8 FILLER_9_944 ();
 sg13g2_decap_8 FILLER_9_951 ();
 sg13g2_decap_8 FILLER_9_958 ();
 sg13g2_decap_8 FILLER_9_965 ();
 sg13g2_decap_8 FILLER_9_972 ();
 sg13g2_decap_8 FILLER_9_979 ();
 sg13g2_decap_8 FILLER_9_986 ();
 sg13g2_decap_8 FILLER_9_993 ();
 sg13g2_decap_8 FILLER_9_1000 ();
 sg13g2_decap_8 FILLER_9_1007 ();
 sg13g2_decap_8 FILLER_9_1014 ();
 sg13g2_decap_8 FILLER_9_1021 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_1 FILLER_10_6 ();
 sg13g2_fill_2 FILLER_10_28 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_136 ();
 sg13g2_fill_1 FILLER_10_138 ();
 sg13g2_fill_2 FILLER_10_157 ();
 sg13g2_fill_1 FILLER_10_228 ();
 sg13g2_decap_4 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_fill_2 FILLER_10_338 ();
 sg13g2_fill_1 FILLER_10_340 ();
 sg13g2_fill_2 FILLER_10_346 ();
 sg13g2_fill_2 FILLER_10_388 ();
 sg13g2_fill_1 FILLER_10_390 ();
 sg13g2_fill_2 FILLER_10_400 ();
 sg13g2_fill_1 FILLER_10_510 ();
 sg13g2_decap_8 FILLER_10_516 ();
 sg13g2_fill_2 FILLER_10_523 ();
 sg13g2_fill_2 FILLER_10_555 ();
 sg13g2_fill_1 FILLER_10_557 ();
 sg13g2_decap_4 FILLER_10_571 ();
 sg13g2_decap_4 FILLER_10_591 ();
 sg13g2_fill_1 FILLER_10_595 ();
 sg13g2_decap_4 FILLER_10_613 ();
 sg13g2_fill_2 FILLER_10_617 ();
 sg13g2_fill_1 FILLER_10_636 ();
 sg13g2_decap_4 FILLER_10_662 ();
 sg13g2_fill_2 FILLER_10_666 ();
 sg13g2_decap_8 FILLER_10_706 ();
 sg13g2_decap_4 FILLER_10_713 ();
 sg13g2_fill_2 FILLER_10_717 ();
 sg13g2_fill_2 FILLER_10_745 ();
 sg13g2_fill_1 FILLER_10_747 ();
 sg13g2_decap_4 FILLER_10_769 ();
 sg13g2_fill_2 FILLER_10_773 ();
 sg13g2_fill_2 FILLER_10_795 ();
 sg13g2_fill_1 FILLER_10_797 ();
 sg13g2_fill_1 FILLER_10_832 ();
 sg13g2_fill_2 FILLER_10_848 ();
 sg13g2_fill_1 FILLER_10_860 ();
 sg13g2_fill_1 FILLER_10_880 ();
 sg13g2_fill_2 FILLER_10_903 ();
 sg13g2_fill_2 FILLER_10_914 ();
 sg13g2_decap_8 FILLER_10_963 ();
 sg13g2_decap_8 FILLER_10_970 ();
 sg13g2_decap_8 FILLER_10_977 ();
 sg13g2_decap_8 FILLER_10_984 ();
 sg13g2_decap_8 FILLER_10_991 ();
 sg13g2_decap_8 FILLER_10_998 ();
 sg13g2_decap_8 FILLER_10_1005 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_fill_2 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_fill_1 FILLER_11_4 ();
 sg13g2_fill_1 FILLER_11_48 ();
 sg13g2_fill_1 FILLER_11_94 ();
 sg13g2_fill_2 FILLER_11_108 ();
 sg13g2_fill_1 FILLER_11_110 ();
 sg13g2_fill_2 FILLER_11_117 ();
 sg13g2_fill_2 FILLER_11_138 ();
 sg13g2_fill_2 FILLER_11_152 ();
 sg13g2_fill_1 FILLER_11_158 ();
 sg13g2_fill_2 FILLER_11_180 ();
 sg13g2_fill_1 FILLER_11_224 ();
 sg13g2_fill_2 FILLER_11_230 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_301 ();
 sg13g2_fill_2 FILLER_11_324 ();
 sg13g2_fill_1 FILLER_11_326 ();
 sg13g2_fill_2 FILLER_11_337 ();
 sg13g2_fill_2 FILLER_11_357 ();
 sg13g2_fill_1 FILLER_11_409 ();
 sg13g2_fill_2 FILLER_11_463 ();
 sg13g2_fill_2 FILLER_11_494 ();
 sg13g2_decap_4 FILLER_11_520 ();
 sg13g2_fill_2 FILLER_11_540 ();
 sg13g2_fill_1 FILLER_11_542 ();
 sg13g2_decap_8 FILLER_11_570 ();
 sg13g2_fill_1 FILLER_11_645 ();
 sg13g2_fill_1 FILLER_11_651 ();
 sg13g2_fill_2 FILLER_11_657 ();
 sg13g2_fill_2 FILLER_11_682 ();
 sg13g2_fill_1 FILLER_11_719 ();
 sg13g2_fill_2 FILLER_11_733 ();
 sg13g2_fill_1 FILLER_11_735 ();
 sg13g2_fill_1 FILLER_11_751 ();
 sg13g2_fill_1 FILLER_11_775 ();
 sg13g2_fill_1 FILLER_11_810 ();
 sg13g2_fill_2 FILLER_11_846 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_fill_1 FILLER_11_874 ();
 sg13g2_fill_2 FILLER_11_901 ();
 sg13g2_fill_1 FILLER_11_948 ();
 sg13g2_decap_8 FILLER_11_965 ();
 sg13g2_decap_8 FILLER_11_972 ();
 sg13g2_decap_8 FILLER_11_979 ();
 sg13g2_decap_8 FILLER_11_986 ();
 sg13g2_decap_8 FILLER_11_993 ();
 sg13g2_decap_8 FILLER_11_1000 ();
 sg13g2_decap_8 FILLER_11_1007 ();
 sg13g2_decap_8 FILLER_11_1014 ();
 sg13g2_decap_8 FILLER_11_1021 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_fill_1 FILLER_12_35 ();
 sg13g2_fill_2 FILLER_12_58 ();
 sg13g2_fill_1 FILLER_12_79 ();
 sg13g2_fill_1 FILLER_12_90 ();
 sg13g2_fill_1 FILLER_12_135 ();
 sg13g2_fill_1 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_158 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_261 ();
 sg13g2_fill_2 FILLER_12_292 ();
 sg13g2_decap_4 FILLER_12_320 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_fill_1 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_436 ();
 sg13g2_fill_2 FILLER_12_452 ();
 sg13g2_fill_2 FILLER_12_504 ();
 sg13g2_fill_2 FILLER_12_548 ();
 sg13g2_fill_1 FILLER_12_559 ();
 sg13g2_decap_4 FILLER_12_578 ();
 sg13g2_fill_2 FILLER_12_582 ();
 sg13g2_decap_4 FILLER_12_588 ();
 sg13g2_fill_2 FILLER_12_601 ();
 sg13g2_fill_1 FILLER_12_603 ();
 sg13g2_fill_2 FILLER_12_626 ();
 sg13g2_fill_1 FILLER_12_628 ();
 sg13g2_fill_2 FILLER_12_657 ();
 sg13g2_fill_2 FILLER_12_684 ();
 sg13g2_fill_2 FILLER_12_695 ();
 sg13g2_fill_1 FILLER_12_706 ();
 sg13g2_fill_2 FILLER_12_731 ();
 sg13g2_fill_2 FILLER_12_822 ();
 sg13g2_fill_1 FILLER_12_824 ();
 sg13g2_fill_1 FILLER_12_864 ();
 sg13g2_fill_1 FILLER_12_891 ();
 sg13g2_fill_2 FILLER_12_920 ();
 sg13g2_fill_1 FILLER_12_922 ();
 sg13g2_fill_2 FILLER_12_942 ();
 sg13g2_decap_8 FILLER_12_977 ();
 sg13g2_decap_8 FILLER_12_984 ();
 sg13g2_decap_8 FILLER_12_991 ();
 sg13g2_decap_8 FILLER_12_998 ();
 sg13g2_decap_8 FILLER_12_1005 ();
 sg13g2_decap_8 FILLER_12_1012 ();
 sg13g2_decap_8 FILLER_12_1019 ();
 sg13g2_fill_2 FILLER_12_1026 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_fill_2 FILLER_13_50 ();
 sg13g2_fill_1 FILLER_13_52 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_100 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_fill_2 FILLER_13_152 ();
 sg13g2_fill_1 FILLER_13_214 ();
 sg13g2_fill_2 FILLER_13_230 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_fill_1 FILLER_13_306 ();
 sg13g2_fill_2 FILLER_13_315 ();
 sg13g2_fill_1 FILLER_13_317 ();
 sg13g2_decap_4 FILLER_13_351 ();
 sg13g2_fill_1 FILLER_13_355 ();
 sg13g2_fill_1 FILLER_13_449 ();
 sg13g2_fill_1 FILLER_13_490 ();
 sg13g2_fill_2 FILLER_13_508 ();
 sg13g2_fill_2 FILLER_13_541 ();
 sg13g2_fill_1 FILLER_13_547 ();
 sg13g2_fill_2 FILLER_13_584 ();
 sg13g2_fill_1 FILLER_13_601 ();
 sg13g2_fill_2 FILLER_13_619 ();
 sg13g2_fill_1 FILLER_13_621 ();
 sg13g2_fill_2 FILLER_13_645 ();
 sg13g2_fill_1 FILLER_13_647 ();
 sg13g2_fill_1 FILLER_13_662 ();
 sg13g2_fill_1 FILLER_13_675 ();
 sg13g2_decap_4 FILLER_13_738 ();
 sg13g2_fill_1 FILLER_13_742 ();
 sg13g2_fill_2 FILLER_13_767 ();
 sg13g2_fill_1 FILLER_13_778 ();
 sg13g2_fill_2 FILLER_13_798 ();
 sg13g2_fill_2 FILLER_13_815 ();
 sg13g2_fill_2 FILLER_13_825 ();
 sg13g2_fill_1 FILLER_13_827 ();
 sg13g2_fill_1 FILLER_13_841 ();
 sg13g2_fill_2 FILLER_13_895 ();
 sg13g2_decap_8 FILLER_13_977 ();
 sg13g2_decap_8 FILLER_13_984 ();
 sg13g2_decap_8 FILLER_13_991 ();
 sg13g2_decap_8 FILLER_13_998 ();
 sg13g2_decap_8 FILLER_13_1005 ();
 sg13g2_decap_8 FILLER_13_1012 ();
 sg13g2_decap_8 FILLER_13_1019 ();
 sg13g2_fill_2 FILLER_13_1026 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_fill_2 FILLER_14_8 ();
 sg13g2_fill_1 FILLER_14_10 ();
 sg13g2_fill_2 FILLER_14_15 ();
 sg13g2_fill_2 FILLER_14_47 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_68 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_101 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_fill_2 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_decap_4 FILLER_14_258 ();
 sg13g2_fill_2 FILLER_14_266 ();
 sg13g2_fill_2 FILLER_14_272 ();
 sg13g2_fill_1 FILLER_14_274 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_fill_2 FILLER_14_354 ();
 sg13g2_fill_2 FILLER_14_373 ();
 sg13g2_fill_2 FILLER_14_415 ();
 sg13g2_fill_1 FILLER_14_417 ();
 sg13g2_fill_1 FILLER_14_428 ();
 sg13g2_fill_2 FILLER_14_437 ();
 sg13g2_fill_1 FILLER_14_439 ();
 sg13g2_fill_1 FILLER_14_491 ();
 sg13g2_decap_4 FILLER_14_502 ();
 sg13g2_fill_1 FILLER_14_506 ();
 sg13g2_fill_2 FILLER_14_554 ();
 sg13g2_fill_1 FILLER_14_585 ();
 sg13g2_fill_1 FILLER_14_614 ();
 sg13g2_fill_1 FILLER_14_662 ();
 sg13g2_fill_2 FILLER_14_708 ();
 sg13g2_fill_1 FILLER_14_726 ();
 sg13g2_fill_2 FILLER_14_747 ();
 sg13g2_fill_2 FILLER_14_791 ();
 sg13g2_fill_1 FILLER_14_819 ();
 sg13g2_fill_1 FILLER_14_837 ();
 sg13g2_fill_1 FILLER_14_856 ();
 sg13g2_fill_1 FILLER_14_906 ();
 sg13g2_fill_1 FILLER_14_921 ();
 sg13g2_decap_8 FILLER_14_983 ();
 sg13g2_decap_8 FILLER_14_990 ();
 sg13g2_decap_8 FILLER_14_997 ();
 sg13g2_decap_8 FILLER_14_1004 ();
 sg13g2_decap_8 FILLER_14_1011 ();
 sg13g2_decap_8 FILLER_14_1018 ();
 sg13g2_decap_4 FILLER_14_1025 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_fill_2 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_75 ();
 sg13g2_fill_2 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_decap_4 FILLER_15_113 ();
 sg13g2_fill_2 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_143 ();
 sg13g2_decap_4 FILLER_15_251 ();
 sg13g2_fill_2 FILLER_15_255 ();
 sg13g2_fill_1 FILLER_15_317 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_fill_2 FILLER_15_410 ();
 sg13g2_fill_1 FILLER_15_428 ();
 sg13g2_fill_1 FILLER_15_434 ();
 sg13g2_fill_2 FILLER_15_445 ();
 sg13g2_fill_1 FILLER_15_447 ();
 sg13g2_fill_1 FILLER_15_475 ();
 sg13g2_fill_1 FILLER_15_487 ();
 sg13g2_fill_1 FILLER_15_495 ();
 sg13g2_fill_2 FILLER_15_506 ();
 sg13g2_fill_1 FILLER_15_540 ();
 sg13g2_fill_2 FILLER_15_561 ();
 sg13g2_fill_1 FILLER_15_603 ();
 sg13g2_fill_2 FILLER_15_633 ();
 sg13g2_fill_1 FILLER_15_635 ();
 sg13g2_fill_1 FILLER_15_663 ();
 sg13g2_fill_1 FILLER_15_688 ();
 sg13g2_fill_2 FILLER_15_697 ();
 sg13g2_fill_1 FILLER_15_729 ();
 sg13g2_fill_2 FILLER_15_802 ();
 sg13g2_fill_1 FILLER_15_829 ();
 sg13g2_fill_1 FILLER_15_896 ();
 sg13g2_fill_2 FILLER_15_910 ();
 sg13g2_fill_1 FILLER_15_912 ();
 sg13g2_decap_8 FILLER_15_917 ();
 sg13g2_fill_1 FILLER_15_929 ();
 sg13g2_fill_2 FILLER_15_935 ();
 sg13g2_fill_1 FILLER_15_937 ();
 sg13g2_fill_1 FILLER_15_943 ();
 sg13g2_decap_8 FILLER_15_967 ();
 sg13g2_decap_8 FILLER_15_974 ();
 sg13g2_decap_8 FILLER_15_981 ();
 sg13g2_decap_8 FILLER_15_988 ();
 sg13g2_decap_8 FILLER_15_995 ();
 sg13g2_decap_8 FILLER_15_1002 ();
 sg13g2_decap_8 FILLER_15_1009 ();
 sg13g2_decap_8 FILLER_15_1016 ();
 sg13g2_decap_4 FILLER_15_1023 ();
 sg13g2_fill_2 FILLER_15_1027 ();
 sg13g2_fill_1 FILLER_16_12 ();
 sg13g2_decap_4 FILLER_16_71 ();
 sg13g2_fill_2 FILLER_16_75 ();
 sg13g2_fill_1 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_1 FILLER_16_187 ();
 sg13g2_decap_8 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_250 ();
 sg13g2_fill_2 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_293 ();
 sg13g2_fill_1 FILLER_16_317 ();
 sg13g2_fill_1 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_385 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_4 FILLER_16_417 ();
 sg13g2_decap_4 FILLER_16_437 ();
 sg13g2_fill_2 FILLER_16_455 ();
 sg13g2_decap_4 FILLER_16_467 ();
 sg13g2_fill_1 FILLER_16_480 ();
 sg13g2_fill_2 FILLER_16_505 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_fill_2 FILLER_16_522 ();
 sg13g2_fill_1 FILLER_16_571 ();
 sg13g2_fill_2 FILLER_16_581 ();
 sg13g2_fill_1 FILLER_16_583 ();
 sg13g2_fill_2 FILLER_16_590 ();
 sg13g2_fill_1 FILLER_16_592 ();
 sg13g2_fill_1 FILLER_16_631 ();
 sg13g2_fill_2 FILLER_16_655 ();
 sg13g2_fill_1 FILLER_16_722 ();
 sg13g2_decap_8 FILLER_16_747 ();
 sg13g2_fill_1 FILLER_16_754 ();
 sg13g2_fill_2 FILLER_16_768 ();
 sg13g2_fill_1 FILLER_16_780 ();
 sg13g2_fill_2 FILLER_16_831 ();
 sg13g2_fill_1 FILLER_16_879 ();
 sg13g2_fill_2 FILLER_16_910 ();
 sg13g2_fill_1 FILLER_16_912 ();
 sg13g2_fill_2 FILLER_16_926 ();
 sg13g2_fill_1 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_976 ();
 sg13g2_decap_8 FILLER_16_983 ();
 sg13g2_decap_8 FILLER_16_990 ();
 sg13g2_decap_8 FILLER_16_997 ();
 sg13g2_decap_8 FILLER_16_1004 ();
 sg13g2_decap_8 FILLER_16_1011 ();
 sg13g2_decap_8 FILLER_16_1018 ();
 sg13g2_decap_4 FILLER_16_1025 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_60 ();
 sg13g2_fill_2 FILLER_17_79 ();
 sg13g2_fill_1 FILLER_17_81 ();
 sg13g2_decap_8 FILLER_17_99 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_137 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_fill_2 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_246 ();
 sg13g2_fill_2 FILLER_17_307 ();
 sg13g2_fill_1 FILLER_17_326 ();
 sg13g2_fill_1 FILLER_17_337 ();
 sg13g2_fill_2 FILLER_17_360 ();
 sg13g2_fill_1 FILLER_17_362 ();
 sg13g2_fill_1 FILLER_17_404 ();
 sg13g2_decap_4 FILLER_17_419 ();
 sg13g2_fill_2 FILLER_17_423 ();
 sg13g2_decap_4 FILLER_17_457 ();
 sg13g2_fill_2 FILLER_17_499 ();
 sg13g2_fill_1 FILLER_17_516 ();
 sg13g2_fill_2 FILLER_17_548 ();
 sg13g2_fill_1 FILLER_17_550 ();
 sg13g2_fill_1 FILLER_17_566 ();
 sg13g2_fill_2 FILLER_17_582 ();
 sg13g2_decap_8 FILLER_17_591 ();
 sg13g2_fill_1 FILLER_17_598 ();
 sg13g2_fill_1 FILLER_17_634 ();
 sg13g2_fill_2 FILLER_17_643 ();
 sg13g2_decap_4 FILLER_17_661 ();
 sg13g2_fill_1 FILLER_17_684 ();
 sg13g2_decap_4 FILLER_17_709 ();
 sg13g2_fill_1 FILLER_17_733 ();
 sg13g2_fill_1 FILLER_17_852 ();
 sg13g2_fill_1 FILLER_17_868 ();
 sg13g2_fill_2 FILLER_17_878 ();
 sg13g2_fill_1 FILLER_17_890 ();
 sg13g2_fill_2 FILLER_17_930 ();
 sg13g2_fill_2 FILLER_17_940 ();
 sg13g2_decap_8 FILLER_17_969 ();
 sg13g2_decap_8 FILLER_17_976 ();
 sg13g2_decap_8 FILLER_17_983 ();
 sg13g2_decap_8 FILLER_17_990 ();
 sg13g2_decap_8 FILLER_17_997 ();
 sg13g2_decap_8 FILLER_17_1004 ();
 sg13g2_decap_8 FILLER_17_1011 ();
 sg13g2_decap_8 FILLER_17_1018 ();
 sg13g2_decap_4 FILLER_17_1025 ();
 sg13g2_fill_2 FILLER_18_8 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_142 ();
 sg13g2_fill_2 FILLER_18_210 ();
 sg13g2_fill_1 FILLER_18_212 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_262 ();
 sg13g2_fill_1 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_284 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_366 ();
 sg13g2_fill_1 FILLER_18_368 ();
 sg13g2_fill_2 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_405 ();
 sg13g2_fill_1 FILLER_18_412 ();
 sg13g2_decap_8 FILLER_18_426 ();
 sg13g2_fill_1 FILLER_18_433 ();
 sg13g2_decap_4 FILLER_18_438 ();
 sg13g2_fill_1 FILLER_18_442 ();
 sg13g2_fill_2 FILLER_18_484 ();
 sg13g2_fill_1 FILLER_18_486 ();
 sg13g2_fill_2 FILLER_18_507 ();
 sg13g2_fill_2 FILLER_18_551 ();
 sg13g2_fill_2 FILLER_18_586 ();
 sg13g2_fill_1 FILLER_18_642 ();
 sg13g2_decap_8 FILLER_18_710 ();
 sg13g2_decap_4 FILLER_18_740 ();
 sg13g2_fill_2 FILLER_18_791 ();
 sg13g2_fill_2 FILLER_18_817 ();
 sg13g2_fill_2 FILLER_18_927 ();
 sg13g2_fill_1 FILLER_18_929 ();
 sg13g2_decap_8 FILLER_18_978 ();
 sg13g2_decap_8 FILLER_18_985 ();
 sg13g2_decap_8 FILLER_18_992 ();
 sg13g2_decap_8 FILLER_18_999 ();
 sg13g2_decap_8 FILLER_18_1006 ();
 sg13g2_decap_8 FILLER_18_1013 ();
 sg13g2_decap_8 FILLER_18_1020 ();
 sg13g2_fill_2 FILLER_18_1027 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_43 ();
 sg13g2_fill_1 FILLER_19_45 ();
 sg13g2_fill_2 FILLER_19_82 ();
 sg13g2_fill_1 FILLER_19_112 ();
 sg13g2_fill_1 FILLER_19_192 ();
 sg13g2_fill_2 FILLER_19_196 ();
 sg13g2_fill_2 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_fill_2 FILLER_19_340 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_decap_4 FILLER_19_380 ();
 sg13g2_fill_2 FILLER_19_384 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_4 FILLER_19_483 ();
 sg13g2_fill_1 FILLER_19_487 ();
 sg13g2_fill_2 FILLER_19_496 ();
 sg13g2_fill_1 FILLER_19_540 ();
 sg13g2_fill_2 FILLER_19_576 ();
 sg13g2_fill_1 FILLER_19_578 ();
 sg13g2_fill_2 FILLER_19_681 ();
 sg13g2_fill_1 FILLER_19_711 ();
 sg13g2_fill_1 FILLER_19_748 ();
 sg13g2_fill_2 FILLER_19_764 ();
 sg13g2_fill_1 FILLER_19_825 ();
 sg13g2_fill_2 FILLER_19_857 ();
 sg13g2_fill_1 FILLER_19_867 ();
 sg13g2_fill_2 FILLER_19_896 ();
 sg13g2_decap_8 FILLER_19_969 ();
 sg13g2_decap_8 FILLER_19_976 ();
 sg13g2_decap_8 FILLER_19_983 ();
 sg13g2_decap_8 FILLER_19_990 ();
 sg13g2_decap_8 FILLER_19_997 ();
 sg13g2_decap_8 FILLER_19_1004 ();
 sg13g2_decap_8 FILLER_19_1011 ();
 sg13g2_decap_8 FILLER_19_1018 ();
 sg13g2_decap_4 FILLER_19_1025 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_2 FILLER_20_10 ();
 sg13g2_fill_2 FILLER_20_36 ();
 sg13g2_decap_8 FILLER_20_79 ();
 sg13g2_fill_2 FILLER_20_111 ();
 sg13g2_fill_2 FILLER_20_132 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_180 ();
 sg13g2_decap_4 FILLER_20_199 ();
 sg13g2_fill_2 FILLER_20_259 ();
 sg13g2_decap_4 FILLER_20_285 ();
 sg13g2_fill_2 FILLER_20_297 ();
 sg13g2_fill_1 FILLER_20_299 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_fill_2 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_363 ();
 sg13g2_fill_1 FILLER_20_422 ();
 sg13g2_decap_4 FILLER_20_454 ();
 sg13g2_fill_1 FILLER_20_458 ();
 sg13g2_fill_1 FILLER_20_480 ();
 sg13g2_fill_2 FILLER_20_517 ();
 sg13g2_fill_1 FILLER_20_569 ();
 sg13g2_fill_2 FILLER_20_596 ();
 sg13g2_fill_1 FILLER_20_598 ();
 sg13g2_fill_2 FILLER_20_627 ();
 sg13g2_decap_4 FILLER_20_642 ();
 sg13g2_fill_1 FILLER_20_646 ();
 sg13g2_fill_2 FILLER_20_691 ();
 sg13g2_fill_1 FILLER_20_693 ();
 sg13g2_fill_1 FILLER_20_721 ();
 sg13g2_fill_1 FILLER_20_726 ();
 sg13g2_decap_8 FILLER_20_741 ();
 sg13g2_fill_2 FILLER_20_748 ();
 sg13g2_fill_1 FILLER_20_802 ();
 sg13g2_fill_2 FILLER_20_816 ();
 sg13g2_fill_2 FILLER_20_831 ();
 sg13g2_fill_1 FILLER_20_833 ();
 sg13g2_fill_2 FILLER_20_847 ();
 sg13g2_fill_1 FILLER_20_849 ();
 sg13g2_fill_1 FILLER_20_886 ();
 sg13g2_fill_2 FILLER_20_901 ();
 sg13g2_fill_1 FILLER_20_910 ();
 sg13g2_decap_8 FILLER_20_986 ();
 sg13g2_decap_8 FILLER_20_993 ();
 sg13g2_decap_8 FILLER_20_1000 ();
 sg13g2_decap_8 FILLER_20_1007 ();
 sg13g2_decap_8 FILLER_20_1014 ();
 sg13g2_decap_8 FILLER_20_1021 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_fill_2 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_153 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_decap_8 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_fill_2 FILLER_21_247 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_277 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_fill_2 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_367 ();
 sg13g2_fill_2 FILLER_21_430 ();
 sg13g2_fill_1 FILLER_21_432 ();
 sg13g2_decap_8 FILLER_21_451 ();
 sg13g2_fill_1 FILLER_21_458 ();
 sg13g2_decap_8 FILLER_21_505 ();
 sg13g2_decap_4 FILLER_21_525 ();
 sg13g2_fill_2 FILLER_21_555 ();
 sg13g2_fill_1 FILLER_21_557 ();
 sg13g2_fill_2 FILLER_21_666 ();
 sg13g2_fill_2 FILLER_21_675 ();
 sg13g2_fill_1 FILLER_21_677 ();
 sg13g2_decap_4 FILLER_21_703 ();
 sg13g2_fill_2 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_743 ();
 sg13g2_fill_2 FILLER_21_750 ();
 sg13g2_fill_1 FILLER_21_752 ();
 sg13g2_decap_4 FILLER_21_775 ();
 sg13g2_fill_2 FILLER_21_779 ();
 sg13g2_fill_2 FILLER_21_841 ();
 sg13g2_fill_2 FILLER_21_867 ();
 sg13g2_fill_2 FILLER_21_937 ();
 sg13g2_fill_1 FILLER_21_939 ();
 sg13g2_decap_8 FILLER_21_970 ();
 sg13g2_decap_8 FILLER_21_977 ();
 sg13g2_decap_8 FILLER_21_984 ();
 sg13g2_decap_8 FILLER_21_991 ();
 sg13g2_decap_8 FILLER_21_998 ();
 sg13g2_decap_8 FILLER_21_1005 ();
 sg13g2_decap_8 FILLER_21_1012 ();
 sg13g2_decap_8 FILLER_21_1019 ();
 sg13g2_fill_2 FILLER_21_1026 ();
 sg13g2_fill_1 FILLER_21_1028 ();
 sg13g2_fill_2 FILLER_22_8 ();
 sg13g2_fill_1 FILLER_22_40 ();
 sg13g2_decap_4 FILLER_22_51 ();
 sg13g2_decap_4 FILLER_22_88 ();
 sg13g2_fill_2 FILLER_22_92 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_decap_4 FILLER_22_278 ();
 sg13g2_fill_1 FILLER_22_346 ();
 sg13g2_fill_1 FILLER_22_360 ();
 sg13g2_fill_2 FILLER_22_438 ();
 sg13g2_fill_1 FILLER_22_468 ();
 sg13g2_decap_8 FILLER_22_506 ();
 sg13g2_fill_1 FILLER_22_513 ();
 sg13g2_decap_8 FILLER_22_527 ();
 sg13g2_fill_2 FILLER_22_534 ();
 sg13g2_fill_1 FILLER_22_539 ();
 sg13g2_decap_4 FILLER_22_571 ();
 sg13g2_fill_1 FILLER_22_575 ();
 sg13g2_decap_8 FILLER_22_589 ();
 sg13g2_fill_1 FILLER_22_596 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_4 FILLER_22_679 ();
 sg13g2_fill_2 FILLER_22_683 ();
 sg13g2_fill_1 FILLER_22_747 ();
 sg13g2_fill_2 FILLER_22_776 ();
 sg13g2_fill_1 FILLER_22_778 ();
 sg13g2_fill_2 FILLER_22_784 ();
 sg13g2_fill_2 FILLER_22_814 ();
 sg13g2_fill_1 FILLER_22_816 ();
 sg13g2_fill_2 FILLER_22_850 ();
 sg13g2_fill_1 FILLER_22_852 ();
 sg13g2_fill_2 FILLER_22_862 ();
 sg13g2_fill_1 FILLER_22_864 ();
 sg13g2_decap_8 FILLER_22_870 ();
 sg13g2_decap_4 FILLER_22_891 ();
 sg13g2_fill_1 FILLER_22_895 ();
 sg13g2_fill_2 FILLER_22_905 ();
 sg13g2_fill_1 FILLER_22_907 ();
 sg13g2_fill_2 FILLER_22_930 ();
 sg13g2_decap_8 FILLER_22_972 ();
 sg13g2_decap_8 FILLER_22_979 ();
 sg13g2_decap_8 FILLER_22_986 ();
 sg13g2_decap_8 FILLER_22_993 ();
 sg13g2_decap_8 FILLER_22_1000 ();
 sg13g2_decap_8 FILLER_22_1007 ();
 sg13g2_decap_8 FILLER_22_1014 ();
 sg13g2_decap_8 FILLER_22_1021 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_13 ();
 sg13g2_decap_4 FILLER_23_20 ();
 sg13g2_fill_2 FILLER_23_24 ();
 sg13g2_fill_2 FILLER_23_36 ();
 sg13g2_decap_8 FILLER_23_58 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_89 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_132 ();
 sg13g2_fill_2 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_196 ();
 sg13g2_fill_2 FILLER_23_209 ();
 sg13g2_fill_1 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_2 FILLER_23_257 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_fill_1 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_311 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_fill_1 FILLER_23_332 ();
 sg13g2_fill_1 FILLER_23_350 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_1 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_448 ();
 sg13g2_fill_2 FILLER_23_473 ();
 sg13g2_fill_1 FILLER_23_475 ();
 sg13g2_decap_8 FILLER_23_522 ();
 sg13g2_fill_2 FILLER_23_534 ();
 sg13g2_fill_2 FILLER_23_568 ();
 sg13g2_fill_2 FILLER_23_575 ();
 sg13g2_fill_1 FILLER_23_722 ();
 sg13g2_fill_2 FILLER_23_736 ();
 sg13g2_decap_4 FILLER_23_746 ();
 sg13g2_fill_1 FILLER_23_750 ();
 sg13g2_fill_1 FILLER_23_766 ();
 sg13g2_fill_2 FILLER_23_854 ();
 sg13g2_fill_1 FILLER_23_856 ();
 sg13g2_fill_2 FILLER_23_919 ();
 sg13g2_fill_2 FILLER_23_951 ();
 sg13g2_fill_1 FILLER_23_953 ();
 sg13g2_decap_8 FILLER_23_982 ();
 sg13g2_decap_8 FILLER_23_989 ();
 sg13g2_decap_8 FILLER_23_996 ();
 sg13g2_decap_8 FILLER_23_1003 ();
 sg13g2_decap_8 FILLER_23_1010 ();
 sg13g2_decap_8 FILLER_23_1017 ();
 sg13g2_decap_4 FILLER_23_1024 ();
 sg13g2_fill_1 FILLER_23_1028 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_56 ();
 sg13g2_fill_1 FILLER_24_58 ();
 sg13g2_fill_1 FILLER_24_64 ();
 sg13g2_fill_1 FILLER_24_86 ();
 sg13g2_fill_1 FILLER_24_133 ();
 sg13g2_decap_4 FILLER_24_170 ();
 sg13g2_decap_4 FILLER_24_184 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_349 ();
 sg13g2_fill_2 FILLER_24_356 ();
 sg13g2_fill_1 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_fill_1 FILLER_24_403 ();
 sg13g2_fill_1 FILLER_24_472 ();
 sg13g2_fill_1 FILLER_24_488 ();
 sg13g2_fill_1 FILLER_24_494 ();
 sg13g2_fill_1 FILLER_24_558 ();
 sg13g2_fill_2 FILLER_24_568 ();
 sg13g2_fill_1 FILLER_24_570 ();
 sg13g2_fill_1 FILLER_24_628 ();
 sg13g2_fill_1 FILLER_24_634 ();
 sg13g2_fill_1 FILLER_24_653 ();
 sg13g2_fill_2 FILLER_24_673 ();
 sg13g2_fill_2 FILLER_24_715 ();
 sg13g2_fill_2 FILLER_24_742 ();
 sg13g2_fill_1 FILLER_24_744 ();
 sg13g2_decap_8 FILLER_24_755 ();
 sg13g2_decap_8 FILLER_24_762 ();
 sg13g2_decap_4 FILLER_24_769 ();
 sg13g2_decap_8 FILLER_24_803 ();
 sg13g2_decap_4 FILLER_24_810 ();
 sg13g2_fill_1 FILLER_24_840 ();
 sg13g2_fill_2 FILLER_24_855 ();
 sg13g2_fill_1 FILLER_24_857 ();
 sg13g2_decap_8 FILLER_24_883 ();
 sg13g2_fill_2 FILLER_24_916 ();
 sg13g2_fill_1 FILLER_24_918 ();
 sg13g2_fill_1 FILLER_24_928 ();
 sg13g2_fill_1 FILLER_24_939 ();
 sg13g2_fill_2 FILLER_24_945 ();
 sg13g2_fill_1 FILLER_24_947 ();
 sg13g2_decap_8 FILLER_24_970 ();
 sg13g2_decap_8 FILLER_24_977 ();
 sg13g2_decap_8 FILLER_24_984 ();
 sg13g2_decap_8 FILLER_24_991 ();
 sg13g2_decap_8 FILLER_24_998 ();
 sg13g2_decap_8 FILLER_24_1005 ();
 sg13g2_decap_8 FILLER_24_1012 ();
 sg13g2_decap_8 FILLER_24_1019 ();
 sg13g2_fill_2 FILLER_24_1026 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_37 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_fill_2 FILLER_25_62 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_143 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_191 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_fill_2 FILLER_25_204 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_237 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_fill_2 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_fill_1 FILLER_25_433 ();
 sg13g2_fill_2 FILLER_25_447 ();
 sg13g2_fill_2 FILLER_25_474 ();
 sg13g2_fill_1 FILLER_25_476 ();
 sg13g2_fill_1 FILLER_25_535 ();
 sg13g2_fill_2 FILLER_25_614 ();
 sg13g2_fill_1 FILLER_25_616 ();
 sg13g2_fill_2 FILLER_25_680 ();
 sg13g2_fill_1 FILLER_25_682 ();
 sg13g2_fill_1 FILLER_25_692 ();
 sg13g2_fill_2 FILLER_25_715 ();
 sg13g2_fill_2 FILLER_25_738 ();
 sg13g2_decap_4 FILLER_25_745 ();
 sg13g2_fill_1 FILLER_25_764 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_fill_2 FILLER_25_851 ();
 sg13g2_decap_8 FILLER_25_872 ();
 sg13g2_decap_8 FILLER_25_879 ();
 sg13g2_fill_1 FILLER_25_926 ();
 sg13g2_fill_2 FILLER_25_953 ();
 sg13g2_fill_1 FILLER_25_955 ();
 sg13g2_decap_8 FILLER_25_983 ();
 sg13g2_decap_8 FILLER_25_990 ();
 sg13g2_decap_8 FILLER_25_997 ();
 sg13g2_decap_8 FILLER_25_1004 ();
 sg13g2_decap_8 FILLER_25_1011 ();
 sg13g2_decap_8 FILLER_25_1018 ();
 sg13g2_decap_4 FILLER_25_1025 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_34 ();
 sg13g2_fill_2 FILLER_26_48 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_108 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_decap_8 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_157 ();
 sg13g2_decap_8 FILLER_26_185 ();
 sg13g2_decap_8 FILLER_26_192 ();
 sg13g2_decap_4 FILLER_26_208 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_282 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_fill_1 FILLER_26_321 ();
 sg13g2_decap_4 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_361 ();
 sg13g2_fill_2 FILLER_26_367 ();
 sg13g2_fill_2 FILLER_26_384 ();
 sg13g2_fill_1 FILLER_26_411 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_2 FILLER_26_443 ();
 sg13g2_fill_1 FILLER_26_445 ();
 sg13g2_decap_8 FILLER_26_487 ();
 sg13g2_decap_8 FILLER_26_494 ();
 sg13g2_fill_2 FILLER_26_501 ();
 sg13g2_fill_1 FILLER_26_503 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_fill_1 FILLER_26_577 ();
 sg13g2_fill_2 FILLER_26_583 ();
 sg13g2_fill_1 FILLER_26_585 ();
 sg13g2_decap_8 FILLER_26_604 ();
 sg13g2_fill_2 FILLER_26_631 ();
 sg13g2_fill_1 FILLER_26_653 ();
 sg13g2_fill_1 FILLER_26_657 ();
 sg13g2_fill_2 FILLER_26_663 ();
 sg13g2_fill_2 FILLER_26_690 ();
 sg13g2_fill_2 FILLER_26_710 ();
 sg13g2_fill_2 FILLER_26_722 ();
 sg13g2_fill_1 FILLER_26_733 ();
 sg13g2_fill_2 FILLER_26_738 ();
 sg13g2_fill_2 FILLER_26_781 ();
 sg13g2_fill_1 FILLER_26_805 ();
 sg13g2_fill_2 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_867 ();
 sg13g2_fill_2 FILLER_26_874 ();
 sg13g2_fill_1 FILLER_26_876 ();
 sg13g2_fill_1 FILLER_26_890 ();
 sg13g2_decap_8 FILLER_26_981 ();
 sg13g2_decap_8 FILLER_26_988 ();
 sg13g2_decap_8 FILLER_26_995 ();
 sg13g2_decap_8 FILLER_26_1002 ();
 sg13g2_decap_8 FILLER_26_1009 ();
 sg13g2_decap_8 FILLER_26_1016 ();
 sg13g2_decap_4 FILLER_26_1023 ();
 sg13g2_fill_2 FILLER_26_1027 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_decap_8 FILLER_27_58 ();
 sg13g2_decap_4 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_fill_1 FILLER_27_97 ();
 sg13g2_fill_1 FILLER_27_183 ();
 sg13g2_fill_2 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_decap_4 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_327 ();
 sg13g2_fill_2 FILLER_27_346 ();
 sg13g2_fill_1 FILLER_27_361 ();
 sg13g2_fill_2 FILLER_27_410 ();
 sg13g2_fill_1 FILLER_27_412 ();
 sg13g2_fill_1 FILLER_27_446 ();
 sg13g2_fill_1 FILLER_27_460 ();
 sg13g2_fill_2 FILLER_27_476 ();
 sg13g2_fill_1 FILLER_27_495 ();
 sg13g2_decap_8 FILLER_27_536 ();
 sg13g2_decap_8 FILLER_27_543 ();
 sg13g2_fill_1 FILLER_27_563 ();
 sg13g2_fill_2 FILLER_27_603 ();
 sg13g2_decap_8 FILLER_27_641 ();
 sg13g2_fill_2 FILLER_27_691 ();
 sg13g2_fill_1 FILLER_27_693 ();
 sg13g2_fill_1 FILLER_27_717 ();
 sg13g2_fill_1 FILLER_27_738 ();
 sg13g2_fill_2 FILLER_27_744 ();
 sg13g2_fill_1 FILLER_27_746 ();
 sg13g2_fill_1 FILLER_27_786 ();
 sg13g2_fill_2 FILLER_27_811 ();
 sg13g2_fill_2 FILLER_27_839 ();
 sg13g2_fill_1 FILLER_27_875 ();
 sg13g2_fill_2 FILLER_27_942 ();
 sg13g2_decap_8 FILLER_27_971 ();
 sg13g2_decap_8 FILLER_27_978 ();
 sg13g2_decap_8 FILLER_27_985 ();
 sg13g2_decap_8 FILLER_27_992 ();
 sg13g2_decap_8 FILLER_27_999 ();
 sg13g2_decap_8 FILLER_27_1006 ();
 sg13g2_decap_8 FILLER_27_1013 ();
 sg13g2_decap_8 FILLER_27_1020 ();
 sg13g2_fill_2 FILLER_27_1027 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_29 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_fill_2 FILLER_28_100 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_decap_4 FILLER_28_131 ();
 sg13g2_fill_1 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_145 ();
 sg13g2_decap_4 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_fill_2 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_290 ();
 sg13g2_fill_1 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_4 FILLER_28_349 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_fill_2 FILLER_28_417 ();
 sg13g2_fill_1 FILLER_28_419 ();
 sg13g2_fill_2 FILLER_28_459 ();
 sg13g2_fill_2 FILLER_28_495 ();
 sg13g2_fill_1 FILLER_28_510 ();
 sg13g2_decap_8 FILLER_28_545 ();
 sg13g2_fill_2 FILLER_28_552 ();
 sg13g2_fill_2 FILLER_28_584 ();
 sg13g2_fill_1 FILLER_28_599 ();
 sg13g2_fill_1 FILLER_28_603 ();
 sg13g2_fill_1 FILLER_28_617 ();
 sg13g2_fill_2 FILLER_28_651 ();
 sg13g2_fill_1 FILLER_28_668 ();
 sg13g2_fill_2 FILLER_28_674 ();
 sg13g2_fill_1 FILLER_28_676 ();
 sg13g2_fill_1 FILLER_28_784 ();
 sg13g2_decap_4 FILLER_28_836 ();
 sg13g2_fill_2 FILLER_28_840 ();
 sg13g2_fill_2 FILLER_28_874 ();
 sg13g2_fill_2 FILLER_28_894 ();
 sg13g2_fill_1 FILLER_28_896 ();
 sg13g2_fill_2 FILLER_28_911 ();
 sg13g2_fill_2 FILLER_28_953 ();
 sg13g2_decap_8 FILLER_28_976 ();
 sg13g2_decap_8 FILLER_28_983 ();
 sg13g2_decap_8 FILLER_28_990 ();
 sg13g2_decap_8 FILLER_28_997 ();
 sg13g2_decap_8 FILLER_28_1004 ();
 sg13g2_decap_8 FILLER_28_1011 ();
 sg13g2_decap_8 FILLER_28_1018 ();
 sg13g2_decap_4 FILLER_28_1025 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_decap_4 FILLER_29_117 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_decap_4 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_2 FILLER_29_299 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_decap_4 FILLER_29_359 ();
 sg13g2_fill_2 FILLER_29_377 ();
 sg13g2_fill_1 FILLER_29_379 ();
 sg13g2_decap_4 FILLER_29_384 ();
 sg13g2_fill_1 FILLER_29_388 ();
 sg13g2_decap_4 FILLER_29_393 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_29_411 ();
 sg13g2_fill_1 FILLER_29_434 ();
 sg13g2_decap_4 FILLER_29_452 ();
 sg13g2_fill_2 FILLER_29_456 ();
 sg13g2_fill_1 FILLER_29_480 ();
 sg13g2_fill_1 FILLER_29_566 ();
 sg13g2_fill_2 FILLER_29_577 ();
 sg13g2_fill_1 FILLER_29_579 ();
 sg13g2_fill_2 FILLER_29_619 ();
 sg13g2_fill_1 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_702 ();
 sg13g2_decap_8 FILLER_29_709 ();
 sg13g2_decap_4 FILLER_29_716 ();
 sg13g2_fill_2 FILLER_29_730 ();
 sg13g2_fill_1 FILLER_29_732 ();
 sg13g2_fill_1 FILLER_29_739 ();
 sg13g2_fill_2 FILLER_29_769 ();
 sg13g2_fill_1 FILLER_29_780 ();
 sg13g2_decap_8 FILLER_29_802 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_fill_1 FILLER_29_847 ();
 sg13g2_fill_2 FILLER_29_877 ();
 sg13g2_fill_2 FILLER_29_889 ();
 sg13g2_fill_2 FILLER_29_902 ();
 sg13g2_fill_1 FILLER_29_904 ();
 sg13g2_fill_2 FILLER_29_918 ();
 sg13g2_fill_1 FILLER_29_920 ();
 sg13g2_decap_8 FILLER_29_976 ();
 sg13g2_decap_8 FILLER_29_983 ();
 sg13g2_decap_8 FILLER_29_990 ();
 sg13g2_decap_8 FILLER_29_997 ();
 sg13g2_decap_8 FILLER_29_1004 ();
 sg13g2_decap_8 FILLER_29_1011 ();
 sg13g2_decap_8 FILLER_29_1018 ();
 sg13g2_decap_4 FILLER_29_1025 ();
 sg13g2_fill_2 FILLER_30_68 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_160 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_fill_2 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_412 ();
 sg13g2_fill_2 FILLER_30_416 ();
 sg13g2_decap_4 FILLER_30_431 ();
 sg13g2_fill_2 FILLER_30_440 ();
 sg13g2_fill_1 FILLER_30_442 ();
 sg13g2_fill_2 FILLER_30_447 ();
 sg13g2_fill_1 FILLER_30_458 ();
 sg13g2_decap_8 FILLER_30_482 ();
 sg13g2_decap_4 FILLER_30_489 ();
 sg13g2_fill_2 FILLER_30_493 ();
 sg13g2_fill_1 FILLER_30_508 ();
 sg13g2_decap_8 FILLER_30_514 ();
 sg13g2_fill_1 FILLER_30_552 ();
 sg13g2_fill_2 FILLER_30_565 ();
 sg13g2_fill_1 FILLER_30_627 ();
 sg13g2_fill_2 FILLER_30_638 ();
 sg13g2_fill_1 FILLER_30_653 ();
 sg13g2_decap_4 FILLER_30_694 ();
 sg13g2_fill_2 FILLER_30_701 ();
 sg13g2_fill_1 FILLER_30_703 ();
 sg13g2_fill_2 FILLER_30_726 ();
 sg13g2_fill_1 FILLER_30_775 ();
 sg13g2_fill_1 FILLER_30_824 ();
 sg13g2_fill_2 FILLER_30_891 ();
 sg13g2_fill_2 FILLER_30_950 ();
 sg13g2_decap_8 FILLER_30_984 ();
 sg13g2_decap_8 FILLER_30_991 ();
 sg13g2_decap_8 FILLER_30_998 ();
 sg13g2_decap_8 FILLER_30_1005 ();
 sg13g2_decap_8 FILLER_30_1012 ();
 sg13g2_decap_8 FILLER_30_1019 ();
 sg13g2_fill_2 FILLER_30_1026 ();
 sg13g2_fill_1 FILLER_30_1028 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_27 ();
 sg13g2_fill_1 FILLER_31_59 ();
 sg13g2_fill_2 FILLER_31_85 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_104 ();
 sg13g2_fill_1 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_312 ();
 sg13g2_decap_4 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_361 ();
 sg13g2_fill_2 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_375 ();
 sg13g2_fill_2 FILLER_31_410 ();
 sg13g2_fill_1 FILLER_31_509 ();
 sg13g2_fill_2 FILLER_31_536 ();
 sg13g2_fill_2 FILLER_31_577 ();
 sg13g2_fill_1 FILLER_31_579 ();
 sg13g2_fill_1 FILLER_31_585 ();
 sg13g2_fill_2 FILLER_31_602 ();
 sg13g2_fill_1 FILLER_31_740 ();
 sg13g2_fill_2 FILLER_31_816 ();
 sg13g2_decap_4 FILLER_31_855 ();
 sg13g2_fill_2 FILLER_31_874 ();
 sg13g2_fill_1 FILLER_31_876 ();
 sg13g2_fill_1 FILLER_31_887 ();
 sg13g2_fill_1 FILLER_31_911 ();
 sg13g2_decap_8 FILLER_31_982 ();
 sg13g2_decap_8 FILLER_31_989 ();
 sg13g2_decap_8 FILLER_31_996 ();
 sg13g2_decap_8 FILLER_31_1003 ();
 sg13g2_decap_8 FILLER_31_1010 ();
 sg13g2_decap_8 FILLER_31_1017 ();
 sg13g2_decap_4 FILLER_31_1024 ();
 sg13g2_fill_1 FILLER_31_1028 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_fill_1 FILLER_32_86 ();
 sg13g2_decap_8 FILLER_32_113 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_decap_8 FILLER_32_233 ();
 sg13g2_fill_2 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_286 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_313 ();
 sg13g2_fill_2 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_380 ();
 sg13g2_fill_1 FILLER_32_420 ();
 sg13g2_decap_4 FILLER_32_442 ();
 sg13g2_fill_1 FILLER_32_446 ();
 sg13g2_decap_4 FILLER_32_480 ();
 sg13g2_fill_1 FILLER_32_484 ();
 sg13g2_decap_8 FILLER_32_489 ();
 sg13g2_fill_2 FILLER_32_509 ();
 sg13g2_fill_1 FILLER_32_511 ();
 sg13g2_fill_1 FILLER_32_557 ();
 sg13g2_fill_2 FILLER_32_571 ();
 sg13g2_fill_1 FILLER_32_573 ();
 sg13g2_fill_1 FILLER_32_595 ();
 sg13g2_fill_2 FILLER_32_627 ();
 sg13g2_fill_2 FILLER_32_633 ();
 sg13g2_fill_2 FILLER_32_651 ();
 sg13g2_fill_2 FILLER_32_712 ();
 sg13g2_fill_1 FILLER_32_714 ();
 sg13g2_fill_2 FILLER_32_742 ();
 sg13g2_fill_1 FILLER_32_796 ();
 sg13g2_fill_2 FILLER_32_814 ();
 sg13g2_fill_2 FILLER_32_825 ();
 sg13g2_decap_4 FILLER_32_843 ();
 sg13g2_fill_2 FILLER_32_847 ();
 sg13g2_fill_1 FILLER_32_863 ();
 sg13g2_fill_1 FILLER_32_874 ();
 sg13g2_fill_2 FILLER_32_939 ();
 sg13g2_fill_1 FILLER_32_941 ();
 sg13g2_decap_8 FILLER_32_982 ();
 sg13g2_decap_8 FILLER_32_989 ();
 sg13g2_decap_8 FILLER_32_996 ();
 sg13g2_decap_8 FILLER_32_1003 ();
 sg13g2_decap_8 FILLER_32_1010 ();
 sg13g2_decap_8 FILLER_32_1017 ();
 sg13g2_decap_4 FILLER_32_1024 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_29 ();
 sg13g2_fill_1 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_41 ();
 sg13g2_fill_2 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_123 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_138 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_decap_4 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_269 ();
 sg13g2_fill_1 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_decap_4 FILLER_33_412 ();
 sg13g2_fill_1 FILLER_33_416 ();
 sg13g2_fill_1 FILLER_33_445 ();
 sg13g2_fill_2 FILLER_33_469 ();
 sg13g2_fill_2 FILLER_33_474 ();
 sg13g2_fill_1 FILLER_33_476 ();
 sg13g2_fill_2 FILLER_33_507 ();
 sg13g2_fill_2 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_fill_1 FILLER_33_574 ();
 sg13g2_fill_1 FILLER_33_622 ();
 sg13g2_fill_2 FILLER_33_680 ();
 sg13g2_fill_2 FILLER_33_704 ();
 sg13g2_fill_1 FILLER_33_706 ();
 sg13g2_fill_2 FILLER_33_719 ();
 sg13g2_fill_1 FILLER_33_721 ();
 sg13g2_fill_1 FILLER_33_727 ();
 sg13g2_fill_1 FILLER_33_734 ();
 sg13g2_fill_1 FILLER_33_775 ();
 sg13g2_fill_2 FILLER_33_781 ();
 sg13g2_fill_1 FILLER_33_796 ();
 sg13g2_decap_4 FILLER_33_861 ();
 sg13g2_fill_2 FILLER_33_865 ();
 sg13g2_fill_1 FILLER_33_916 ();
 sg13g2_fill_2 FILLER_33_933 ();
 sg13g2_fill_1 FILLER_33_958 ();
 sg13g2_decap_8 FILLER_33_981 ();
 sg13g2_decap_8 FILLER_33_988 ();
 sg13g2_decap_8 FILLER_33_995 ();
 sg13g2_decap_8 FILLER_33_1002 ();
 sg13g2_decap_8 FILLER_33_1009 ();
 sg13g2_decap_8 FILLER_33_1016 ();
 sg13g2_decap_4 FILLER_33_1023 ();
 sg13g2_fill_2 FILLER_33_1027 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_29 ();
 sg13g2_fill_1 FILLER_34_102 ();
 sg13g2_fill_2 FILLER_34_108 ();
 sg13g2_fill_1 FILLER_34_110 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_fill_2 FILLER_34_135 ();
 sg13g2_fill_1 FILLER_34_177 ();
 sg13g2_fill_1 FILLER_34_210 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_243 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_273 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_decap_4 FILLER_34_354 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_440 ();
 sg13g2_fill_2 FILLER_34_457 ();
 sg13g2_fill_2 FILLER_34_473 ();
 sg13g2_fill_1 FILLER_34_503 ();
 sg13g2_fill_2 FILLER_34_542 ();
 sg13g2_fill_1 FILLER_34_636 ();
 sg13g2_fill_1 FILLER_34_650 ();
 sg13g2_fill_1 FILLER_34_713 ();
 sg13g2_fill_1 FILLER_34_719 ();
 sg13g2_fill_1 FILLER_34_757 ();
 sg13g2_fill_1 FILLER_34_805 ();
 sg13g2_fill_2 FILLER_34_814 ();
 sg13g2_fill_2 FILLER_34_841 ();
 sg13g2_fill_1 FILLER_34_843 ();
 sg13g2_fill_1 FILLER_34_895 ();
 sg13g2_fill_2 FILLER_34_961 ();
 sg13g2_fill_1 FILLER_34_963 ();
 sg13g2_decap_8 FILLER_34_977 ();
 sg13g2_decap_8 FILLER_34_984 ();
 sg13g2_decap_8 FILLER_34_991 ();
 sg13g2_decap_8 FILLER_34_998 ();
 sg13g2_decap_8 FILLER_34_1005 ();
 sg13g2_decap_8 FILLER_34_1012 ();
 sg13g2_decap_8 FILLER_34_1019 ();
 sg13g2_fill_2 FILLER_34_1026 ();
 sg13g2_fill_1 FILLER_34_1028 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_10 ();
 sg13g2_fill_2 FILLER_35_41 ();
 sg13g2_fill_2 FILLER_35_53 ();
 sg13g2_fill_1 FILLER_35_55 ();
 sg13g2_fill_2 FILLER_35_61 ();
 sg13g2_fill_2 FILLER_35_85 ();
 sg13g2_fill_2 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_122 ();
 sg13g2_fill_2 FILLER_35_187 ();
 sg13g2_fill_1 FILLER_35_203 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_decap_4 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_decap_4 FILLER_35_329 ();
 sg13g2_fill_2 FILLER_35_392 ();
 sg13g2_fill_1 FILLER_35_394 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_1 FILLER_35_446 ();
 sg13g2_fill_1 FILLER_35_462 ();
 sg13g2_decap_4 FILLER_35_475 ();
 sg13g2_fill_2 FILLER_35_479 ();
 sg13g2_fill_1 FILLER_35_508 ();
 sg13g2_fill_2 FILLER_35_546 ();
 sg13g2_fill_2 FILLER_35_557 ();
 sg13g2_fill_2 FILLER_35_585 ();
 sg13g2_fill_1 FILLER_35_619 ();
 sg13g2_fill_2 FILLER_35_669 ();
 sg13g2_fill_1 FILLER_35_689 ();
 sg13g2_fill_2 FILLER_35_720 ();
 sg13g2_fill_1 FILLER_35_722 ();
 sg13g2_fill_2 FILLER_35_748 ();
 sg13g2_fill_1 FILLER_35_808 ();
 sg13g2_fill_2 FILLER_35_814 ();
 sg13g2_fill_2 FILLER_35_820 ();
 sg13g2_fill_1 FILLER_35_822 ();
 sg13g2_fill_1 FILLER_35_846 ();
 sg13g2_fill_1 FILLER_35_852 ();
 sg13g2_fill_1 FILLER_35_862 ();
 sg13g2_fill_2 FILLER_35_882 ();
 sg13g2_fill_1 FILLER_35_894 ();
 sg13g2_fill_2 FILLER_35_909 ();
 sg13g2_decap_8 FILLER_35_975 ();
 sg13g2_decap_8 FILLER_35_982 ();
 sg13g2_decap_8 FILLER_35_989 ();
 sg13g2_decap_8 FILLER_35_996 ();
 sg13g2_decap_8 FILLER_35_1003 ();
 sg13g2_decap_8 FILLER_35_1010 ();
 sg13g2_decap_8 FILLER_35_1017 ();
 sg13g2_decap_4 FILLER_35_1024 ();
 sg13g2_fill_1 FILLER_35_1028 ();
 sg13g2_fill_1 FILLER_36_76 ();
 sg13g2_fill_2 FILLER_36_115 ();
 sg13g2_fill_1 FILLER_36_136 ();
 sg13g2_fill_1 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_238 ();
 sg13g2_fill_1 FILLER_36_240 ();
 sg13g2_decap_4 FILLER_36_316 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_fill_2 FILLER_36_396 ();
 sg13g2_fill_2 FILLER_36_415 ();
 sg13g2_fill_1 FILLER_36_417 ();
 sg13g2_decap_8 FILLER_36_422 ();
 sg13g2_fill_2 FILLER_36_429 ();
 sg13g2_fill_1 FILLER_36_431 ();
 sg13g2_fill_2 FILLER_36_464 ();
 sg13g2_fill_2 FILLER_36_474 ();
 sg13g2_fill_1 FILLER_36_476 ();
 sg13g2_fill_2 FILLER_36_486 ();
 sg13g2_fill_1 FILLER_36_488 ();
 sg13g2_fill_1 FILLER_36_531 ();
 sg13g2_fill_1 FILLER_36_573 ();
 sg13g2_fill_2 FILLER_36_579 ();
 sg13g2_fill_1 FILLER_36_581 ();
 sg13g2_fill_2 FILLER_36_608 ();
 sg13g2_fill_1 FILLER_36_610 ();
 sg13g2_fill_1 FILLER_36_639 ();
 sg13g2_fill_2 FILLER_36_686 ();
 sg13g2_fill_1 FILLER_36_711 ();
 sg13g2_fill_1 FILLER_36_749 ();
 sg13g2_fill_2 FILLER_36_792 ();
 sg13g2_fill_2 FILLER_36_856 ();
 sg13g2_fill_1 FILLER_36_858 ();
 sg13g2_fill_1 FILLER_36_874 ();
 sg13g2_fill_2 FILLER_36_932 ();
 sg13g2_fill_2 FILLER_36_939 ();
 sg13g2_decap_4 FILLER_36_955 ();
 sg13g2_fill_2 FILLER_36_959 ();
 sg13g2_decap_8 FILLER_36_965 ();
 sg13g2_decap_8 FILLER_36_972 ();
 sg13g2_decap_8 FILLER_36_979 ();
 sg13g2_decap_8 FILLER_36_986 ();
 sg13g2_decap_8 FILLER_36_993 ();
 sg13g2_decap_8 FILLER_36_1000 ();
 sg13g2_decap_8 FILLER_36_1007 ();
 sg13g2_decap_8 FILLER_36_1014 ();
 sg13g2_decap_8 FILLER_36_1021 ();
 sg13g2_fill_1 FILLER_36_1028 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_2 FILLER_37_31 ();
 sg13g2_decap_4 FILLER_37_68 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_fill_2 FILLER_37_146 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_fill_2 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_decap_4 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_307 ();
 sg13g2_decap_4 FILLER_37_317 ();
 sg13g2_fill_2 FILLER_37_334 ();
 sg13g2_fill_1 FILLER_37_336 ();
 sg13g2_fill_2 FILLER_37_429 ();
 sg13g2_fill_2 FILLER_37_478 ();
 sg13g2_fill_2 FILLER_37_517 ();
 sg13g2_fill_1 FILLER_37_519 ();
 sg13g2_fill_2 FILLER_37_530 ();
 sg13g2_fill_1 FILLER_37_532 ();
 sg13g2_fill_1 FILLER_37_598 ();
 sg13g2_fill_1 FILLER_37_639 ();
 sg13g2_decap_4 FILLER_37_695 ();
 sg13g2_fill_2 FILLER_37_729 ();
 sg13g2_fill_1 FILLER_37_744 ();
 sg13g2_fill_2 FILLER_37_798 ();
 sg13g2_fill_1 FILLER_37_800 ();
 sg13g2_fill_2 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_834 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_fill_2 FILLER_37_854 ();
 sg13g2_fill_1 FILLER_37_869 ();
 sg13g2_fill_2 FILLER_37_875 ();
 sg13g2_fill_1 FILLER_37_877 ();
 sg13g2_fill_2 FILLER_37_887 ();
 sg13g2_decap_8 FILLER_37_962 ();
 sg13g2_decap_8 FILLER_37_969 ();
 sg13g2_decap_8 FILLER_37_976 ();
 sg13g2_decap_8 FILLER_37_983 ();
 sg13g2_decap_8 FILLER_37_990 ();
 sg13g2_decap_8 FILLER_37_997 ();
 sg13g2_decap_8 FILLER_37_1004 ();
 sg13g2_decap_8 FILLER_37_1011 ();
 sg13g2_decap_8 FILLER_37_1018 ();
 sg13g2_decap_4 FILLER_37_1025 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_2 FILLER_38_51 ();
 sg13g2_fill_1 FILLER_38_53 ();
 sg13g2_fill_1 FILLER_38_64 ();
 sg13g2_fill_2 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_78 ();
 sg13g2_decap_4 FILLER_38_95 ();
 sg13g2_fill_1 FILLER_38_99 ();
 sg13g2_fill_1 FILLER_38_104 ();
 sg13g2_decap_8 FILLER_38_110 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_decap_4 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_214 ();
 sg13g2_decap_4 FILLER_38_233 ();
 sg13g2_fill_1 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_272 ();
 sg13g2_fill_2 FILLER_38_292 ();
 sg13g2_fill_1 FILLER_38_294 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_2 FILLER_38_389 ();
 sg13g2_fill_1 FILLER_38_407 ();
 sg13g2_fill_2 FILLER_38_418 ();
 sg13g2_decap_4 FILLER_38_502 ();
 sg13g2_fill_2 FILLER_38_506 ();
 sg13g2_fill_1 FILLER_38_568 ();
 sg13g2_fill_2 FILLER_38_587 ();
 sg13g2_decap_4 FILLER_38_677 ();
 sg13g2_fill_2 FILLER_38_729 ();
 sg13g2_fill_1 FILLER_38_731 ();
 sg13g2_fill_2 FILLER_38_760 ();
 sg13g2_fill_2 FILLER_38_767 ();
 sg13g2_fill_2 FILLER_38_796 ();
 sg13g2_decap_4 FILLER_38_850 ();
 sg13g2_fill_2 FILLER_38_854 ();
 sg13g2_fill_1 FILLER_38_879 ();
 sg13g2_decap_4 FILLER_38_936 ();
 sg13g2_decap_8 FILLER_38_944 ();
 sg13g2_decap_8 FILLER_38_951 ();
 sg13g2_decap_8 FILLER_38_958 ();
 sg13g2_decap_8 FILLER_38_965 ();
 sg13g2_decap_8 FILLER_38_972 ();
 sg13g2_decap_8 FILLER_38_979 ();
 sg13g2_decap_8 FILLER_38_986 ();
 sg13g2_decap_8 FILLER_38_993 ();
 sg13g2_decap_8 FILLER_38_1000 ();
 sg13g2_decap_8 FILLER_38_1007 ();
 sg13g2_decap_8 FILLER_38_1014 ();
 sg13g2_decap_8 FILLER_38_1021 ();
 sg13g2_fill_1 FILLER_38_1028 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_30 ();
 sg13g2_fill_2 FILLER_39_71 ();
 sg13g2_fill_1 FILLER_39_73 ();
 sg13g2_fill_1 FILLER_39_84 ();
 sg13g2_fill_2 FILLER_39_106 ();
 sg13g2_decap_8 FILLER_39_138 ();
 sg13g2_decap_8 FILLER_39_145 ();
 sg13g2_decap_4 FILLER_39_163 ();
 sg13g2_fill_2 FILLER_39_167 ();
 sg13g2_fill_2 FILLER_39_181 ();
 sg13g2_fill_2 FILLER_39_199 ();
 sg13g2_fill_1 FILLER_39_227 ();
 sg13g2_fill_1 FILLER_39_241 ();
 sg13g2_fill_2 FILLER_39_293 ();
 sg13g2_decap_4 FILLER_39_333 ();
 sg13g2_fill_2 FILLER_39_350 ();
 sg13g2_fill_1 FILLER_39_352 ();
 sg13g2_fill_1 FILLER_39_363 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_decap_8 FILLER_39_386 ();
 sg13g2_fill_2 FILLER_39_393 ();
 sg13g2_fill_1 FILLER_39_395 ();
 sg13g2_fill_1 FILLER_39_405 ();
 sg13g2_fill_2 FILLER_39_418 ();
 sg13g2_fill_2 FILLER_39_425 ();
 sg13g2_fill_1 FILLER_39_452 ();
 sg13g2_decap_8 FILLER_39_481 ();
 sg13g2_fill_2 FILLER_39_488 ();
 sg13g2_fill_1 FILLER_39_522 ();
 sg13g2_fill_2 FILLER_39_535 ();
 sg13g2_fill_1 FILLER_39_537 ();
 sg13g2_fill_2 FILLER_39_570 ();
 sg13g2_fill_2 FILLER_39_615 ();
 sg13g2_fill_2 FILLER_39_651 ();
 sg13g2_fill_2 FILLER_39_738 ();
 sg13g2_fill_2 FILLER_39_762 ();
 sg13g2_fill_1 FILLER_39_764 ();
 sg13g2_fill_2 FILLER_39_796 ();
 sg13g2_fill_1 FILLER_39_809 ();
 sg13g2_decap_4 FILLER_39_856 ();
 sg13g2_fill_2 FILLER_39_900 ();
 sg13g2_fill_1 FILLER_39_920 ();
 sg13g2_decap_8 FILLER_39_930 ();
 sg13g2_decap_8 FILLER_39_937 ();
 sg13g2_decap_8 FILLER_39_944 ();
 sg13g2_decap_8 FILLER_39_951 ();
 sg13g2_decap_8 FILLER_39_958 ();
 sg13g2_decap_8 FILLER_39_965 ();
 sg13g2_decap_8 FILLER_39_972 ();
 sg13g2_decap_8 FILLER_39_979 ();
 sg13g2_decap_8 FILLER_39_986 ();
 sg13g2_decap_8 FILLER_39_993 ();
 sg13g2_decap_8 FILLER_39_1000 ();
 sg13g2_decap_8 FILLER_39_1007 ();
 sg13g2_decap_8 FILLER_39_1014 ();
 sg13g2_decap_8 FILLER_39_1021 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_fill_2 FILLER_40_54 ();
 sg13g2_fill_2 FILLER_40_65 ();
 sg13g2_fill_1 FILLER_40_67 ();
 sg13g2_decap_8 FILLER_40_82 ();
 sg13g2_fill_2 FILLER_40_89 ();
 sg13g2_fill_1 FILLER_40_104 ();
 sg13g2_decap_4 FILLER_40_127 ();
 sg13g2_fill_1 FILLER_40_131 ();
 sg13g2_decap_4 FILLER_40_145 ();
 sg13g2_fill_1 FILLER_40_149 ();
 sg13g2_fill_1 FILLER_40_157 ();
 sg13g2_decap_4 FILLER_40_168 ();
 sg13g2_fill_1 FILLER_40_198 ();
 sg13g2_fill_1 FILLER_40_263 ();
 sg13g2_fill_1 FILLER_40_269 ();
 sg13g2_fill_1 FILLER_40_302 ();
 sg13g2_fill_2 FILLER_40_327 ();
 sg13g2_fill_2 FILLER_40_333 ();
 sg13g2_fill_1 FILLER_40_335 ();
 sg13g2_fill_2 FILLER_40_340 ();
 sg13g2_fill_1 FILLER_40_342 ();
 sg13g2_fill_2 FILLER_40_358 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_fill_2 FILLER_40_366 ();
 sg13g2_fill_1 FILLER_40_368 ();
 sg13g2_fill_2 FILLER_40_378 ();
 sg13g2_fill_2 FILLER_40_397 ();
 sg13g2_fill_1 FILLER_40_399 ();
 sg13g2_decap_4 FILLER_40_432 ();
 sg13g2_fill_2 FILLER_40_436 ();
 sg13g2_decap_4 FILLER_40_506 ();
 sg13g2_fill_1 FILLER_40_510 ();
 sg13g2_fill_2 FILLER_40_524 ();
 sg13g2_fill_1 FILLER_40_536 ();
 sg13g2_fill_2 FILLER_40_574 ();
 sg13g2_fill_2 FILLER_40_586 ();
 sg13g2_fill_1 FILLER_40_598 ();
 sg13g2_fill_1 FILLER_40_641 ();
 sg13g2_fill_2 FILLER_40_659 ();
 sg13g2_fill_2 FILLER_40_677 ();
 sg13g2_fill_1 FILLER_40_696 ();
 sg13g2_fill_1 FILLER_40_701 ();
 sg13g2_fill_1 FILLER_40_715 ();
 sg13g2_fill_2 FILLER_40_720 ();
 sg13g2_fill_2 FILLER_40_734 ();
 sg13g2_fill_2 FILLER_40_741 ();
 sg13g2_fill_1 FILLER_40_743 ();
 sg13g2_fill_2 FILLER_40_793 ();
 sg13g2_fill_1 FILLER_40_795 ();
 sg13g2_fill_1 FILLER_40_877 ();
 sg13g2_decap_8 FILLER_40_924 ();
 sg13g2_decap_8 FILLER_40_931 ();
 sg13g2_decap_8 FILLER_40_938 ();
 sg13g2_decap_8 FILLER_40_945 ();
 sg13g2_decap_8 FILLER_40_952 ();
 sg13g2_decap_8 FILLER_40_959 ();
 sg13g2_decap_8 FILLER_40_966 ();
 sg13g2_decap_8 FILLER_40_973 ();
 sg13g2_decap_8 FILLER_40_980 ();
 sg13g2_decap_8 FILLER_40_987 ();
 sg13g2_decap_8 FILLER_40_994 ();
 sg13g2_decap_8 FILLER_40_1001 ();
 sg13g2_decap_8 FILLER_40_1008 ();
 sg13g2_decap_8 FILLER_40_1015 ();
 sg13g2_decap_8 FILLER_40_1022 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_4 ();
 sg13g2_fill_1 FILLER_41_12 ();
 sg13g2_fill_2 FILLER_41_67 ();
 sg13g2_fill_1 FILLER_41_69 ();
 sg13g2_fill_2 FILLER_41_80 ();
 sg13g2_fill_1 FILLER_41_87 ();
 sg13g2_fill_2 FILLER_41_93 ();
 sg13g2_fill_1 FILLER_41_95 ();
 sg13g2_fill_1 FILLER_41_101 ();
 sg13g2_fill_2 FILLER_41_141 ();
 sg13g2_fill_1 FILLER_41_203 ();
 sg13g2_fill_2 FILLER_41_251 ();
 sg13g2_fill_1 FILLER_41_253 ();
 sg13g2_fill_1 FILLER_41_265 ();
 sg13g2_fill_2 FILLER_41_290 ();
 sg13g2_fill_2 FILLER_41_302 ();
 sg13g2_fill_2 FILLER_41_325 ();
 sg13g2_fill_2 FILLER_41_331 ();
 sg13g2_fill_1 FILLER_41_333 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_fill_2 FILLER_41_399 ();
 sg13g2_fill_1 FILLER_41_426 ();
 sg13g2_decap_8 FILLER_41_508 ();
 sg13g2_decap_4 FILLER_41_519 ();
 sg13g2_fill_2 FILLER_41_542 ();
 sg13g2_fill_2 FILLER_41_561 ();
 sg13g2_fill_1 FILLER_41_563 ();
 sg13g2_fill_1 FILLER_41_577 ();
 sg13g2_fill_1 FILLER_41_591 ();
 sg13g2_fill_2 FILLER_41_706 ();
 sg13g2_fill_2 FILLER_41_740 ();
 sg13g2_fill_2 FILLER_41_747 ();
 sg13g2_fill_1 FILLER_41_749 ();
 sg13g2_fill_1 FILLER_41_755 ();
 sg13g2_fill_2 FILLER_41_761 ();
 sg13g2_fill_2 FILLER_41_795 ();
 sg13g2_fill_1 FILLER_41_797 ();
 sg13g2_fill_1 FILLER_41_803 ();
 sg13g2_fill_1 FILLER_41_822 ();
 sg13g2_decap_4 FILLER_41_878 ();
 sg13g2_fill_2 FILLER_41_882 ();
 sg13g2_fill_1 FILLER_41_892 ();
 sg13g2_decap_8 FILLER_41_902 ();
 sg13g2_decap_8 FILLER_41_913 ();
 sg13g2_decap_8 FILLER_41_920 ();
 sg13g2_decap_8 FILLER_41_927 ();
 sg13g2_decap_8 FILLER_41_934 ();
 sg13g2_decap_8 FILLER_41_941 ();
 sg13g2_decap_8 FILLER_41_948 ();
 sg13g2_decap_8 FILLER_41_955 ();
 sg13g2_decap_8 FILLER_41_962 ();
 sg13g2_decap_8 FILLER_41_969 ();
 sg13g2_decap_8 FILLER_41_976 ();
 sg13g2_decap_8 FILLER_41_983 ();
 sg13g2_decap_8 FILLER_41_990 ();
 sg13g2_decap_8 FILLER_41_997 ();
 sg13g2_decap_8 FILLER_41_1004 ();
 sg13g2_decap_8 FILLER_41_1011 ();
 sg13g2_decap_8 FILLER_41_1018 ();
 sg13g2_decap_4 FILLER_41_1025 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_2 ();
 sg13g2_fill_1 FILLER_42_31 ();
 sg13g2_fill_1 FILLER_42_71 ();
 sg13g2_fill_2 FILLER_42_88 ();
 sg13g2_decap_4 FILLER_42_95 ();
 sg13g2_fill_2 FILLER_42_99 ();
 sg13g2_fill_1 FILLER_42_106 ();
 sg13g2_decap_4 FILLER_42_139 ();
 sg13g2_fill_1 FILLER_42_143 ();
 sg13g2_fill_1 FILLER_42_151 ();
 sg13g2_fill_1 FILLER_42_178 ();
 sg13g2_fill_2 FILLER_42_240 ();
 sg13g2_fill_1 FILLER_42_324 ();
 sg13g2_fill_1 FILLER_42_356 ();
 sg13g2_fill_2 FILLER_42_371 ();
 sg13g2_fill_1 FILLER_42_373 ();
 sg13g2_fill_1 FILLER_42_398 ();
 sg13g2_decap_4 FILLER_42_403 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_fill_2 FILLER_42_435 ();
 sg13g2_fill_1 FILLER_42_437 ();
 sg13g2_decap_8 FILLER_42_441 ();
 sg13g2_decap_4 FILLER_42_448 ();
 sg13g2_fill_1 FILLER_42_452 ();
 sg13g2_fill_2 FILLER_42_470 ();
 sg13g2_fill_1 FILLER_42_472 ();
 sg13g2_fill_1 FILLER_42_482 ();
 sg13g2_decap_8 FILLER_42_500 ();
 sg13g2_decap_4 FILLER_42_507 ();
 sg13g2_decap_4 FILLER_42_524 ();
 sg13g2_fill_2 FILLER_42_533 ();
 sg13g2_decap_8 FILLER_42_577 ();
 sg13g2_fill_1 FILLER_42_638 ();
 sg13g2_fill_1 FILLER_42_652 ();
 sg13g2_fill_2 FILLER_42_663 ();
 sg13g2_fill_2 FILLER_42_719 ();
 sg13g2_fill_1 FILLER_42_721 ();
 sg13g2_fill_1 FILLER_42_766 ();
 sg13g2_fill_1 FILLER_42_799 ();
 sg13g2_fill_2 FILLER_42_824 ();
 sg13g2_fill_2 FILLER_42_834 ();
 sg13g2_decap_4 FILLER_42_859 ();
 sg13g2_fill_2 FILLER_42_863 ();
 sg13g2_decap_4 FILLER_42_868 ();
 sg13g2_decap_4 FILLER_42_881 ();
 sg13g2_fill_2 FILLER_42_885 ();
 sg13g2_decap_8 FILLER_42_892 ();
 sg13g2_decap_8 FILLER_42_899 ();
 sg13g2_decap_8 FILLER_42_906 ();
 sg13g2_decap_8 FILLER_42_913 ();
 sg13g2_decap_8 FILLER_42_920 ();
 sg13g2_decap_8 FILLER_42_927 ();
 sg13g2_decap_8 FILLER_42_934 ();
 sg13g2_decap_8 FILLER_42_941 ();
 sg13g2_decap_8 FILLER_42_948 ();
 sg13g2_decap_8 FILLER_42_955 ();
 sg13g2_decap_8 FILLER_42_962 ();
 sg13g2_decap_8 FILLER_42_969 ();
 sg13g2_decap_8 FILLER_42_976 ();
 sg13g2_decap_8 FILLER_42_983 ();
 sg13g2_decap_8 FILLER_42_990 ();
 sg13g2_decap_8 FILLER_42_997 ();
 sg13g2_decap_8 FILLER_42_1004 ();
 sg13g2_decap_8 FILLER_42_1011 ();
 sg13g2_decap_8 FILLER_42_1018 ();
 sg13g2_decap_4 FILLER_42_1025 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_31 ();
 sg13g2_fill_1 FILLER_43_33 ();
 sg13g2_fill_1 FILLER_43_61 ();
 sg13g2_fill_2 FILLER_43_66 ();
 sg13g2_fill_2 FILLER_43_75 ();
 sg13g2_fill_2 FILLER_43_82 ();
 sg13g2_fill_2 FILLER_43_158 ();
 sg13g2_fill_1 FILLER_43_160 ();
 sg13g2_fill_1 FILLER_43_171 ();
 sg13g2_fill_2 FILLER_43_182 ();
 sg13g2_fill_2 FILLER_43_208 ();
 sg13g2_fill_1 FILLER_43_227 ();
 sg13g2_fill_1 FILLER_43_256 ();
 sg13g2_fill_2 FILLER_43_292 ();
 sg13g2_decap_4 FILLER_43_304 ();
 sg13g2_fill_1 FILLER_43_308 ();
 sg13g2_fill_2 FILLER_43_322 ();
 sg13g2_fill_1 FILLER_43_389 ();
 sg13g2_decap_4 FILLER_43_450 ();
 sg13g2_decap_4 FILLER_43_495 ();
 sg13g2_fill_2 FILLER_43_516 ();
 sg13g2_fill_2 FILLER_43_550 ();
 sg13g2_fill_2 FILLER_43_602 ();
 sg13g2_fill_1 FILLER_43_604 ();
 sg13g2_fill_2 FILLER_43_617 ();
 sg13g2_fill_1 FILLER_43_629 ();
 sg13g2_fill_2 FILLER_43_639 ();
 sg13g2_fill_1 FILLER_43_659 ();
 sg13g2_fill_1 FILLER_43_710 ();
 sg13g2_decap_8 FILLER_43_823 ();
 sg13g2_decap_8 FILLER_43_830 ();
 sg13g2_decap_8 FILLER_43_837 ();
 sg13g2_decap_4 FILLER_43_844 ();
 sg13g2_fill_2 FILLER_43_848 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_decap_8 FILLER_43_875 ();
 sg13g2_decap_8 FILLER_43_882 ();
 sg13g2_decap_8 FILLER_43_889 ();
 sg13g2_decap_8 FILLER_43_896 ();
 sg13g2_decap_8 FILLER_43_903 ();
 sg13g2_decap_8 FILLER_43_910 ();
 sg13g2_decap_8 FILLER_43_917 ();
 sg13g2_decap_8 FILLER_43_924 ();
 sg13g2_decap_8 FILLER_43_931 ();
 sg13g2_decap_8 FILLER_43_938 ();
 sg13g2_decap_8 FILLER_43_945 ();
 sg13g2_decap_8 FILLER_43_952 ();
 sg13g2_decap_8 FILLER_43_959 ();
 sg13g2_decap_8 FILLER_43_966 ();
 sg13g2_decap_8 FILLER_43_973 ();
 sg13g2_decap_8 FILLER_43_980 ();
 sg13g2_decap_8 FILLER_43_987 ();
 sg13g2_decap_8 FILLER_43_994 ();
 sg13g2_decap_8 FILLER_43_1001 ();
 sg13g2_decap_8 FILLER_43_1008 ();
 sg13g2_decap_8 FILLER_43_1015 ();
 sg13g2_decap_8 FILLER_43_1022 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_13 ();
 sg13g2_fill_2 FILLER_44_20 ();
 sg13g2_fill_1 FILLER_44_22 ();
 sg13g2_fill_1 FILLER_44_37 ();
 sg13g2_fill_2 FILLER_44_68 ();
 sg13g2_fill_1 FILLER_44_70 ();
 sg13g2_fill_2 FILLER_44_86 ();
 sg13g2_fill_2 FILLER_44_106 ();
 sg13g2_fill_1 FILLER_44_108 ();
 sg13g2_fill_2 FILLER_44_113 ();
 sg13g2_fill_1 FILLER_44_115 ();
 sg13g2_fill_1 FILLER_44_178 ();
 sg13g2_fill_1 FILLER_44_233 ();
 sg13g2_fill_1 FILLER_44_238 ();
 sg13g2_fill_1 FILLER_44_306 ();
 sg13g2_fill_2 FILLER_44_379 ();
 sg13g2_fill_2 FILLER_44_398 ();
 sg13g2_fill_1 FILLER_44_400 ();
 sg13g2_fill_1 FILLER_44_411 ();
 sg13g2_fill_2 FILLER_44_419 ();
 sg13g2_fill_2 FILLER_44_438 ();
 sg13g2_fill_1 FILLER_44_481 ();
 sg13g2_fill_1 FILLER_44_496 ();
 sg13g2_decap_8 FILLER_44_502 ();
 sg13g2_decap_8 FILLER_44_509 ();
 sg13g2_fill_2 FILLER_44_516 ();
 sg13g2_decap_4 FILLER_44_553 ();
 sg13g2_decap_8 FILLER_44_561 ();
 sg13g2_decap_4 FILLER_44_568 ();
 sg13g2_fill_1 FILLER_44_664 ();
 sg13g2_fill_2 FILLER_44_698 ();
 sg13g2_fill_2 FILLER_44_733 ();
 sg13g2_fill_1 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_739 ();
 sg13g2_decap_4 FILLER_44_746 ();
 sg13g2_fill_1 FILLER_44_750 ();
 sg13g2_fill_2 FILLER_44_755 ();
 sg13g2_fill_1 FILLER_44_757 ();
 sg13g2_fill_2 FILLER_44_767 ();
 sg13g2_decap_8 FILLER_44_800 ();
 sg13g2_decap_8 FILLER_44_807 ();
 sg13g2_decap_8 FILLER_44_814 ();
 sg13g2_decap_8 FILLER_44_821 ();
 sg13g2_decap_8 FILLER_44_828 ();
 sg13g2_decap_8 FILLER_44_835 ();
 sg13g2_decap_8 FILLER_44_842 ();
 sg13g2_decap_8 FILLER_44_849 ();
 sg13g2_decap_8 FILLER_44_856 ();
 sg13g2_decap_8 FILLER_44_863 ();
 sg13g2_decap_8 FILLER_44_870 ();
 sg13g2_decap_8 FILLER_44_877 ();
 sg13g2_decap_8 FILLER_44_884 ();
 sg13g2_decap_8 FILLER_44_891 ();
 sg13g2_decap_8 FILLER_44_898 ();
 sg13g2_decap_8 FILLER_44_905 ();
 sg13g2_decap_8 FILLER_44_912 ();
 sg13g2_decap_8 FILLER_44_919 ();
 sg13g2_decap_8 FILLER_44_926 ();
 sg13g2_decap_8 FILLER_44_933 ();
 sg13g2_decap_8 FILLER_44_940 ();
 sg13g2_decap_8 FILLER_44_947 ();
 sg13g2_decap_8 FILLER_44_954 ();
 sg13g2_decap_8 FILLER_44_961 ();
 sg13g2_decap_8 FILLER_44_968 ();
 sg13g2_decap_8 FILLER_44_975 ();
 sg13g2_decap_8 FILLER_44_982 ();
 sg13g2_decap_8 FILLER_44_989 ();
 sg13g2_decap_8 FILLER_44_996 ();
 sg13g2_decap_8 FILLER_44_1003 ();
 sg13g2_decap_8 FILLER_44_1010 ();
 sg13g2_decap_8 FILLER_44_1017 ();
 sg13g2_decap_4 FILLER_44_1024 ();
 sg13g2_fill_1 FILLER_44_1028 ();
 sg13g2_decap_4 FILLER_45_42 ();
 sg13g2_decap_4 FILLER_45_56 ();
 sg13g2_fill_2 FILLER_45_106 ();
 sg13g2_fill_2 FILLER_45_113 ();
 sg13g2_fill_2 FILLER_45_148 ();
 sg13g2_fill_1 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_246 ();
 sg13g2_fill_2 FILLER_45_336 ();
 sg13g2_fill_2 FILLER_45_371 ();
 sg13g2_fill_2 FILLER_45_383 ();
 sg13g2_fill_1 FILLER_45_385 ();
 sg13g2_fill_2 FILLER_45_421 ();
 sg13g2_fill_2 FILLER_45_437 ();
 sg13g2_decap_4 FILLER_45_463 ();
 sg13g2_fill_2 FILLER_45_479 ();
 sg13g2_fill_1 FILLER_45_481 ();
 sg13g2_fill_1 FILLER_45_513 ();
 sg13g2_fill_1 FILLER_45_549 ();
 sg13g2_fill_1 FILLER_45_565 ();
 sg13g2_fill_2 FILLER_45_610 ();
 sg13g2_fill_1 FILLER_45_612 ();
 sg13g2_fill_1 FILLER_45_631 ();
 sg13g2_fill_2 FILLER_45_660 ();
 sg13g2_decap_4 FILLER_45_674 ();
 sg13g2_decap_8 FILLER_45_683 ();
 sg13g2_fill_1 FILLER_45_690 ();
 sg13g2_fill_2 FILLER_45_695 ();
 sg13g2_fill_1 FILLER_45_697 ();
 sg13g2_fill_2 FILLER_45_706 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_decap_8 FILLER_45_746 ();
 sg13g2_decap_8 FILLER_45_753 ();
 sg13g2_decap_8 FILLER_45_760 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_fill_1 FILLER_45_777 ();
 sg13g2_fill_2 FILLER_45_788 ();
 sg13g2_fill_1 FILLER_45_790 ();
 sg13g2_decap_8 FILLER_45_795 ();
 sg13g2_decap_8 FILLER_45_802 ();
 sg13g2_decap_8 FILLER_45_809 ();
 sg13g2_decap_8 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_823 ();
 sg13g2_decap_8 FILLER_45_830 ();
 sg13g2_decap_8 FILLER_45_837 ();
 sg13g2_decap_8 FILLER_45_844 ();
 sg13g2_decap_8 FILLER_45_851 ();
 sg13g2_decap_8 FILLER_45_858 ();
 sg13g2_decap_8 FILLER_45_865 ();
 sg13g2_decap_8 FILLER_45_872 ();
 sg13g2_decap_8 FILLER_45_879 ();
 sg13g2_decap_8 FILLER_45_886 ();
 sg13g2_decap_8 FILLER_45_893 ();
 sg13g2_decap_8 FILLER_45_900 ();
 sg13g2_decap_8 FILLER_45_907 ();
 sg13g2_decap_8 FILLER_45_914 ();
 sg13g2_decap_8 FILLER_45_921 ();
 sg13g2_decap_8 FILLER_45_928 ();
 sg13g2_decap_8 FILLER_45_935 ();
 sg13g2_decap_8 FILLER_45_942 ();
 sg13g2_decap_8 FILLER_45_949 ();
 sg13g2_decap_8 FILLER_45_956 ();
 sg13g2_decap_8 FILLER_45_963 ();
 sg13g2_decap_8 FILLER_45_970 ();
 sg13g2_decap_8 FILLER_45_977 ();
 sg13g2_decap_8 FILLER_45_984 ();
 sg13g2_decap_8 FILLER_45_991 ();
 sg13g2_decap_8 FILLER_45_998 ();
 sg13g2_decap_8 FILLER_45_1005 ();
 sg13g2_decap_8 FILLER_45_1012 ();
 sg13g2_decap_8 FILLER_45_1019 ();
 sg13g2_fill_2 FILLER_45_1026 ();
 sg13g2_fill_1 FILLER_45_1028 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_fill_2 FILLER_46_45 ();
 sg13g2_fill_1 FILLER_46_47 ();
 sg13g2_fill_2 FILLER_46_99 ();
 sg13g2_fill_1 FILLER_46_101 ();
 sg13g2_fill_2 FILLER_46_141 ();
 sg13g2_fill_1 FILLER_46_143 ();
 sg13g2_fill_1 FILLER_46_161 ();
 sg13g2_fill_2 FILLER_46_177 ();
 sg13g2_fill_1 FILLER_46_207 ();
 sg13g2_fill_2 FILLER_46_213 ();
 sg13g2_decap_8 FILLER_46_228 ();
 sg13g2_fill_2 FILLER_46_235 ();
 sg13g2_fill_2 FILLER_46_265 ();
 sg13g2_fill_2 FILLER_46_340 ();
 sg13g2_fill_2 FILLER_46_364 ();
 sg13g2_fill_2 FILLER_46_487 ();
 sg13g2_fill_1 FILLER_46_503 ();
 sg13g2_fill_2 FILLER_46_555 ();
 sg13g2_fill_1 FILLER_46_557 ();
 sg13g2_fill_2 FILLER_46_598 ();
 sg13g2_fill_1 FILLER_46_600 ();
 sg13g2_decap_8 FILLER_46_653 ();
 sg13g2_decap_8 FILLER_46_660 ();
 sg13g2_decap_8 FILLER_46_667 ();
 sg13g2_decap_8 FILLER_46_674 ();
 sg13g2_decap_8 FILLER_46_681 ();
 sg13g2_decap_8 FILLER_46_688 ();
 sg13g2_decap_8 FILLER_46_695 ();
 sg13g2_decap_8 FILLER_46_702 ();
 sg13g2_decap_8 FILLER_46_709 ();
 sg13g2_decap_8 FILLER_46_716 ();
 sg13g2_decap_8 FILLER_46_723 ();
 sg13g2_decap_8 FILLER_46_730 ();
 sg13g2_decap_8 FILLER_46_737 ();
 sg13g2_decap_8 FILLER_46_744 ();
 sg13g2_decap_8 FILLER_46_751 ();
 sg13g2_decap_8 FILLER_46_758 ();
 sg13g2_decap_8 FILLER_46_765 ();
 sg13g2_decap_8 FILLER_46_772 ();
 sg13g2_decap_8 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_793 ();
 sg13g2_decap_8 FILLER_46_800 ();
 sg13g2_decap_8 FILLER_46_807 ();
 sg13g2_decap_8 FILLER_46_814 ();
 sg13g2_decap_8 FILLER_46_821 ();
 sg13g2_decap_8 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_835 ();
 sg13g2_decap_8 FILLER_46_842 ();
 sg13g2_decap_8 FILLER_46_849 ();
 sg13g2_decap_8 FILLER_46_856 ();
 sg13g2_decap_8 FILLER_46_863 ();
 sg13g2_decap_8 FILLER_46_870 ();
 sg13g2_decap_8 FILLER_46_877 ();
 sg13g2_decap_8 FILLER_46_884 ();
 sg13g2_decap_8 FILLER_46_891 ();
 sg13g2_decap_8 FILLER_46_898 ();
 sg13g2_decap_8 FILLER_46_905 ();
 sg13g2_decap_8 FILLER_46_912 ();
 sg13g2_decap_8 FILLER_46_919 ();
 sg13g2_decap_8 FILLER_46_926 ();
 sg13g2_decap_8 FILLER_46_933 ();
 sg13g2_decap_8 FILLER_46_940 ();
 sg13g2_decap_8 FILLER_46_947 ();
 sg13g2_decap_8 FILLER_46_954 ();
 sg13g2_decap_8 FILLER_46_961 ();
 sg13g2_decap_8 FILLER_46_968 ();
 sg13g2_decap_8 FILLER_46_975 ();
 sg13g2_decap_8 FILLER_46_982 ();
 sg13g2_decap_8 FILLER_46_989 ();
 sg13g2_decap_8 FILLER_46_996 ();
 sg13g2_decap_8 FILLER_46_1003 ();
 sg13g2_decap_8 FILLER_46_1010 ();
 sg13g2_decap_8 FILLER_46_1017 ();
 sg13g2_decap_4 FILLER_46_1024 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_11 ();
 sg13g2_fill_2 FILLER_47_17 ();
 sg13g2_fill_1 FILLER_47_61 ();
 sg13g2_fill_2 FILLER_47_126 ();
 sg13g2_fill_1 FILLER_47_165 ();
 sg13g2_fill_1 FILLER_47_282 ();
 sg13g2_fill_1 FILLER_47_323 ();
 sg13g2_fill_2 FILLER_47_337 ();
 sg13g2_fill_2 FILLER_47_376 ();
 sg13g2_fill_2 FILLER_47_410 ();
 sg13g2_fill_1 FILLER_47_412 ();
 sg13g2_fill_2 FILLER_47_445 ();
 sg13g2_fill_1 FILLER_47_562 ();
 sg13g2_fill_2 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_591 ();
 sg13g2_decap_8 FILLER_47_598 ();
 sg13g2_fill_1 FILLER_47_605 ();
 sg13g2_decap_8 FILLER_47_610 ();
 sg13g2_decap_8 FILLER_47_617 ();
 sg13g2_decap_4 FILLER_47_624 ();
 sg13g2_decap_4 FILLER_47_632 ();
 sg13g2_fill_1 FILLER_47_636 ();
 sg13g2_decap_8 FILLER_47_641 ();
 sg13g2_decap_8 FILLER_47_648 ();
 sg13g2_decap_8 FILLER_47_655 ();
 sg13g2_decap_8 FILLER_47_662 ();
 sg13g2_decap_8 FILLER_47_669 ();
 sg13g2_decap_8 FILLER_47_676 ();
 sg13g2_decap_8 FILLER_47_683 ();
 sg13g2_decap_8 FILLER_47_690 ();
 sg13g2_decap_8 FILLER_47_697 ();
 sg13g2_decap_8 FILLER_47_704 ();
 sg13g2_decap_8 FILLER_47_711 ();
 sg13g2_decap_8 FILLER_47_718 ();
 sg13g2_decap_8 FILLER_47_725 ();
 sg13g2_decap_8 FILLER_47_732 ();
 sg13g2_decap_8 FILLER_47_739 ();
 sg13g2_decap_8 FILLER_47_746 ();
 sg13g2_decap_8 FILLER_47_753 ();
 sg13g2_decap_8 FILLER_47_760 ();
 sg13g2_decap_8 FILLER_47_767 ();
 sg13g2_decap_8 FILLER_47_774 ();
 sg13g2_decap_8 FILLER_47_781 ();
 sg13g2_decap_8 FILLER_47_788 ();
 sg13g2_decap_8 FILLER_47_795 ();
 sg13g2_decap_8 FILLER_47_802 ();
 sg13g2_decap_8 FILLER_47_809 ();
 sg13g2_decap_8 FILLER_47_816 ();
 sg13g2_decap_8 FILLER_47_823 ();
 sg13g2_decap_8 FILLER_47_830 ();
 sg13g2_decap_8 FILLER_47_837 ();
 sg13g2_decap_8 FILLER_47_844 ();
 sg13g2_decap_8 FILLER_47_851 ();
 sg13g2_decap_8 FILLER_47_858 ();
 sg13g2_decap_8 FILLER_47_865 ();
 sg13g2_decap_8 FILLER_47_872 ();
 sg13g2_decap_8 FILLER_47_879 ();
 sg13g2_decap_8 FILLER_47_886 ();
 sg13g2_decap_8 FILLER_47_893 ();
 sg13g2_decap_8 FILLER_47_900 ();
 sg13g2_decap_8 FILLER_47_907 ();
 sg13g2_decap_8 FILLER_47_914 ();
 sg13g2_decap_8 FILLER_47_921 ();
 sg13g2_decap_8 FILLER_47_928 ();
 sg13g2_decap_8 FILLER_47_935 ();
 sg13g2_decap_8 FILLER_47_942 ();
 sg13g2_decap_8 FILLER_47_949 ();
 sg13g2_decap_8 FILLER_47_956 ();
 sg13g2_decap_8 FILLER_47_963 ();
 sg13g2_decap_8 FILLER_47_970 ();
 sg13g2_decap_8 FILLER_47_977 ();
 sg13g2_decap_8 FILLER_47_984 ();
 sg13g2_decap_8 FILLER_47_991 ();
 sg13g2_decap_8 FILLER_47_998 ();
 sg13g2_decap_8 FILLER_47_1005 ();
 sg13g2_decap_8 FILLER_47_1012 ();
 sg13g2_decap_8 FILLER_47_1019 ();
 sg13g2_fill_2 FILLER_47_1026 ();
 sg13g2_fill_1 FILLER_47_1028 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_fill_1 FILLER_48_21 ();
 sg13g2_fill_2 FILLER_48_159 ();
 sg13g2_fill_1 FILLER_48_166 ();
 sg13g2_decap_8 FILLER_48_232 ();
 sg13g2_fill_1 FILLER_48_239 ();
 sg13g2_fill_1 FILLER_48_298 ();
 sg13g2_fill_2 FILLER_48_332 ();
 sg13g2_fill_1 FILLER_48_334 ();
 sg13g2_fill_1 FILLER_48_423 ();
 sg13g2_fill_1 FILLER_48_464 ();
 sg13g2_decap_8 FILLER_48_562 ();
 sg13g2_fill_2 FILLER_48_569 ();
 sg13g2_decap_8 FILLER_48_575 ();
 sg13g2_decap_8 FILLER_48_582 ();
 sg13g2_decap_8 FILLER_48_589 ();
 sg13g2_decap_8 FILLER_48_596 ();
 sg13g2_decap_8 FILLER_48_603 ();
 sg13g2_decap_8 FILLER_48_610 ();
 sg13g2_decap_8 FILLER_48_617 ();
 sg13g2_decap_8 FILLER_48_624 ();
 sg13g2_decap_8 FILLER_48_631 ();
 sg13g2_decap_8 FILLER_48_638 ();
 sg13g2_decap_8 FILLER_48_645 ();
 sg13g2_decap_8 FILLER_48_652 ();
 sg13g2_decap_8 FILLER_48_659 ();
 sg13g2_decap_8 FILLER_48_666 ();
 sg13g2_decap_8 FILLER_48_673 ();
 sg13g2_decap_8 FILLER_48_680 ();
 sg13g2_decap_8 FILLER_48_687 ();
 sg13g2_decap_8 FILLER_48_694 ();
 sg13g2_decap_8 FILLER_48_701 ();
 sg13g2_decap_8 FILLER_48_708 ();
 sg13g2_decap_8 FILLER_48_715 ();
 sg13g2_decap_8 FILLER_48_722 ();
 sg13g2_decap_8 FILLER_48_729 ();
 sg13g2_decap_8 FILLER_48_736 ();
 sg13g2_decap_8 FILLER_48_743 ();
 sg13g2_decap_8 FILLER_48_750 ();
 sg13g2_decap_8 FILLER_48_757 ();
 sg13g2_decap_8 FILLER_48_764 ();
 sg13g2_decap_8 FILLER_48_771 ();
 sg13g2_decap_8 FILLER_48_778 ();
 sg13g2_decap_8 FILLER_48_785 ();
 sg13g2_decap_8 FILLER_48_792 ();
 sg13g2_decap_8 FILLER_48_799 ();
 sg13g2_decap_8 FILLER_48_806 ();
 sg13g2_decap_8 FILLER_48_813 ();
 sg13g2_decap_8 FILLER_48_820 ();
 sg13g2_decap_8 FILLER_48_827 ();
 sg13g2_decap_8 FILLER_48_834 ();
 sg13g2_decap_8 FILLER_48_841 ();
 sg13g2_decap_8 FILLER_48_848 ();
 sg13g2_decap_8 FILLER_48_855 ();
 sg13g2_decap_8 FILLER_48_862 ();
 sg13g2_decap_8 FILLER_48_869 ();
 sg13g2_decap_8 FILLER_48_876 ();
 sg13g2_decap_8 FILLER_48_883 ();
 sg13g2_decap_8 FILLER_48_890 ();
 sg13g2_decap_8 FILLER_48_897 ();
 sg13g2_decap_8 FILLER_48_904 ();
 sg13g2_decap_8 FILLER_48_911 ();
 sg13g2_decap_8 FILLER_48_918 ();
 sg13g2_decap_8 FILLER_48_925 ();
 sg13g2_decap_8 FILLER_48_932 ();
 sg13g2_decap_8 FILLER_48_939 ();
 sg13g2_decap_8 FILLER_48_946 ();
 sg13g2_decap_8 FILLER_48_953 ();
 sg13g2_decap_8 FILLER_48_960 ();
 sg13g2_decap_8 FILLER_48_967 ();
 sg13g2_decap_8 FILLER_48_974 ();
 sg13g2_decap_8 FILLER_48_981 ();
 sg13g2_decap_8 FILLER_48_988 ();
 sg13g2_decap_8 FILLER_48_995 ();
 sg13g2_decap_8 FILLER_48_1002 ();
 sg13g2_decap_8 FILLER_48_1009 ();
 sg13g2_decap_8 FILLER_48_1016 ();
 sg13g2_decap_4 FILLER_48_1023 ();
 sg13g2_fill_2 FILLER_48_1027 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_1 FILLER_49_21 ();
 sg13g2_fill_2 FILLER_49_134 ();
 sg13g2_fill_1 FILLER_49_161 ();
 sg13g2_fill_1 FILLER_49_172 ();
 sg13g2_fill_2 FILLER_49_195 ();
 sg13g2_fill_1 FILLER_49_205 ();
 sg13g2_decap_8 FILLER_49_219 ();
 sg13g2_decap_8 FILLER_49_226 ();
 sg13g2_decap_8 FILLER_49_233 ();
 sg13g2_decap_8 FILLER_49_240 ();
 sg13g2_fill_1 FILLER_49_277 ();
 sg13g2_fill_1 FILLER_49_301 ();
 sg13g2_fill_1 FILLER_49_315 ();
 sg13g2_fill_1 FILLER_49_378 ();
 sg13g2_fill_1 FILLER_49_392 ();
 sg13g2_fill_2 FILLER_49_440 ();
 sg13g2_decap_4 FILLER_49_455 ();
 sg13g2_fill_2 FILLER_49_459 ();
 sg13g2_decap_8 FILLER_49_465 ();
 sg13g2_fill_1 FILLER_49_472 ();
 sg13g2_fill_2 FILLER_49_481 ();
 sg13g2_fill_1 FILLER_49_483 ();
 sg13g2_fill_2 FILLER_49_488 ();
 sg13g2_decap_4 FILLER_49_503 ();
 sg13g2_fill_1 FILLER_49_507 ();
 sg13g2_decap_8 FILLER_49_512 ();
 sg13g2_fill_2 FILLER_49_519 ();
 sg13g2_decap_8 FILLER_49_530 ();
 sg13g2_fill_2 FILLER_49_537 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_decap_8 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_8 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_8 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_decap_8 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_882 ();
 sg13g2_decap_8 FILLER_49_889 ();
 sg13g2_decap_8 FILLER_49_896 ();
 sg13g2_decap_8 FILLER_49_903 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_917 ();
 sg13g2_decap_8 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_8 FILLER_49_959 ();
 sg13g2_decap_8 FILLER_49_966 ();
 sg13g2_decap_8 FILLER_49_973 ();
 sg13g2_decap_8 FILLER_49_980 ();
 sg13g2_decap_8 FILLER_49_987 ();
 sg13g2_decap_8 FILLER_49_994 ();
 sg13g2_decap_8 FILLER_49_1001 ();
 sg13g2_decap_8 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1015 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 assign uio_oe[0] = net11;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net368;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net369;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
endmodule
