module heichips25_top_sorter (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire \s0.data_new_delayed[0] ;
 wire \s0.data_new_delayed[1] ;
 wire \s0.data_new_delayed[2] ;
 wire \s0.data_new_delayed[3] ;
 wire \s0.data_new_delayed[4] ;
 wire \s0.data_new_delayed[5] ;
 wire \s0.data_new_delayed[6] ;
 wire \s0.data_new_delayed[7] ;
 wire \s0.data_out[0][0] ;
 wire \s0.data_out[0][1] ;
 wire \s0.data_out[0][2] ;
 wire \s0.data_out[0][3] ;
 wire \s0.data_out[0][4] ;
 wire \s0.data_out[0][5] ;
 wire \s0.data_out[0][6] ;
 wire \s0.data_out[0][7] ;
 wire \s0.data_out[10][0] ;
 wire \s0.data_out[10][1] ;
 wire \s0.data_out[10][2] ;
 wire \s0.data_out[10][3] ;
 wire \s0.data_out[10][4] ;
 wire \s0.data_out[10][5] ;
 wire \s0.data_out[10][6] ;
 wire \s0.data_out[10][7] ;
 wire \s0.data_out[11][0] ;
 wire \s0.data_out[11][1] ;
 wire \s0.data_out[11][2] ;
 wire \s0.data_out[11][3] ;
 wire \s0.data_out[11][4] ;
 wire \s0.data_out[11][5] ;
 wire \s0.data_out[11][6] ;
 wire \s0.data_out[11][7] ;
 wire \s0.data_out[12][0] ;
 wire \s0.data_out[12][1] ;
 wire \s0.data_out[12][2] ;
 wire \s0.data_out[12][3] ;
 wire \s0.data_out[12][4] ;
 wire \s0.data_out[12][5] ;
 wire \s0.data_out[12][6] ;
 wire \s0.data_out[12][7] ;
 wire \s0.data_out[13][0] ;
 wire \s0.data_out[13][1] ;
 wire \s0.data_out[13][2] ;
 wire \s0.data_out[13][3] ;
 wire \s0.data_out[13][4] ;
 wire \s0.data_out[13][5] ;
 wire \s0.data_out[13][6] ;
 wire \s0.data_out[13][7] ;
 wire \s0.data_out[14][0] ;
 wire \s0.data_out[14][1] ;
 wire \s0.data_out[14][2] ;
 wire \s0.data_out[14][3] ;
 wire \s0.data_out[14][4] ;
 wire \s0.data_out[14][5] ;
 wire \s0.data_out[14][6] ;
 wire \s0.data_out[14][7] ;
 wire \s0.data_out[15][0] ;
 wire \s0.data_out[15][1] ;
 wire \s0.data_out[15][2] ;
 wire \s0.data_out[15][3] ;
 wire \s0.data_out[15][4] ;
 wire \s0.data_out[15][5] ;
 wire \s0.data_out[15][6] ;
 wire \s0.data_out[15][7] ;
 wire \s0.data_out[16][0] ;
 wire \s0.data_out[16][1] ;
 wire \s0.data_out[16][2] ;
 wire \s0.data_out[16][3] ;
 wire \s0.data_out[16][4] ;
 wire \s0.data_out[16][5] ;
 wire \s0.data_out[16][6] ;
 wire \s0.data_out[16][7] ;
 wire \s0.data_out[17][0] ;
 wire \s0.data_out[17][1] ;
 wire \s0.data_out[17][2] ;
 wire \s0.data_out[17][3] ;
 wire \s0.data_out[17][4] ;
 wire \s0.data_out[17][5] ;
 wire \s0.data_out[17][6] ;
 wire \s0.data_out[17][7] ;
 wire \s0.data_out[18][0] ;
 wire \s0.data_out[18][1] ;
 wire \s0.data_out[18][2] ;
 wire \s0.data_out[18][3] ;
 wire \s0.data_out[18][4] ;
 wire \s0.data_out[18][5] ;
 wire \s0.data_out[18][6] ;
 wire \s0.data_out[18][7] ;
 wire \s0.data_out[19][0] ;
 wire \s0.data_out[19][1] ;
 wire \s0.data_out[19][2] ;
 wire \s0.data_out[19][3] ;
 wire \s0.data_out[19][4] ;
 wire \s0.data_out[19][5] ;
 wire \s0.data_out[19][6] ;
 wire \s0.data_out[19][7] ;
 wire \s0.data_out[1][0] ;
 wire \s0.data_out[1][1] ;
 wire \s0.data_out[1][2] ;
 wire \s0.data_out[1][3] ;
 wire \s0.data_out[1][4] ;
 wire \s0.data_out[1][5] ;
 wire \s0.data_out[1][6] ;
 wire \s0.data_out[1][7] ;
 wire \s0.data_out[20][0] ;
 wire \s0.data_out[20][1] ;
 wire \s0.data_out[20][2] ;
 wire \s0.data_out[20][3] ;
 wire \s0.data_out[20][4] ;
 wire \s0.data_out[20][5] ;
 wire \s0.data_out[20][6] ;
 wire \s0.data_out[20][7] ;
 wire \s0.data_out[21][0] ;
 wire \s0.data_out[21][1] ;
 wire \s0.data_out[21][2] ;
 wire \s0.data_out[21][3] ;
 wire \s0.data_out[21][4] ;
 wire \s0.data_out[21][5] ;
 wire \s0.data_out[21][6] ;
 wire \s0.data_out[21][7] ;
 wire \s0.data_out[22][0] ;
 wire \s0.data_out[22][1] ;
 wire \s0.data_out[22][2] ;
 wire \s0.data_out[22][3] ;
 wire \s0.data_out[22][4] ;
 wire \s0.data_out[22][5] ;
 wire \s0.data_out[22][6] ;
 wire \s0.data_out[22][7] ;
 wire \s0.data_out[23][0] ;
 wire \s0.data_out[23][1] ;
 wire \s0.data_out[23][2] ;
 wire \s0.data_out[23][3] ;
 wire \s0.data_out[23][4] ;
 wire \s0.data_out[23][5] ;
 wire \s0.data_out[23][6] ;
 wire \s0.data_out[23][7] ;
 wire \s0.data_out[2][0] ;
 wire \s0.data_out[2][1] ;
 wire \s0.data_out[2][2] ;
 wire \s0.data_out[2][3] ;
 wire \s0.data_out[2][4] ;
 wire \s0.data_out[2][5] ;
 wire \s0.data_out[2][6] ;
 wire \s0.data_out[2][7] ;
 wire \s0.data_out[3][0] ;
 wire \s0.data_out[3][1] ;
 wire \s0.data_out[3][2] ;
 wire \s0.data_out[3][3] ;
 wire \s0.data_out[3][4] ;
 wire \s0.data_out[3][5] ;
 wire \s0.data_out[3][6] ;
 wire \s0.data_out[3][7] ;
 wire \s0.data_out[4][0] ;
 wire \s0.data_out[4][1] ;
 wire \s0.data_out[4][2] ;
 wire \s0.data_out[4][3] ;
 wire \s0.data_out[4][4] ;
 wire \s0.data_out[4][5] ;
 wire \s0.data_out[4][6] ;
 wire \s0.data_out[4][7] ;
 wire \s0.data_out[5][0] ;
 wire \s0.data_out[5][1] ;
 wire \s0.data_out[5][2] ;
 wire \s0.data_out[5][3] ;
 wire \s0.data_out[5][4] ;
 wire \s0.data_out[5][5] ;
 wire \s0.data_out[5][6] ;
 wire \s0.data_out[5][7] ;
 wire \s0.data_out[6][0] ;
 wire \s0.data_out[6][1] ;
 wire \s0.data_out[6][2] ;
 wire \s0.data_out[6][3] ;
 wire \s0.data_out[6][4] ;
 wire \s0.data_out[6][5] ;
 wire \s0.data_out[6][6] ;
 wire \s0.data_out[6][7] ;
 wire \s0.data_out[7][0] ;
 wire \s0.data_out[7][1] ;
 wire \s0.data_out[7][2] ;
 wire \s0.data_out[7][3] ;
 wire \s0.data_out[7][4] ;
 wire \s0.data_out[7][5] ;
 wire \s0.data_out[7][6] ;
 wire \s0.data_out[7][7] ;
 wire \s0.data_out[8][0] ;
 wire \s0.data_out[8][1] ;
 wire \s0.data_out[8][2] ;
 wire \s0.data_out[8][3] ;
 wire \s0.data_out[8][4] ;
 wire \s0.data_out[8][5] ;
 wire \s0.data_out[8][6] ;
 wire \s0.data_out[8][7] ;
 wire \s0.data_out[9][0] ;
 wire \s0.data_out[9][1] ;
 wire \s0.data_out[9][2] ;
 wire \s0.data_out[9][3] ;
 wire \s0.data_out[9][4] ;
 wire \s0.data_out[9][5] ;
 wire \s0.data_out[9][6] ;
 wire \s0.data_out[9][7] ;
 wire \s0.genblk1[10].modules.bubble ;
 wire \s0.genblk1[11].modules.bubble ;
 wire \s0.genblk1[12].modules.bubble ;
 wire \s0.genblk1[13].modules.bubble ;
 wire \s0.genblk1[14].modules.bubble ;
 wire \s0.genblk1[15].modules.bubble ;
 wire \s0.genblk1[16].modules.bubble ;
 wire \s0.genblk1[17].modules.bubble ;
 wire \s0.genblk1[18].modules.bubble ;
 wire \s0.genblk1[19].modules.bubble ;
 wire \s0.genblk1[1].modules.bubble ;
 wire \s0.genblk1[20].modules.bubble ;
 wire \s0.genblk1[21].modules.bubble ;
 wire \s0.genblk1[22].modules.bubble ;
 wire \s0.genblk1[23].modules.bubble ;
 wire \s0.genblk1[2].modules.bubble ;
 wire \s0.genblk1[3].modules.bubble ;
 wire \s0.genblk1[4].modules.bubble ;
 wire \s0.genblk1[5].modules.bubble ;
 wire \s0.genblk1[6].modules.bubble ;
 wire \s0.genblk1[7].modules.bubble ;
 wire \s0.genblk1[8].modules.bubble ;
 wire \s0.genblk1[9].modules.bubble ;
 wire \s0.module0.bubble ;
 wire net11;
 wire net12;
 wire net320;
 wire net13;
 wire net14;
 wire clknet_leaf_0_clk;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net1;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net10;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire [0:0] \s0.shift_out[0] ;
 wire [0:0] \s0.shift_out[10] ;
 wire [0:0] \s0.shift_out[11] ;
 wire [0:0] \s0.shift_out[12] ;
 wire [0:0] \s0.shift_out[13] ;
 wire [0:0] \s0.shift_out[14] ;
 wire [0:0] \s0.shift_out[15] ;
 wire [0:0] \s0.shift_out[16] ;
 wire [0:0] \s0.shift_out[17] ;
 wire [0:0] \s0.shift_out[18] ;
 wire [0:0] \s0.shift_out[19] ;
 wire [0:0] \s0.shift_out[1] ;
 wire [0:0] \s0.shift_out[20] ;
 wire [0:0] \s0.shift_out[21] ;
 wire [0:0] \s0.shift_out[22] ;
 wire [0:0] \s0.shift_out[23] ;
 wire [0:0] \s0.shift_out[2] ;
 wire [0:0] \s0.shift_out[3] ;
 wire [0:0] \s0.shift_out[4] ;
 wire [0:0] \s0.shift_out[5] ;
 wire [0:0] \s0.shift_out[6] ;
 wire [0:0] \s0.shift_out[7] ;
 wire [0:0] \s0.shift_out[8] ;
 wire [0:0] \s0.shift_out[9] ;
 wire [0:0] \s0.valid_out[0] ;
 wire [0:0] \s0.valid_out[10] ;
 wire [0:0] \s0.valid_out[11] ;
 wire [0:0] \s0.valid_out[12] ;
 wire [0:0] \s0.valid_out[13] ;
 wire [0:0] \s0.valid_out[14] ;
 wire [0:0] \s0.valid_out[15] ;
 wire [0:0] \s0.valid_out[16] ;
 wire [0:0] \s0.valid_out[17] ;
 wire [0:0] \s0.valid_out[18] ;
 wire [0:0] \s0.valid_out[19] ;
 wire [0:0] \s0.valid_out[1] ;
 wire [0:0] \s0.valid_out[20] ;
 wire [0:0] \s0.valid_out[21] ;
 wire [0:0] \s0.valid_out[22] ;
 wire [0:0] \s0.valid_out[23] ;
 wire [0:0] \s0.valid_out[2] ;
 wire [0:0] \s0.valid_out[3] ;
 wire [0:0] \s0.valid_out[4] ;
 wire [0:0] \s0.valid_out[5] ;
 wire [0:0] \s0.valid_out[6] ;
 wire [0:0] \s0.valid_out[7] ;
 wire [0:0] \s0.valid_out[8] ;
 wire [0:0] \s0.valid_out[9] ;
 wire [0:0] \s0.was_valid_out[0] ;
 wire [0:0] \s0.was_valid_out[10] ;
 wire [0:0] \s0.was_valid_out[11] ;
 wire [0:0] \s0.was_valid_out[12] ;
 wire [0:0] \s0.was_valid_out[13] ;
 wire [0:0] \s0.was_valid_out[14] ;
 wire [0:0] \s0.was_valid_out[15] ;
 wire [0:0] \s0.was_valid_out[16] ;
 wire [0:0] \s0.was_valid_out[17] ;
 wire [0:0] \s0.was_valid_out[18] ;
 wire [0:0] \s0.was_valid_out[19] ;
 wire [0:0] \s0.was_valid_out[1] ;
 wire [0:0] \s0.was_valid_out[20] ;
 wire [0:0] \s0.was_valid_out[21] ;
 wire [0:0] \s0.was_valid_out[22] ;
 wire [0:0] \s0.was_valid_out[23] ;
 wire [0:0] \s0.was_valid_out[2] ;
 wire [0:0] \s0.was_valid_out[3] ;
 wire [0:0] \s0.was_valid_out[4] ;
 wire [0:0] \s0.was_valid_out[5] ;
 wire [0:0] \s0.was_valid_out[6] ;
 wire [0:0] \s0.was_valid_out[7] ;
 wire [0:0] \s0.was_valid_out[8] ;
 wire [0:0] \s0.was_valid_out[9] ;

 sg13g2_and2_1 _3389_ (.A(net328),
    .B(net1485),
    .X(_0099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3390_ (.Y(_1004_),
    .A(net1220),
    .B(net548),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3391_ (.A0(\s0.data_out[15][2] ),
    .A1(\s0.data_out[14][2] ),
    .S(net1219),
    .X(_1005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3392_ (.A(net1213),
    .B_N(net1164),
    .Y(_1006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3393_ (.A2(_1005_),
    .A1(net1215),
    .B1(_1006_),
    .X(_1007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3394_ (.Y(_1008_),
    .B(\s0.data_out[14][2] ),
    .A_N(net1232),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3395_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0893_),
    .A2(_1008_),
    .Y(_1009_),
    .B1(net1227));
 sg13g2_a21oi_1 _3396_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1227),
    .A2(_1007_),
    .Y(_1010_),
    .B1(_1009_));
 sg13g2_or2_1 _3397_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1011_),
    .B(_1010_),
    .A(net1445));
 sg13g2_nor2b_1 _3398_ (.A(net1213),
    .B_N(net1168),
    .Y(_1012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3399_ (.Y(_1013_),
    .A(net1219),
    .B(net647),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3400_ (.B1(_1013_),
    .VDD(VPWR),
    .Y(_1014_),
    .VSS(VGND),
    .A1(net1220),
    .A2(_2818_));
 sg13g2_a21o_1 _3401_ (.A2(_1014_),
    .A1(net1213),
    .B1(_1012_),
    .X(_1015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3402_ (.Y(_1016_),
    .B(\s0.data_out[14][1] ),
    .A_N(net1235),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3403_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0901_),
    .A2(_1016_),
    .Y(_1017_),
    .B1(net1225));
 sg13g2_a21oi_1 _3404_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1227),
    .A2(_1015_),
    .Y(_1018_),
    .B1(_1017_));
 sg13g2_mux2_1 _3405_ (.A0(\s0.data_out[15][0] ),
    .A1(\s0.data_out[14][0] ),
    .S(net1219),
    .X(_1019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3406_ (.A(net1213),
    .B_N(net1171),
    .Y(_1020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3407_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1213),
    .A2(_1019_),
    .Y(_1021_),
    .B1(_1020_));
 sg13g2_nand2b_1 _3408_ (.Y(_1022_),
    .B(net1228),
    .A_N(_1021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3409_ (.A0(\s0.data_out[14][0] ),
    .A1(\s0.data_out[15][0] ),
    .S(net1232),
    .X(_1023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3410_ (.Y(_1024_),
    .B(_1023_),
    .A_N(net1228),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3411_ (.B1(_1011_),
    .VDD(VPWR),
    .Y(_1025_),
    .VSS(VGND),
    .A1(net1454),
    .A2(_1018_));
 sg13g2_a221oi_1 _3412_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1024_),
    .C1(net1460),
    .B1(_1022_),
    .A1(net1454),
    .Y(_1026_),
    .A2(_1018_));
 sg13g2_nand2_1 _3413_ (.Y(_1027_),
    .A(net1219),
    .B(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3414_ (.B1(_1027_),
    .VDD(VPWR),
    .Y(_1028_),
    .VSS(VGND),
    .A1(net1219),
    .A2(_2816_));
 sg13g2_nor2_1 _3415_ (.A(net1213),
    .B(net993),
    .Y(_1029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3416_ (.A2(_1028_),
    .A1(net1213),
    .B1(_1029_),
    .X(_1030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3417_ (.Y(_1031_),
    .B(\s0.data_out[14][3] ),
    .A_N(net1235),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3418_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0916_),
    .A2(_1031_),
    .Y(_1032_),
    .B1(net1227));
 sg13g2_a21oi_1 _3419_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1227),
    .A2(_1030_),
    .Y(_1033_),
    .B1(_1032_));
 sg13g2_a22oi_1 _3420_ (.Y(_1034_),
    .B1(_1033_),
    .B2(net1440),
    .A2(_1010_),
    .A1(net1445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3421_ (.B1(_1034_),
    .VDD(VPWR),
    .Y(_1035_),
    .VSS(VGND),
    .A1(_1025_),
    .A2(_1026_));
 sg13g2_nand2_1 _3422_ (.Y(_1036_),
    .A(net1222),
    .B(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3423_ (.A0(\s0.data_out[15][7] ),
    .A1(\s0.data_out[14][7] ),
    .S(net1221),
    .X(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3424_ (.A(net1217),
    .B_N(net1145),
    .Y(_1038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3425_ (.A2(_1037_),
    .A1(net1217),
    .B1(_1038_),
    .X(_1039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3426_ (.Y(_1040_),
    .B(\s0.data_out[14][7] ),
    .A_N(net1234),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3427_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0932_),
    .A2(_1040_),
    .Y(_1041_),
    .B1(net1229));
 sg13g2_a21oi_1 _3428_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1229),
    .A2(_1039_),
    .Y(_1042_),
    .B1(_1041_));
 sg13g2_nand2_1 _3429_ (.Y(_1043_),
    .A(net1221),
    .B(net545),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3430_ (.A0(\s0.data_out[15][6] ),
    .A1(\s0.data_out[14][6] ),
    .S(net1221),
    .X(_1044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3431_ (.A(net1217),
    .B_N(net1150),
    .Y(_1045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3432_ (.A2(_1044_),
    .A1(net1217),
    .B1(_1045_),
    .X(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3433_ (.Y(_1047_),
    .B(net545),
    .A_N(net1234),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3434_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0925_),
    .A2(_1047_),
    .Y(_1048_),
    .B1(net1230));
 sg13g2_a21oi_1 _3435_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1229),
    .A2(_1046_),
    .Y(_1049_),
    .B1(_1048_));
 sg13g2_a22oi_1 _3436_ (.Y(_1050_),
    .B1(_1049_),
    .B2(net1413),
    .A2(_1042_),
    .A1(net1404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3437_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1051_),
    .B(_1049_),
    .A(net1413));
 sg13g2_or2_1 _3438_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1052_),
    .B(_1042_),
    .A(net1404));
 sg13g2_inv_1 _3439_ (.VDD(VPWR),
    .Y(_1053_),
    .A(_1052_),
    .VSS(VGND));
 sg13g2_and3_1 _3440_ (.X(_1054_),
    .A(_1050_),
    .B(_1051_),
    .C(_1052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3441_ (.B(_1051_),
    .C(_1052_),
    .A(_1050_),
    .Y(_1055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3442_ (.A0(\s0.data_out[15][5] ),
    .A1(\s0.data_out[14][5] ),
    .S(net1219),
    .X(_1056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3443_ (.A(net1215),
    .B_N(net1154),
    .Y(_1057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3444_ (.A2(_1056_),
    .A1(net1215),
    .B1(_1057_),
    .X(_1058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3445_ (.Y(_1059_),
    .B(\s0.data_out[14][5] ),
    .A_N(net1234),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3446_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0953_),
    .A2(_1059_),
    .Y(_1060_),
    .B1(net1230));
 sg13g2_a21oi_1 _3447_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1230),
    .A2(_1058_),
    .Y(_1061_),
    .B1(_1060_));
 sg13g2_nor2_1 _3448_ (.A(net1423),
    .B(_1061_),
    .Y(_1062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3449_ (.Y(_1063_),
    .A(net1221),
    .B(\s0.data_out[14][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3450_ (.A0(\s0.data_out[15][4] ),
    .A1(\s0.data_out[14][4] ),
    .S(net1220),
    .X(_1064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3451_ (.A(net1216),
    .B_N(net1159),
    .Y(_1065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3452_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1216),
    .A2(_1064_),
    .Y(_1066_),
    .B1(_1065_));
 sg13g2_nand2b_1 _3453_ (.Y(_1067_),
    .B(net1230),
    .A_N(_1066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3454_ (.B1(_0945_),
    .VDD(VPWR),
    .Y(_1068_),
    .VSS(VGND),
    .A1(net1234),
    .A2(_2821_));
 sg13g2_nand2b_1 _3455_ (.Y(_1069_),
    .B(_1068_),
    .A_N(net1230),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3456_ (.B(_1067_),
    .C(_1069_),
    .A(net1432),
    .Y(_1070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3457_ (.Y(_1071_),
    .A(net1423),
    .B(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3458_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1067_),
    .A2(_1069_),
    .Y(_1072_),
    .B1(net1432));
 sg13g2_o21ai_1 _3459_ (.B1(_1071_),
    .VDD(VPWR),
    .Y(_1073_),
    .VSS(VGND),
    .A1(net1440),
    .A2(_1033_));
 sg13g2_nand2b_1 _3460_ (.Y(_1074_),
    .B(_1070_),
    .A_N(_1062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3461_ (.A(_1055_),
    .B(_1072_),
    .C(_1073_),
    .D(_1074_),
    .Y(_1075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3462_ (.B1(_1071_),
    .VDD(VPWR),
    .Y(_1076_),
    .VSS(VGND),
    .A1(_1062_),
    .A2(_1070_));
 sg13g2_o21ai_1 _3463_ (.B1(_0998_),
    .VDD(VPWR),
    .Y(_1077_),
    .VSS(VGND),
    .A1(_1050_),
    .A2(_1053_));
 sg13g2_a221oi_1 _3464_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1054_),
    .C1(_1077_),
    .B1(_1076_),
    .A1(_1035_),
    .Y(_1078_),
    .A2(_1075_));
 sg13g2_nor3_1 _3465_ (.A(net323),
    .B(net1332),
    .C(_1078_),
    .Y(_0100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3466_ (.A(net1213),
    .B(\s0.data_out[14][0] ),
    .X(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3467_ (.B1(net1228),
    .VDD(VPWR),
    .Y(_1080_),
    .VSS(VGND),
    .A1(_1020_),
    .A2(_1079_));
 sg13g2_nand3_1 _3468_ (.B(_1024_),
    .C(_1080_),
    .A(net1477),
    .Y(_1081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3469_ (.B1(_1081_),
    .VDD(VPWR),
    .Y(_1082_),
    .VSS(VGND),
    .A1(net1477),
    .A2(net607));
 sg13g2_inv_1 _3470_ (.VDD(VPWR),
    .Y(_0101_),
    .A(_1082_),
    .VSS(VGND));
 sg13g2_nor2_1 _3471_ (.A(net1018),
    .B(_2824_),
    .Y(_1083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3472_ (.B1(net1227),
    .VDD(VPWR),
    .Y(_1084_),
    .VSS(VGND),
    .A1(_1012_),
    .A2(_1083_));
 sg13g2_nor2_1 _3473_ (.A(net1369),
    .B(_1017_),
    .Y(_1085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3474_ (.Y(_0102_),
    .B1(_1084_),
    .B2(_1085_),
    .A2(_2818_),
    .A1(net1369),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3475_ (.A(net1018),
    .B(_2823_),
    .Y(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3476_ (.B1(net1227),
    .VDD(VPWR),
    .Y(_1087_),
    .VSS(VGND),
    .A1(_1006_),
    .A2(_1086_));
 sg13g2_nor2_1 _3477_ (.A(net1367),
    .B(_1009_),
    .Y(_1088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3478_ (.Y(_0103_),
    .B1(_1087_),
    .B2(_1088_),
    .A2(_2817_),
    .A1(net1368),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3479_ (.A(net1018),
    .B(_2822_),
    .Y(_1089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3480_ (.B1(net1227),
    .VDD(VPWR),
    .Y(_1090_),
    .VSS(VGND),
    .A1(_1029_),
    .A2(_1089_));
 sg13g2_nor2_1 _3481_ (.A(net1367),
    .B(_1032_),
    .Y(_1091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3482_ (.Y(_0104_),
    .B1(_1090_),
    .B2(_1091_),
    .A2(_2816_),
    .A1(net1367),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3483_ (.A(net1018),
    .B(_2821_),
    .Y(_1092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3484_ (.B1(net1230),
    .VDD(VPWR),
    .Y(_1093_),
    .VSS(VGND),
    .A1(_1065_),
    .A2(_1092_));
 sg13g2_nand3_1 _3485_ (.B(_1069_),
    .C(_1093_),
    .A(net1484),
    .Y(_1094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3486_ (.B1(_1094_),
    .VDD(VPWR),
    .Y(_1095_),
    .VSS(VGND),
    .A1(net1484),
    .A2(net643));
 sg13g2_inv_1 _3487_ (.VDD(VPWR),
    .Y(_0105_),
    .A(_1095_),
    .VSS(VGND));
 sg13g2_and2_1 _3488_ (.A(net1215),
    .B(\s0.data_out[14][5] ),
    .X(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3489_ (.B1(net1230),
    .VDD(VPWR),
    .Y(_1097_),
    .VSS(VGND),
    .A1(_1057_),
    .A2(_1096_));
 sg13g2_nor2_1 _3490_ (.A(net1380),
    .B(_1060_),
    .Y(_1098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3491_ (.Y(_0106_),
    .B1(_1097_),
    .B2(_1098_),
    .A2(_2815_),
    .A1(net1380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3492_ (.A(net1017),
    .B(_2820_),
    .Y(_1099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3493_ (.B1(net1229),
    .VDD(VPWR),
    .Y(_1100_),
    .VSS(VGND),
    .A1(_1045_),
    .A2(_1099_));
 sg13g2_nand3b_1 _3494_ (.B(_1100_),
    .C(net1485),
    .Y(_1101_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1048_));
 sg13g2_o21ai_1 _3495_ (.B1(_1101_),
    .VDD(VPWR),
    .Y(_1102_),
    .VSS(VGND),
    .A1(net1485),
    .A2(net693));
 sg13g2_inv_1 _3496_ (.VDD(VPWR),
    .Y(_0107_),
    .A(net694),
    .VSS(VGND));
 sg13g2_nor2_1 _3497_ (.A(net1017),
    .B(_2819_),
    .Y(_1103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3498_ (.B1(net1229),
    .VDD(VPWR),
    .Y(_1104_),
    .VSS(VGND),
    .A1(_1038_),
    .A2(_1103_));
 sg13g2_nor2_1 _3499_ (.A(net1380),
    .B(_1041_),
    .Y(_1105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3500_ (.Y(_0108_),
    .B1(_1104_),
    .B2(_1105_),
    .A2(_2814_),
    .A1(net1380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3501_ (.B1(net1218),
    .VDD(VPWR),
    .Y(_1106_),
    .VSS(VGND),
    .A1(net1205),
    .A2(net1395));
 sg13g2_nor2_1 _3502_ (.A(_2740_),
    .B(net1395),
    .Y(_1107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3503_ (.A(_1106_),
    .B(_1107_),
    .Y(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3504_ (.VDD(VPWR),
    .Y(_1109_),
    .A(_1108_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3505_ (.B1(_1109_),
    .VDD(VPWR),
    .Y(_1110_),
    .VSS(VGND),
    .A1(net1217),
    .A2(_0995_));
 sg13g2_or2_1 _3506_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1111_),
    .B(net1211),
    .A(net566));
 sg13g2_o21ai_1 _3507_ (.B1(net1018),
    .VDD(VPWR),
    .Y(_1112_),
    .VSS(VGND),
    .A1(net566),
    .A2(net1222));
 sg13g2_o21ai_1 _3508_ (.B1(_1112_),
    .VDD(VPWR),
    .Y(_1113_),
    .VSS(VGND),
    .A1(net1205),
    .A2(_1106_));
 sg13g2_a21oi_1 _3509_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1108_),
    .A2(_1111_),
    .Y(_1114_),
    .B1(_1113_));
 sg13g2_o21ai_1 _3510_ (.B1(net1485),
    .VDD(VPWR),
    .Y(_1115_),
    .VSS(VGND),
    .A1(net615),
    .A2(_1110_));
 sg13g2_nor2_1 _3511_ (.A(_1114_),
    .B(_1115_),
    .Y(_0109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3512_ (.A(net1381),
    .B(_1110_),
    .Y(_0110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3513_ (.A(net1485),
    .B(net343),
    .X(_0111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3514_ (.Y(_1116_),
    .A(net1212),
    .B(net457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3515_ (.A0(\s0.data_out[14][2] ),
    .A1(\s0.data_out[13][2] ),
    .S(net1210),
    .X(_1117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3516_ (.A(net1203),
    .B_N(net1164),
    .Y(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3517_ (.A2(_1117_),
    .A1(net1203),
    .B1(_1118_),
    .X(_1119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3518_ (.Y(_1120_),
    .B(net457),
    .A_N(net1220),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3519_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1004_),
    .A2(_1120_),
    .Y(_1121_),
    .B1(net1216));
 sg13g2_a21oi_1 _3520_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1216),
    .A2(_1119_),
    .Y(_1122_),
    .B1(_1121_));
 sg13g2_or2_1 _3521_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1123_),
    .B(_1122_),
    .A(net1445));
 sg13g2_nand2_1 _3522_ (.Y(_1124_),
    .A(net1210),
    .B(net481),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3523_ (.B1(_1124_),
    .VDD(VPWR),
    .Y(_1125_),
    .VSS(VGND),
    .A1(net1210),
    .A2(_2824_));
 sg13g2_nor2b_1 _3524_ (.A(net1201),
    .B_N(net1169),
    .Y(_1126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3525_ (.A2(_1125_),
    .A1(net1201),
    .B1(_1126_),
    .X(_1127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3526_ (.Y(_1128_),
    .B(net481),
    .A_N(net1219),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3527_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1013_),
    .A2(_1128_),
    .Y(_1129_),
    .B1(net1214));
 sg13g2_a21oi_1 _3528_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1214),
    .A2(_1127_),
    .Y(_1130_),
    .B1(_1129_));
 sg13g2_mux2_1 _3529_ (.A0(\s0.data_out[14][0] ),
    .A1(\s0.data_out[13][0] ),
    .S(net1210),
    .X(_1131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3530_ (.A(net1201),
    .B_N(net1172),
    .Y(_1132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3531_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1201),
    .A2(_1131_),
    .Y(_1133_),
    .B1(_1132_));
 sg13g2_nand2b_1 _3532_ (.Y(_1134_),
    .B(net1214),
    .A_N(_1133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3533_ (.A0(\s0.data_out[13][0] ),
    .A1(\s0.data_out[14][0] ),
    .S(net1219),
    .X(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3534_ (.Y(_1136_),
    .A(net1018),
    .B(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3535_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1136_),
    .C1(net1459),
    .B1(_1134_),
    .A1(net1454),
    .Y(_1137_),
    .A2(_1130_));
 sg13g2_o21ai_1 _3536_ (.B1(_1123_),
    .VDD(VPWR),
    .Y(_1138_),
    .VSS(VGND),
    .A1(net1454),
    .A2(_1130_));
 sg13g2_nand2_1 _3537_ (.Y(_1139_),
    .A(net1210),
    .B(net532),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3538_ (.B1(_1139_),
    .VDD(VPWR),
    .Y(_1140_),
    .VSS(VGND),
    .A1(net1210),
    .A2(_2822_));
 sg13g2_nor2_1 _3539_ (.A(net1203),
    .B(net994),
    .Y(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3540_ (.A2(_1140_),
    .A1(net1203),
    .B1(_1141_),
    .X(_1142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3541_ (.Y(_1143_),
    .B(net532),
    .A_N(net1220),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3542_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1027_),
    .A2(_1143_),
    .Y(_1144_),
    .B1(net1214));
 sg13g2_a21oi_1 _3543_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1216),
    .A2(_1142_),
    .Y(_1145_),
    .B1(_1144_));
 sg13g2_a22oi_1 _3544_ (.Y(_1146_),
    .B1(_1145_),
    .B2(net1441),
    .A2(_1122_),
    .A1(net1445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3545_ (.B1(_1146_),
    .VDD(VPWR),
    .Y(_1147_),
    .VSS(VGND),
    .A1(_1137_),
    .A2(_1138_));
 sg13g2_nand2_1 _3546_ (.Y(_1148_),
    .A(net1211),
    .B(net406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3547_ (.B1(_1148_),
    .VDD(VPWR),
    .Y(_1149_),
    .VSS(VGND),
    .A1(net1211),
    .A2(_2819_));
 sg13g2_nor2b_1 _3548_ (.A(net1206),
    .B_N(net1145),
    .Y(_1150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3549_ (.A2(_1149_),
    .A1(net1206),
    .B1(_1150_),
    .X(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3550_ (.Y(_1152_),
    .B(net406),
    .A_N(net1222),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3551_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1036_),
    .A2(_1152_),
    .Y(_1153_),
    .B1(net1218));
 sg13g2_a21oi_1 _3552_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1218),
    .A2(_1151_),
    .Y(_1154_),
    .B1(_1153_));
 sg13g2_nand2_1 _3553_ (.Y(_1155_),
    .A(net1211),
    .B(\s0.data_out[13][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3554_ (.B1(_1155_),
    .VDD(VPWR),
    .Y(_1156_),
    .VSS(VGND),
    .A1(net1211),
    .A2(_2820_));
 sg13g2_nor2b_1 _3555_ (.A(net1206),
    .B_N(net1150),
    .Y(_1157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3556_ (.A2(_1156_),
    .A1(net1206),
    .B1(_1157_),
    .X(_1158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3557_ (.Y(_1159_),
    .B(\s0.data_out[13][6] ),
    .A_N(net1222),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3558_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1043_),
    .A2(_1159_),
    .Y(_1160_),
    .B1(net1218));
 sg13g2_a21oi_1 _3559_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\s0.shift_out[14] [0]),
    .A2(_1158_),
    .Y(_1161_),
    .B1(_1160_));
 sg13g2_a22oi_1 _3560_ (.Y(_1162_),
    .B1(_1161_),
    .B2(net1413),
    .A2(_1154_),
    .A1(net1404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3561_ (.VDD(VPWR),
    .Y(_1163_),
    .A(_1162_),
    .VSS(VGND));
 sg13g2_or2_1 _3562_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1164_),
    .B(_1161_),
    .A(net1413));
 sg13g2_or2_1 _3563_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1165_),
    .B(_1154_),
    .A(net1404));
 sg13g2_and3_1 _3564_ (.X(_1166_),
    .A(_1162_),
    .B(_1164_),
    .C(_1165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3565_ (.A0(\s0.data_out[14][5] ),
    .A1(\s0.data_out[13][5] ),
    .S(net1211),
    .X(_1167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3566_ (.A(net1205),
    .B_N(net1154),
    .Y(_1168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3567_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1205),
    .A2(_1167_),
    .Y(_1169_),
    .B1(_1168_));
 sg13g2_nand2b_1 _3568_ (.Y(_1170_),
    .B(net1218),
    .A_N(_1169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3569_ (.A0(\s0.data_out[13][5] ),
    .A1(\s0.data_out[14][5] ),
    .S(net1221),
    .X(_1171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3570_ (.Y(_1172_),
    .A(_2741_),
    .B(_1171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3571_ (.B(_1170_),
    .C(_1172_),
    .A(net1423),
    .Y(_1173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3572_ (.B1(_1173_),
    .VDD(VPWR),
    .Y(_1174_),
    .VSS(VGND),
    .A1(net1441),
    .A2(_1145_));
 sg13g2_a21oi_1 _3573_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1170_),
    .A2(_1172_),
    .Y(_1175_),
    .B1(net1423));
 sg13g2_nor2b_1 _3574_ (.A(net1204),
    .B_N(net1159),
    .Y(_1176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3575_ (.Y(_1177_),
    .A(net1211),
    .B(\s0.data_out[13][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3576_ (.B1(_1177_),
    .VDD(VPWR),
    .Y(_1178_),
    .VSS(VGND),
    .A1(net1210),
    .A2(_2821_));
 sg13g2_a21oi_1 _3577_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1204),
    .A2(_1178_),
    .Y(_1179_),
    .B1(_1176_));
 sg13g2_o21ai_1 _3578_ (.B1(_1063_),
    .VDD(VPWR),
    .Y(_1180_),
    .VSS(VGND),
    .A1(net1221),
    .A2(_2826_));
 sg13g2_nand2_1 _3579_ (.Y(_1181_),
    .A(net1017),
    .B(_1180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3580_ (.B1(_1181_),
    .VDD(VPWR),
    .Y(_1182_),
    .VSS(VGND),
    .A1(net1017),
    .A2(_1179_));
 sg13g2_or2_1 _3581_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1183_),
    .B(_1182_),
    .A(_2768_));
 sg13g2_xnor2_1 _3582_ (.Y(_1184_),
    .A(_2768_),
    .B(_1182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3583_ (.A(_1174_),
    .B(_1175_),
    .C(_1184_),
    .Y(_1185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3584_ (.B(_1166_),
    .C(_1185_),
    .A(_1147_),
    .Y(_1186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3585_ (.B1(_1173_),
    .VDD(VPWR),
    .Y(_1187_),
    .VSS(VGND),
    .A1(_1175_),
    .A2(_1183_));
 sg13g2_a221oi_1 _3586_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1187_),
    .C1(_1110_),
    .B1(_1166_),
    .A1(_1163_),
    .Y(_1188_),
    .A2(_1165_));
 sg13g2_or2_1 _3587_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1189_),
    .B(net1332),
    .A(net328));
 sg13g2_a21oi_1 _3588_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1186_),
    .A2(_1188_),
    .Y(_0112_),
    .B1(_1189_));
 sg13g2_a21oi_1 _3589_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1201),
    .A2(\s0.data_out[13][0] ),
    .Y(_1190_),
    .B1(_1132_));
 sg13g2_a21oi_1 _3590_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1018),
    .A2(_1135_),
    .Y(_1191_),
    .B1(net1378));
 sg13g2_o21ai_1 _3591_ (.B1(_1191_),
    .VDD(VPWR),
    .Y(_1192_),
    .VSS(VGND),
    .A1(net1018),
    .A2(_1190_));
 sg13g2_o21ai_1 _3592_ (.B1(_1192_),
    .VDD(VPWR),
    .Y(_1193_),
    .VSS(VGND),
    .A1(net1477),
    .A2(net591));
 sg13g2_inv_1 _3593_ (.VDD(VPWR),
    .Y(_0113_),
    .A(net592),
    .VSS(VGND));
 sg13g2_and2_1 _3594_ (.A(net1201),
    .B(net481),
    .X(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3595_ (.B1(net1214),
    .VDD(VPWR),
    .Y(_1195_),
    .VSS(VGND),
    .A1(_1126_),
    .A2(_1194_));
 sg13g2_nor2_1 _3596_ (.A(net1378),
    .B(_1129_),
    .Y(_1196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3597_ (.Y(_0114_),
    .B1(_1195_),
    .B2(_1196_),
    .A2(_2824_),
    .A1(net1378),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3598_ (.A(net1203),
    .B(net457),
    .X(_1197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3599_ (.B1(net1216),
    .VDD(VPWR),
    .Y(_1198_),
    .VSS(VGND),
    .A1(_1118_),
    .A2(_1197_));
 sg13g2_nor2_1 _3600_ (.A(net1380),
    .B(_1121_),
    .Y(_1199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3601_ (.Y(_0115_),
    .B1(_1198_),
    .B2(_1199_),
    .A2(_2823_),
    .A1(net1380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3602_ (.A(net1203),
    .B(net532),
    .X(_1200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3603_ (.B1(net1216),
    .VDD(VPWR),
    .Y(_1201_),
    .VSS(VGND),
    .A1(_1141_),
    .A2(_1200_));
 sg13g2_nor2_1 _3604_ (.A(net1378),
    .B(_1144_),
    .Y(_1202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3605_ (.Y(_0116_),
    .B1(_1201_),
    .B2(_1202_),
    .A2(_2822_),
    .A1(net1378),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3606_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1204),
    .A2(net491),
    .Y(_1203_),
    .B1(_1176_));
 sg13g2_a21oi_1 _3607_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1017),
    .A2(_1180_),
    .Y(_1204_),
    .B1(net1380));
 sg13g2_o21ai_1 _3608_ (.B1(_1204_),
    .VDD(VPWR),
    .Y(_1205_),
    .VSS(VGND),
    .A1(net1017),
    .A2(_1203_));
 sg13g2_o21ai_1 _3609_ (.B1(_1205_),
    .VDD(VPWR),
    .Y(_1206_),
    .VSS(VGND),
    .A1(net1484),
    .A2(net522));
 sg13g2_inv_1 _3610_ (.VDD(VPWR),
    .Y(_0117_),
    .A(net523),
    .VSS(VGND));
 sg13g2_a21oi_1 _3611_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1205),
    .A2(\s0.data_out[13][5] ),
    .Y(_1207_),
    .B1(_1168_));
 sg13g2_a21oi_1 _3612_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1017),
    .A2(_1171_),
    .Y(_1208_),
    .B1(net1381));
 sg13g2_o21ai_1 _3613_ (.B1(_1208_),
    .VDD(VPWR),
    .Y(_1209_),
    .VSS(VGND),
    .A1(net1017),
    .A2(_1207_));
 sg13g2_o21ai_1 _3614_ (.B1(_1209_),
    .VDD(VPWR),
    .Y(_1210_),
    .VSS(VGND),
    .A1(net1485),
    .A2(net684));
 sg13g2_inv_1 _3615_ (.VDD(VPWR),
    .Y(_0118_),
    .A(net685),
    .VSS(VGND));
 sg13g2_and2_1 _3616_ (.A(net1206),
    .B(\s0.data_out[13][6] ),
    .X(_1211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3617_ (.B1(net1218),
    .VDD(VPWR),
    .Y(_1212_),
    .VSS(VGND),
    .A1(_1157_),
    .A2(_1211_));
 sg13g2_nor2_1 _3618_ (.A(net1381),
    .B(_1160_),
    .Y(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3619_ (.Y(_0119_),
    .B1(_1212_),
    .B2(_1213_),
    .A2(_2820_),
    .A1(net1381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3620_ (.A(net1206),
    .B(net406),
    .X(_1214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3621_ (.B1(net1218),
    .VDD(VPWR),
    .Y(_1215_),
    .VSS(VGND),
    .A1(_1150_),
    .A2(_1214_));
 sg13g2_nor2_1 _3622_ (.A(net1381),
    .B(_1153_),
    .Y(_1216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3623_ (.Y(_0120_),
    .B1(_1215_),
    .B2(_1216_),
    .A2(_2819_),
    .A1(net1381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3624_ (.B1(net1208),
    .VDD(VPWR),
    .Y(_1217_),
    .VSS(VGND),
    .A1(net1395),
    .A2(net1196));
 sg13g2_nand2_1 _3625_ (.Y(_1218_),
    .A(net1337),
    .B(net1198),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3626_ (.Y(_1219_),
    .B(_1218_),
    .A_N(_1217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3627_ (.B1(_1219_),
    .VDD(VPWR),
    .Y(_1220_),
    .VSS(VGND),
    .A1(net1208),
    .A2(_1107_));
 sg13g2_nor2_1 _3628_ (.A(net348),
    .B(net1198),
    .Y(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3629_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1222_),
    .B(_1221_),
    .A(_1219_));
 sg13g2_nor2_1 _3630_ (.A(net1196),
    .B(_1217_),
    .Y(_1223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3631_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2734_),
    .A2(_2740_),
    .Y(_1224_),
    .B1(net1208));
 sg13g2_nor2_1 _3632_ (.A(_1223_),
    .B(_1224_),
    .Y(_1225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3633_ (.B1(net1486),
    .VDD(VPWR),
    .Y(_1226_),
    .VSS(VGND),
    .A1(net566),
    .A2(_1220_));
 sg13g2_a21oi_1 _3634_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1222_),
    .A2(_1225_),
    .Y(_0121_),
    .B1(_1226_));
 sg13g2_nor2_1 _3635_ (.A(net1382),
    .B(_1220_),
    .Y(_0122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3636_ (.A(net1490),
    .B(net342),
    .X(_0123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3637_ (.A0(\s0.data_out[13][2] ),
    .A1(\s0.data_out[12][2] ),
    .S(net1200),
    .X(_1227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3638_ (.A(net1193),
    .B_N(net1165),
    .Y(_1228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3639_ (.A2(_1227_),
    .A1(net1193),
    .B1(_1228_),
    .X(_1229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3640_ (.Y(_1230_),
    .B(\s0.data_out[12][2] ),
    .A_N(net1212),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3641_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1116_),
    .A2(_1230_),
    .Y(_1231_),
    .B1(net1204));
 sg13g2_a21oi_1 _3642_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1204),
    .A2(_1229_),
    .Y(_1232_),
    .B1(_1231_));
 sg13g2_or2_1 _3643_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1233_),
    .B(_1232_),
    .A(net1445));
 sg13g2_nand2_1 _3644_ (.Y(_1234_),
    .A(net1197),
    .B(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3645_ (.B1(_1234_),
    .VDD(VPWR),
    .Y(_1235_),
    .VSS(VGND),
    .A1(net1197),
    .A2(_2829_));
 sg13g2_nor2b_1 _3646_ (.A(net1191),
    .B_N(net1168),
    .Y(_1236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3647_ (.A2(_1235_),
    .A1(net1191),
    .B1(_1236_),
    .X(_1237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3648_ (.Y(_1238_),
    .A(_2740_),
    .B(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3649_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1124_),
    .A2(_1238_),
    .Y(_1239_),
    .B1(net1202));
 sg13g2_a21oi_1 _3650_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1202),
    .A2(_1237_),
    .Y(_1240_),
    .B1(_1239_));
 sg13g2_mux2_1 _3651_ (.A0(\s0.data_out[13][0] ),
    .A1(\s0.data_out[12][0] ),
    .S(net1197),
    .X(_1241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3652_ (.A(net1191),
    .B_N(net1171),
    .Y(_1242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3653_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1192),
    .A2(_1241_),
    .Y(_1243_),
    .B1(_1242_));
 sg13g2_nand2b_1 _3654_ (.Y(_1244_),
    .B(net1201),
    .A_N(_1243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3655_ (.A0(\s0.data_out[12][0] ),
    .A1(\s0.data_out[13][0] ),
    .S(net1210),
    .X(_1245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3656_ (.Y(_1246_),
    .B(_1245_),
    .A_N(net1201),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3657_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1246_),
    .C1(net1459),
    .B1(_1244_),
    .A1(net1454),
    .Y(_1247_),
    .A2(_1240_));
 sg13g2_o21ai_1 _3658_ (.B1(_1233_),
    .VDD(VPWR),
    .Y(_1248_),
    .VSS(VGND),
    .A1(net1454),
    .A2(_1240_));
 sg13g2_nand2_1 _3659_ (.Y(_1249_),
    .A(net1197),
    .B(net467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3660_ (.B1(_1249_),
    .VDD(VPWR),
    .Y(_1250_),
    .VSS(VGND),
    .A1(net1197),
    .A2(_2827_));
 sg13g2_nor2_1 _3661_ (.A(net1192),
    .B(net994),
    .Y(_1251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3662_ (.A2(_1250_),
    .A1(net1193),
    .B1(_1251_),
    .X(_1252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3663_ (.Y(_1253_),
    .A(_2740_),
    .B(net467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3664_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1139_),
    .A2(_1253_),
    .Y(_1254_),
    .B1(net1204));
 sg13g2_a21oi_1 _3665_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1204),
    .A2(_1252_),
    .Y(_1255_),
    .B1(_1254_));
 sg13g2_a22oi_1 _3666_ (.Y(_1256_),
    .B1(_1255_),
    .B2(net1440),
    .A2(_1232_),
    .A1(net1445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3667_ (.B1(_1256_),
    .VDD(VPWR),
    .Y(_1257_),
    .VSS(VGND),
    .A1(_1247_),
    .A2(_1248_));
 sg13g2_nand2_1 _3668_ (.Y(_1258_),
    .A(net1199),
    .B(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3669_ (.A0(\s0.data_out[13][7] ),
    .A1(\s0.data_out[12][7] ),
    .S(net1198),
    .X(_1259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3670_ (.A(net1194),
    .B_N(net1145),
    .Y(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3671_ (.A2(_1259_),
    .A1(net1194),
    .B1(_1260_),
    .X(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3672_ (.Y(_1262_),
    .B(\s0.data_out[12][7] ),
    .A_N(net1212),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3673_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1148_),
    .A2(_1262_),
    .Y(_1263_),
    .B1(net1206));
 sg13g2_a21oi_1 _3674_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1207),
    .A2(_1261_),
    .Y(_1264_),
    .B1(_1263_));
 sg13g2_nand2_1 _3675_ (.Y(_1265_),
    .A(net1199),
    .B(net619),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3676_ (.A0(\s0.data_out[13][6] ),
    .A1(\s0.data_out[12][6] ),
    .S(net1199),
    .X(_1266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3677_ (.A(net1194),
    .B_N(net1150),
    .Y(_1267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3678_ (.A2(_1266_),
    .A1(net1194),
    .B1(_1267_),
    .X(_1268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3679_ (.Y(_1269_),
    .B(\s0.data_out[12][6] ),
    .A_N(net1212),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3680_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1155_),
    .A2(_1269_),
    .Y(_1270_),
    .B1(net1206));
 sg13g2_a21oi_1 _3681_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1207),
    .A2(_1268_),
    .Y(_1271_),
    .B1(_1270_));
 sg13g2_a22oi_1 _3682_ (.Y(_1272_),
    .B1(_1271_),
    .B2(net1413),
    .A2(_1264_),
    .A1(net1404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3683_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1273_),
    .B(_1271_),
    .A(net1413));
 sg13g2_or2_1 _3684_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1274_),
    .B(_1264_),
    .A(net1404));
 sg13g2_and3_1 _3685_ (.X(_1275_),
    .A(_1272_),
    .B(_1273_),
    .C(_1274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3686_ (.A0(\s0.data_out[13][5] ),
    .A1(\s0.data_out[12][5] ),
    .S(net1198),
    .X(_1276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3687_ (.A(net1194),
    .B_N(net1154),
    .Y(_1277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3688_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1194),
    .A2(_1276_),
    .Y(_1278_),
    .B1(_1277_));
 sg13g2_nand2b_1 _3689_ (.Y(_1279_),
    .B(net1207),
    .A_N(_1278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3690_ (.A0(\s0.data_out[12][5] ),
    .A1(\s0.data_out[13][5] ),
    .S(net1212),
    .X(_1280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3691_ (.Y(_1281_),
    .B(_1280_),
    .A_N(net1207),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3692_ (.B(_1279_),
    .C(_1281_),
    .A(net1423),
    .Y(_1282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3693_ (.Y(_1283_),
    .A(net1198),
    .B(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3694_ (.A0(\s0.data_out[13][4] ),
    .A1(\s0.data_out[12][4] ),
    .S(net1198),
    .X(_1284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3695_ (.A(net1196),
    .B_N(net1159),
    .Y(_1285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3696_ (.A2(_1284_),
    .A1(net1196),
    .B1(_1285_),
    .X(_1286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3697_ (.Y(_1287_),
    .B(net414),
    .A_N(net1211),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3698_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1177_),
    .A2(_1287_),
    .Y(_1288_),
    .B1(net1205));
 sg13g2_a21oi_1 _3699_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1205),
    .A2(_1286_),
    .Y(_1289_),
    .B1(_1288_));
 sg13g2_nand2_1 _3700_ (.Y(_1290_),
    .A(net1432),
    .B(_1289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3701_ (.Y(_1291_),
    .A(_1282_),
    .B(_1290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3702_ (.A(net1440),
    .B(_1255_),
    .Y(_1292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3703_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1279_),
    .A2(_1281_),
    .Y(_1293_),
    .B1(net1423));
 sg13g2_nor2_1 _3704_ (.A(net1432),
    .B(_1289_),
    .Y(_1294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3705_ (.A(_1291_),
    .B(_1292_),
    .C(_1293_),
    .D(_1294_),
    .Y(_1295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3706_ (.B(_1275_),
    .C(_1295_),
    .A(_1257_),
    .Y(_1296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3707_ (.B1(_1282_),
    .VDD(VPWR),
    .Y(_1297_),
    .VSS(VGND),
    .A1(_1290_),
    .A2(_1293_));
 sg13g2_and2_1 _3708_ (.A(_1275_),
    .B(_1297_),
    .X(_1298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3709_ (.A(_1272_),
    .B_N(_1274_),
    .Y(_1299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3710_ (.A(_1220_),
    .B(_1298_),
    .C(_1299_),
    .Y(_1300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3711_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1301_),
    .B(net1332),
    .A(net343));
 sg13g2_a21oi_1 _3712_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1296_),
    .A2(_1300_),
    .Y(_0124_),
    .B1(_1301_));
 sg13g2_and2_1 _3713_ (.A(net1191),
    .B(\s0.data_out[12][0] ),
    .X(_1302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3714_ (.B1(net1202),
    .VDD(VPWR),
    .Y(_1303_),
    .VSS(VGND),
    .A1(_1242_),
    .A2(_1302_));
 sg13g2_nand3_1 _3715_ (.B(_1246_),
    .C(_1303_),
    .A(net1484),
    .Y(_1304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3716_ (.B1(_1304_),
    .VDD(VPWR),
    .Y(_1305_),
    .VSS(VGND),
    .A1(net1487),
    .A2(net679));
 sg13g2_inv_1 _3717_ (.VDD(VPWR),
    .Y(_0125_),
    .A(_1305_),
    .VSS(VGND));
 sg13g2_nor2_1 _3718_ (.A(net1016),
    .B(_2833_),
    .Y(_1306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3719_ (.B1(net1202),
    .VDD(VPWR),
    .Y(_1307_),
    .VSS(VGND),
    .A1(_1236_),
    .A2(_1306_));
 sg13g2_nor2_1 _3720_ (.A(net1378),
    .B(_1239_),
    .Y(_1308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3721_ (.Y(_0126_),
    .B1(_1307_),
    .B2(_1308_),
    .A2(_2829_),
    .A1(net1378),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3722_ (.A(net1193),
    .B(\s0.data_out[12][2] ),
    .X(_1309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3723_ (.B1(net1204),
    .VDD(VPWR),
    .Y(_1310_),
    .VSS(VGND),
    .A1(_1228_),
    .A2(_1309_));
 sg13g2_nor2_1 _3724_ (.A(net1379),
    .B(_1231_),
    .Y(_1311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3725_ (.Y(_0127_),
    .B1(_1310_),
    .B2(_1311_),
    .A2(_2828_),
    .A1(net1379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3726_ (.A(net1016),
    .B(_2832_),
    .Y(_1312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3727_ (.B1(net1209),
    .VDD(VPWR),
    .Y(_1313_),
    .VSS(VGND),
    .A1(_1251_),
    .A2(_1312_));
 sg13g2_nor2_1 _3728_ (.A(net1379),
    .B(_1254_),
    .Y(_1314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3729_ (.Y(_0128_),
    .B1(_1313_),
    .B2(_1314_),
    .A2(_2827_),
    .A1(net1379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3730_ (.A(net1196),
    .B(net414),
    .X(_1315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3731_ (.B1(net1205),
    .VDD(VPWR),
    .Y(_1316_),
    .VSS(VGND),
    .A1(_1285_),
    .A2(_1315_));
 sg13g2_nor2_1 _3732_ (.A(net1382),
    .B(net415),
    .Y(_1317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3733_ (.Y(_0129_),
    .B1(_1316_),
    .B2(_1317_),
    .A2(_2826_),
    .A1(net1381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3734_ (.A(net1194),
    .B(\s0.data_out[12][5] ),
    .X(_1318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3735_ (.B1(net1207),
    .VDD(VPWR),
    .Y(_1319_),
    .VSS(VGND),
    .A1(_1277_),
    .A2(_1318_));
 sg13g2_nand3_1 _3736_ (.B(_1281_),
    .C(_1319_),
    .A(net1486),
    .Y(_1320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3737_ (.B1(_1320_),
    .VDD(VPWR),
    .Y(_1321_),
    .VSS(VGND),
    .A1(net1486),
    .A2(net686));
 sg13g2_inv_1 _3738_ (.VDD(VPWR),
    .Y(_0130_),
    .A(_1321_),
    .VSS(VGND));
 sg13g2_nor2_1 _3739_ (.A(net1015),
    .B(_2831_),
    .Y(_1322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3740_ (.B1(net1207),
    .VDD(VPWR),
    .Y(_1323_),
    .VSS(VGND),
    .A1(_1267_),
    .A2(_1322_));
 sg13g2_nand3b_1 _3741_ (.B(_1323_),
    .C(net1486),
    .Y(_1324_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1270_));
 sg13g2_o21ai_1 _3742_ (.B1(_1324_),
    .VDD(VPWR),
    .Y(_1325_),
    .VSS(VGND),
    .A1(net1486),
    .A2(net550));
 sg13g2_inv_1 _3743_ (.VDD(VPWR),
    .Y(_0131_),
    .A(net551),
    .VSS(VGND));
 sg13g2_nor2_1 _3744_ (.A(net1015),
    .B(_2830_),
    .Y(_1326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3745_ (.B1(net1207),
    .VDD(VPWR),
    .Y(_1327_),
    .VSS(VGND),
    .A1(_1260_),
    .A2(_1326_));
 sg13g2_nor2_1 _3746_ (.A(net1382),
    .B(_1263_),
    .Y(_1328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3747_ (.Y(_0132_),
    .B1(_1327_),
    .B2(_1328_),
    .A2(_2825_),
    .A1(net1382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3748_ (.B1(net1196),
    .VDD(VPWR),
    .Y(_1329_),
    .VSS(VGND),
    .A1(net1395),
    .A2(net1183));
 sg13g2_nor2_1 _3749_ (.A(net1395),
    .B(_2745_),
    .Y(_1330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3750_ (.A(_1329_),
    .B(_1330_),
    .Y(_1331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3751_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1015),
    .A2(_1218_),
    .Y(_1332_),
    .B1(_1331_));
 sg13g2_o21ai_1 _3752_ (.B1(_1331_),
    .VDD(VPWR),
    .Y(_1333_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[11] [0]),
    .A2(net1188));
 sg13g2_nor2_1 _3753_ (.A(net1183),
    .B(_1329_),
    .Y(_1334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3754_ (.B1(net1015),
    .VDD(VPWR),
    .Y(_1335_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[11] [0]),
    .A2(net1198));
 sg13g2_nand2_1 _3755_ (.Y(_1336_),
    .A(_1333_),
    .B(_1335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3756_ (.B1(net1485),
    .VDD(VPWR),
    .Y(_1337_),
    .VSS(VGND),
    .A1(_1334_),
    .A2(_1336_));
 sg13g2_a21oi_1 _3757_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2734_),
    .A2(_1332_),
    .Y(_0133_),
    .B1(_1337_));
 sg13g2_and2_1 _3758_ (.A(net1485),
    .B(_1332_),
    .X(_0134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3759_ (.Y(_1338_),
    .A(net1187),
    .B(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3760_ (.A0(\s0.data_out[12][1] ),
    .A1(\s0.data_out[11][1] ),
    .S(net1187),
    .X(_1339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3761_ (.A(net1178),
    .B_N(net1168),
    .Y(_1340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3762_ (.A2(_1339_),
    .A1(net1178),
    .B1(_1340_),
    .X(_1341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3763_ (.Y(_1342_),
    .B(\s0.data_out[11][1] ),
    .A_N(net1197),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3764_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1234_),
    .A2(_1342_),
    .Y(_1343_),
    .B1(net1191));
 sg13g2_a21oi_1 _3765_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1192),
    .A2(_1341_),
    .Y(_1344_),
    .B1(_1343_));
 sg13g2_mux2_1 _3766_ (.A0(\s0.data_out[11][0] ),
    .A1(\s0.data_out[12][0] ),
    .S(net1197),
    .X(_1345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3767_ (.Y(_1346_),
    .A(net1016),
    .B(_1345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3768_ (.A(net1178),
    .B_N(net1171),
    .Y(_1347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3769_ (.A0(\s0.data_out[12][0] ),
    .A1(\s0.data_out[11][0] ),
    .S(net1187),
    .X(_1348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3770_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1178),
    .A2(_1348_),
    .Y(_1349_),
    .B1(_1347_));
 sg13g2_nand2b_1 _3771_ (.Y(_1350_),
    .B(net1191),
    .A_N(_1349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3772_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1350_),
    .C1(net1459),
    .B1(_1346_),
    .A1(net1455),
    .Y(_1351_),
    .A2(_1344_));
 sg13g2_nand2_1 _3773_ (.Y(_1352_),
    .A(net1190),
    .B(net422),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3774_ (.A0(\s0.data_out[12][2] ),
    .A1(\s0.data_out[11][2] ),
    .S(net1187),
    .X(_1353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3775_ (.A(net1180),
    .B_N(net1164),
    .Y(_1354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1180),
    .A2(_1353_),
    .Y(_1355_),
    .B1(_1354_));
 sg13g2_mux2_1 _3777_ (.A0(\s0.data_out[11][2] ),
    .A1(\s0.data_out[12][2] ),
    .S(net1200),
    .X(_1356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3778_ (.Y(_1357_),
    .A(net1016),
    .B(_1356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3779_ (.B1(_1357_),
    .VDD(VPWR),
    .Y(_1358_),
    .VSS(VGND),
    .A1(net1016),
    .A2(_1355_));
 sg13g2_or2_1 _3780_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1359_),
    .B(_1358_),
    .A(net1335));
 sg13g2_xnor2_1 _3781_ (.Y(_1360_),
    .A(net1335),
    .B(_1358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3782_ (.A(net1455),
    .B(_1344_),
    .Y(_1361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3783_ (.Y(_1362_),
    .A(net1187),
    .B(net461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3784_ (.A0(\s0.data_out[12][3] ),
    .A1(\s0.data_out[11][3] ),
    .S(net1187),
    .X(_1363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3785_ (.A(net1180),
    .B_N(net1161),
    .Y(_1364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3786_ (.A2(_1363_),
    .A1(net1180),
    .B1(_1364_),
    .X(_1365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3787_ (.Y(_1366_),
    .B(net461),
    .A_N(net1197),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3788_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1249_),
    .A2(_1366_),
    .Y(_1367_),
    .B1(net1193));
 sg13g2_a21oi_1 _3789_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1193),
    .A2(_1365_),
    .Y(_1368_),
    .B1(_1367_));
 sg13g2_nor2_1 _3790_ (.A(net1440),
    .B(_1368_),
    .Y(_1369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3791_ (.A(_1351_),
    .B(_1360_),
    .C(_1361_),
    .D(_1369_),
    .Y(_1370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3792_ (.Y(_1371_),
    .A(net1440),
    .B(_1368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3793_ (.B1(_1371_),
    .VDD(VPWR),
    .Y(_1372_),
    .VSS(VGND),
    .A1(_1359_),
    .A2(_1369_));
 sg13g2_nor2_1 _3794_ (.A(_1370_),
    .B(_1372_),
    .Y(_1373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3795_ (.Y(_1374_),
    .A(net1188),
    .B(net451),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3796_ (.A0(\s0.data_out[12][7] ),
    .A1(\s0.data_out[11][7] ),
    .S(net1188),
    .X(_1375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3797_ (.A(net1182),
    .B_N(net1144),
    .Y(_1376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3798_ (.A2(_1375_),
    .A1(net1182),
    .B1(_1376_),
    .X(_1377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3799_ (.Y(_1378_),
    .B(net451),
    .A_N(net1199),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3800_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1258_),
    .A2(_1378_),
    .Y(_1379_),
    .B1(net1195));
 sg13g2_a21oi_1 _3801_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1195),
    .A2(_1377_),
    .Y(_1380_),
    .B1(_1379_));
 sg13g2_nand2_1 _3802_ (.Y(_1381_),
    .A(net1188),
    .B(\s0.data_out[11][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3803_ (.A0(\s0.data_out[12][6] ),
    .A1(\s0.data_out[11][6] ),
    .S(net1188),
    .X(_1382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3804_ (.A(net1182),
    .B_N(net1149),
    .Y(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3805_ (.A2(_1382_),
    .A1(net1182),
    .B1(_1383_),
    .X(_1384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3806_ (.Y(_1385_),
    .B(\s0.data_out[11][6] ),
    .A_N(net1199),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3807_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1265_),
    .A2(_1385_),
    .Y(_1386_),
    .B1(net1194));
 sg13g2_a21oi_1 _3808_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1195),
    .A2(_1384_),
    .Y(_1387_),
    .B1(_1386_));
 sg13g2_a22oi_1 _3809_ (.Y(_1388_),
    .B1(_1387_),
    .B2(net1413),
    .A2(_1380_),
    .A1(net1404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3810_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1389_),
    .B(_1387_),
    .A(net1413));
 sg13g2_nor2_1 _3811_ (.A(net1404),
    .B(_1380_),
    .Y(_1390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3812_ (.B(_1388_),
    .C(_1389_),
    .Y(_1391_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1390_));
 sg13g2_nor2b_1 _3813_ (.A(net1183),
    .B_N(net1158),
    .Y(_1392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3814_ (.Y(_1393_),
    .A(net1188),
    .B(net373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3815_ (.A0(\s0.data_out[12][4] ),
    .A1(\s0.data_out[11][4] ),
    .S(net1188),
    .X(_1394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3816_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1183),
    .A2(_1394_),
    .Y(_1395_),
    .B1(_1392_));
 sg13g2_nand2b_1 _3817_ (.Y(_1396_),
    .B(net1196),
    .A_N(_1395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3818_ (.B1(_1283_),
    .VDD(VPWR),
    .Y(_1397_),
    .VSS(VGND),
    .A1(net1198),
    .A2(_2835_));
 sg13g2_nand2_1 _3819_ (.Y(_1398_),
    .A(net1015),
    .B(_1397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3820_ (.B(_1396_),
    .C(_1398_),
    .A(net1432),
    .Y(_1399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3821_ (.A0(\s0.data_out[12][5] ),
    .A1(\s0.data_out[11][5] ),
    .S(net1188),
    .X(_1400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3822_ (.A(net1186),
    .B_N(net1153),
    .Y(_1401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1182),
    .A2(_1400_),
    .Y(_1402_),
    .B1(_1401_));
 sg13g2_nand2b_1 _3824_ (.Y(_1403_),
    .B(net1195),
    .A_N(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3825_ (.A0(\s0.data_out[11][5] ),
    .A1(\s0.data_out[12][5] ),
    .S(net1199),
    .X(_1404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3826_ (.Y(_1405_),
    .A(net1015),
    .B(_1404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3827_ (.B(_1403_),
    .C(_1405_),
    .A(net1423),
    .Y(_1406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3828_ (.Y(_1407_),
    .A(_1399_),
    .B(_1406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3829_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1396_),
    .A2(_1398_),
    .Y(_1408_),
    .B1(net1432));
 sg13g2_a21oi_1 _3830_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1403_),
    .A2(_1405_),
    .Y(_1409_),
    .B1(net1423));
 sg13g2_or2_1 _3831_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1410_),
    .B(_1409_),
    .A(_1408_));
 sg13g2_or4_1 _3832_ (.A(_1373_),
    .B(_1391_),
    .C(_1407_),
    .D(_1410_),
    .X(_1411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3833_ (.B1(_1406_),
    .VDD(VPWR),
    .Y(_1412_),
    .VSS(VGND),
    .A1(_1399_),
    .A2(_1409_));
 sg13g2_nor2b_1 _3834_ (.A(_1391_),
    .B_N(_1412_),
    .Y(_1413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3835_ (.B1(_1332_),
    .VDD(VPWR),
    .Y(_1414_),
    .VSS(VGND),
    .A1(_1388_),
    .A2(_1390_));
 sg13g2_nor2_1 _3836_ (.A(_1413_),
    .B(_1414_),
    .Y(_1415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3837_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1416_),
    .B(net1331),
    .A(net342));
 sg13g2_a21oi_1 _3838_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1411_),
    .A2(_1415_),
    .Y(_0135_),
    .B1(_1416_));
 sg13g2_and2_1 _3839_ (.A(net1178),
    .B(\s0.data_out[11][0] ),
    .X(_1417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3840_ (.B1(net1191),
    .VDD(VPWR),
    .Y(_1418_),
    .VSS(VGND),
    .A1(_1347_),
    .A2(_1417_));
 sg13g2_nand3_1 _3841_ (.B(_1346_),
    .C(_1418_),
    .A(net1484),
    .Y(_1419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3842_ (.B1(_1419_),
    .VDD(VPWR),
    .Y(_1420_),
    .VSS(VGND),
    .A1(net1484),
    .A2(net621));
 sg13g2_inv_1 _3843_ (.VDD(VPWR),
    .Y(_0136_),
    .A(_1420_),
    .VSS(VGND));
 sg13g2_and2_1 _3844_ (.A(net1178),
    .B(\s0.data_out[11][1] ),
    .X(_1421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3845_ (.B1(net1191),
    .VDD(VPWR),
    .Y(_1422_),
    .VSS(VGND),
    .A1(_1340_),
    .A2(_1421_));
 sg13g2_nor2_1 _3846_ (.A(net1379),
    .B(_1343_),
    .Y(_1423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3847_ (.Y(_0137_),
    .B1(_1422_),
    .B2(_1423_),
    .A2(_2833_),
    .A1(net1378),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3848_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1180),
    .A2(net422),
    .Y(_1424_),
    .B1(_1354_));
 sg13g2_a21oi_1 _3849_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1016),
    .A2(_1356_),
    .Y(_1425_),
    .B1(net1385));
 sg13g2_o21ai_1 _3850_ (.B1(_1425_),
    .VDD(VPWR),
    .Y(_1426_),
    .VSS(VGND),
    .A1(net1016),
    .A2(_1424_));
 sg13g2_o21ai_1 _3851_ (.B1(_1426_),
    .VDD(VPWR),
    .Y(_1427_),
    .VSS(VGND),
    .A1(net1488),
    .A2(net651));
 sg13g2_inv_1 _3852_ (.VDD(VPWR),
    .Y(_0138_),
    .A(_1427_),
    .VSS(VGND));
 sg13g2_and2_1 _3853_ (.A(net1180),
    .B(net461),
    .X(_1428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3854_ (.B1(net1193),
    .VDD(VPWR),
    .Y(_1429_),
    .VSS(VGND),
    .A1(_1364_),
    .A2(_1428_));
 sg13g2_nor2_1 _3855_ (.A(net1379),
    .B(_1367_),
    .Y(_1430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3856_ (.Y(_0139_),
    .B1(_1429_),
    .B2(_1430_),
    .A2(_2832_),
    .A1(net1379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3857_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1183),
    .A2(net373),
    .Y(_1431_),
    .B1(_1392_));
 sg13g2_a21oi_1 _3858_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1015),
    .A2(_1397_),
    .Y(_1432_),
    .B1(net1386));
 sg13g2_o21ai_1 _3859_ (.B1(_1432_),
    .VDD(VPWR),
    .Y(_1433_),
    .VSS(VGND),
    .A1(net1015),
    .A2(_1431_));
 sg13g2_o21ai_1 _3860_ (.B1(_1433_),
    .VDD(VPWR),
    .Y(_1434_),
    .VSS(VGND),
    .A1(net1486),
    .A2(net414));
 sg13g2_inv_1 _3861_ (.VDD(VPWR),
    .Y(_0140_),
    .A(_1434_),
    .VSS(VGND));
 sg13g2_a21oi_1 _3862_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1182),
    .A2(\s0.data_out[11][5] ),
    .Y(_1435_),
    .B1(_1401_));
 sg13g2_a21oi_1 _3863_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2744_),
    .A2(_1404_),
    .Y(_1436_),
    .B1(net1386));
 sg13g2_o21ai_1 _3864_ (.B1(_1436_),
    .VDD(VPWR),
    .Y(_1437_),
    .VSS(VGND),
    .A1(_2744_),
    .A2(_1435_));
 sg13g2_o21ai_1 _3865_ (.B1(_1437_),
    .VDD(VPWR),
    .Y(_1438_),
    .VSS(VGND),
    .A1(net1490),
    .A2(net616));
 sg13g2_inv_1 _3866_ (.VDD(VPWR),
    .Y(_0141_),
    .A(net617),
    .VSS(VGND));
 sg13g2_and2_1 _3867_ (.A(net1182),
    .B(\s0.data_out[11][6] ),
    .X(_1439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3868_ (.B1(net1195),
    .VDD(VPWR),
    .Y(_1440_),
    .VSS(VGND),
    .A1(_1383_),
    .A2(_1439_));
 sg13g2_nor2_1 _3869_ (.A(net1381),
    .B(_1386_),
    .Y(_1441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3870_ (.Y(_0142_),
    .B1(_1440_),
    .B2(_1441_),
    .A2(_2831_),
    .A1(net1382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3871_ (.A(net1182),
    .B(net451),
    .X(_1442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3872_ (.B1(net1195),
    .VDD(VPWR),
    .Y(_1443_),
    .VSS(VGND),
    .A1(_1376_),
    .A2(_1442_));
 sg13g2_nor2_1 _3873_ (.A(net1382),
    .B(_1379_),
    .Y(_1444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3874_ (.Y(_0143_),
    .B1(_1443_),
    .B2(_1444_),
    .A2(_2830_),
    .A1(net1382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3875_ (.B1(net1185),
    .VDD(VPWR),
    .Y(_1445_),
    .VSS(VGND),
    .A1(net1395),
    .A2(net1140));
 sg13g2_nand2_1 _3876_ (.Y(_1446_),
    .A(net1338),
    .B(net1175),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3877_ (.Y(_1447_),
    .B(_1446_),
    .A_N(_1445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3878_ (.B1(_1447_),
    .VDD(VPWR),
    .Y(_1448_),
    .VSS(VGND),
    .A1(net1185),
    .A2(_1330_));
 sg13g2_nor2_1 _3879_ (.A(net350),
    .B(net1176),
    .Y(_1449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3880_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1450_),
    .B(_1449_),
    .A(_1447_));
 sg13g2_nor2_1 _3881_ (.A(net1140),
    .B(_1445_),
    .Y(_1451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3882_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2733_),
    .A2(_2745_),
    .Y(_1452_),
    .B1(net1185));
 sg13g2_nor2_1 _3883_ (.A(_1451_),
    .B(_1452_),
    .Y(_1453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3884_ (.B1(net1490),
    .VDD(VPWR),
    .Y(_1454_),
    .VSS(VGND),
    .A1(net644),
    .A2(_1448_));
 sg13g2_a21oi_1 _3885_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1450_),
    .A2(_1453_),
    .Y(_0144_),
    .B1(_1454_));
 sg13g2_nor2_1 _3886_ (.A(net1386),
    .B(_1448_),
    .Y(_0145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3887_ (.A(net1490),
    .B(net341),
    .X(_0146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3888_ (.A(net1490),
    .B(net329),
    .X(_0147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3889_ (.A0(\s0.data_out[11][2] ),
    .A1(\s0.data_out[10][2] ),
    .S(net1174),
    .X(_1455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3890_ (.A(net1136),
    .B_N(net1164),
    .Y(_1456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3891_ (.A2(_1455_),
    .A1(net1136),
    .B1(_1456_),
    .X(_1457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3892_ (.Y(_1458_),
    .B(\s0.data_out[10][2] ),
    .A_N(net1190),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3893_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1352_),
    .A2(_1458_),
    .Y(_1459_),
    .B1(net1181));
 sg13g2_a21oi_1 _3894_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1181),
    .A2(_1457_),
    .Y(_1460_),
    .B1(_1459_));
 sg13g2_or2_1 _3895_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1461_),
    .B(_1460_),
    .A(net1445));
 sg13g2_nand2_1 _3896_ (.Y(_1462_),
    .A(net1174),
    .B(net489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3897_ (.B1(_1462_),
    .VDD(VPWR),
    .Y(_1463_),
    .VSS(VGND),
    .A1(net1174),
    .A2(_2838_));
 sg13g2_nor2b_1 _3898_ (.A(net1135),
    .B_N(net1168),
    .Y(_1464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3899_ (.A2(_1463_),
    .A1(net1136),
    .B1(_1464_),
    .X(_1465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3900_ (.Y(_1466_),
    .A(_2745_),
    .B(net489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3901_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1338_),
    .A2(_1466_),
    .Y(_1467_),
    .B1(net1178));
 sg13g2_a21oi_1 _3902_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1179),
    .A2(_1465_),
    .Y(_1468_),
    .B1(_1467_));
 sg13g2_mux2_1 _3903_ (.A0(\s0.data_out[11][0] ),
    .A1(\s0.data_out[10][0] ),
    .S(net1174),
    .X(_1469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3904_ (.A(net1135),
    .B_N(net1171),
    .Y(_1470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3905_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1135),
    .A2(_1469_),
    .Y(_1471_),
    .B1(_1470_));
 sg13g2_nand2b_1 _3906_ (.Y(_1472_),
    .B(net1179),
    .A_N(_1471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3907_ (.A0(\s0.data_out[10][0] ),
    .A1(\s0.data_out[11][0] ),
    .S(net1187),
    .X(_1473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3908_ (.Y(_1474_),
    .B(_1473_),
    .A_N(net1179),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3909_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1474_),
    .C1(net1459),
    .B1(_1472_),
    .A1(net1454),
    .Y(_1475_),
    .A2(_1468_));
 sg13g2_o21ai_1 _3910_ (.B1(_1461_),
    .VDD(VPWR),
    .Y(_1476_),
    .VSS(VGND),
    .A1(net1454),
    .A2(_1468_));
 sg13g2_nand2_1 _3911_ (.Y(_1477_),
    .A(net1177),
    .B(net477),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3912_ (.A0(\s0.data_out[11][3] ),
    .A1(\s0.data_out[10][3] ),
    .S(net1177),
    .X(_1478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3913_ (.A(net1136),
    .B_N(net1161),
    .Y(_1479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3914_ (.A2(_1478_),
    .A1(net1137),
    .B1(_1479_),
    .X(_1480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3915_ (.Y(_1481_),
    .B(\s0.data_out[10][3] ),
    .A_N(net1190),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3916_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1362_),
    .A2(_1481_),
    .Y(_1482_),
    .B1(net1181));
 sg13g2_a21oi_1 _3917_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1181),
    .A2(_1480_),
    .Y(_1483_),
    .B1(_1482_));
 sg13g2_a22oi_1 _3918_ (.Y(_1484_),
    .B1(_1483_),
    .B2(net1441),
    .A2(_1460_),
    .A1(net1445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3919_ (.B1(_1484_),
    .VDD(VPWR),
    .Y(_1485_),
    .VSS(VGND),
    .A1(_1475_),
    .A2(_1476_));
 sg13g2_nand2_1 _3920_ (.Y(_1486_),
    .A(net1175),
    .B(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3921_ (.A0(\s0.data_out[11][7] ),
    .A1(\s0.data_out[10][7] ),
    .S(net1175),
    .X(_1487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3922_ (.A(net1138),
    .B_N(net1144),
    .Y(_1488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3923_ (.A2(_1487_),
    .A1(net1138),
    .B1(_1488_),
    .X(_1489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3924_ (.Y(_1490_),
    .B(\s0.data_out[10][7] ),
    .A_N(net1189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3925_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1374_),
    .A2(_1490_),
    .Y(_1491_),
    .B1(net1185));
 sg13g2_a21oi_1 _3926_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1184),
    .A2(_1489_),
    .Y(_1492_),
    .B1(_1491_));
 sg13g2_nand2_1 _3927_ (.Y(_1493_),
    .A(net1175),
    .B(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3928_ (.A0(\s0.data_out[11][6] ),
    .A1(\s0.data_out[10][6] ),
    .S(net1176),
    .X(_1494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3929_ (.A(net1138),
    .B_N(net1149),
    .Y(_1495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3930_ (.A2(_1494_),
    .A1(net1138),
    .B1(_1495_),
    .X(_1496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3931_ (.Y(_1497_),
    .B(net636),
    .A_N(net1189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3932_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1381_),
    .A2(_1497_),
    .Y(_1498_),
    .B1(net1184));
 sg13g2_a21oi_1 _3933_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1184),
    .A2(_1496_),
    .Y(_1499_),
    .B1(_1498_));
 sg13g2_a22oi_1 _3934_ (.Y(_1500_),
    .B1(_1499_),
    .B2(net1414),
    .A2(_1492_),
    .A1(net1405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3935_ (.A(net1414),
    .B(_1499_),
    .Y(_1501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3936_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1502_),
    .B(_1492_),
    .A(net1405));
 sg13g2_nand3b_1 _3937_ (.B(_1502_),
    .C(_1500_),
    .Y(_1503_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1501_));
 sg13g2_mux2_1 _3938_ (.A0(\s0.data_out[11][5] ),
    .A1(\s0.data_out[10][5] ),
    .S(net1176),
    .X(_1504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3939_ (.A(net1140),
    .B_N(net1153),
    .Y(_1505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3940_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1140),
    .A2(_1504_),
    .Y(_1506_),
    .B1(_1505_));
 sg13g2_nand2b_1 _3941_ (.Y(_1507_),
    .B(net1184),
    .A_N(_1506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3942_ (.A0(\s0.data_out[10][5] ),
    .A1(\s0.data_out[11][5] ),
    .S(net1189),
    .X(_1508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3943_ (.Y(_1509_),
    .B(_1508_),
    .A_N(net1184),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3944_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1507_),
    .A2(_1509_),
    .Y(_1510_),
    .B1(net1424));
 sg13g2_mux2_1 _3945_ (.A0(\s0.data_out[11][4] ),
    .A1(\s0.data_out[10][4] ),
    .S(net1176),
    .X(_1511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3946_ (.A(net1140),
    .B_N(net1158),
    .Y(_1512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3947_ (.A2(_1511_),
    .A1(net1140),
    .B1(_1512_),
    .X(_1513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3948_ (.Y(_1514_),
    .B(\s0.data_out[10][4] ),
    .A_N(net1189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3949_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1393_),
    .A2(_1514_),
    .Y(_1515_),
    .B1(net1183));
 sg13g2_a21oi_1 _3950_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1185),
    .A2(_1513_),
    .Y(_1516_),
    .B1(_1515_));
 sg13g2_nor2_1 _3951_ (.A(net1432),
    .B(_1516_),
    .Y(_1517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3952_ (.Y(_1518_),
    .A(net1432),
    .B(_1516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3953_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1519_),
    .B(_1483_),
    .A(net1441));
 sg13g2_nand3_1 _3954_ (.B(_1507_),
    .C(_1509_),
    .A(net1424),
    .Y(_1520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3955_ (.B(_1519_),
    .C(_1520_),
    .A(_1518_),
    .Y(_1521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3956_ (.A(_1503_),
    .B(_1510_),
    .C(_1517_),
    .D(_1521_),
    .Y(_1522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3957_ (.Y(_1523_),
    .A(_1485_),
    .B(_1522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3958_ (.B1(_1520_),
    .VDD(VPWR),
    .Y(_1524_),
    .VSS(VGND),
    .A1(_1510_),
    .A2(_1518_));
 sg13g2_nor2b_1 _3959_ (.A(_1503_),
    .B_N(_1524_),
    .Y(_1525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3960_ (.A(_1500_),
    .B_N(_1502_),
    .Y(_1526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3961_ (.A(_1448_),
    .B(_1525_),
    .C(_1526_),
    .Y(_1527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3962_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1528_),
    .B(net1331),
    .A(net341));
 sg13g2_a21oi_1 _3963_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1523_),
    .A2(_1527_),
    .Y(_0148_),
    .B1(_1528_));
 sg13g2_and2_1 _3964_ (.A(net1135),
    .B(\s0.data_out[10][0] ),
    .X(_1529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3965_ (.B1(net1179),
    .VDD(VPWR),
    .Y(_1530_),
    .VSS(VGND),
    .A1(_1470_),
    .A2(_1529_));
 sg13g2_nand3_1 _3966_ (.B(_1474_),
    .C(_1530_),
    .A(net1488),
    .Y(_1531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3967_ (.B1(_1531_),
    .VDD(VPWR),
    .Y(_1532_),
    .VSS(VGND),
    .A1(net1488),
    .A2(net661));
 sg13g2_inv_1 _3968_ (.VDD(VPWR),
    .Y(_0149_),
    .A(_1532_),
    .VSS(VGND));
 sg13g2_nor2_1 _3969_ (.A(net1014),
    .B(_2839_),
    .Y(_1533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3970_ (.B1(net1178),
    .VDD(VPWR),
    .Y(_1534_),
    .VSS(VGND),
    .A1(_1464_),
    .A2(_1533_));
 sg13g2_nor2_1 _3971_ (.A(net1385),
    .B(_1467_),
    .Y(_1535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3972_ (.Y(_0150_),
    .B1(_1534_),
    .B2(_1535_),
    .A2(_2838_),
    .A1(net1385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3973_ (.A(net1136),
    .B(\s0.data_out[10][2] ),
    .X(_1536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3974_ (.B1(net1181),
    .VDD(VPWR),
    .Y(_1537_),
    .VSS(VGND),
    .A1(_1456_),
    .A2(_1536_));
 sg13g2_nor2_1 _3975_ (.A(net1385),
    .B(_1459_),
    .Y(_1538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3976_ (.Y(_0151_),
    .B1(_1537_),
    .B2(_1538_),
    .A2(_2837_),
    .A1(net1385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3977_ (.A(net1014),
    .B(_2840_),
    .Y(_1539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3978_ (.B1(net1181),
    .VDD(VPWR),
    .Y(_1540_),
    .VSS(VGND),
    .A1(_1479_),
    .A2(_1539_));
 sg13g2_nor2_1 _3979_ (.A(net1384),
    .B(_1482_),
    .Y(_1541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3980_ (.Y(_0152_),
    .B1(_1540_),
    .B2(_1541_),
    .A2(_2836_),
    .A1(net1384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3981_ (.A(net1140),
    .B(net610),
    .X(_1542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3982_ (.B1(net1183),
    .VDD(VPWR),
    .Y(_1543_),
    .VSS(VGND),
    .A1(_1512_),
    .A2(_1542_));
 sg13g2_nor2_1 _3983_ (.A(net1386),
    .B(net374),
    .Y(_1544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3984_ (.Y(_0153_),
    .B1(net611),
    .B2(_1544_),
    .A2(_2835_),
    .A1(net1386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3985_ (.A(net1140),
    .B(\s0.data_out[10][5] ),
    .X(_1545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3986_ (.B1(net1184),
    .VDD(VPWR),
    .Y(_1546_),
    .VSS(VGND),
    .A1(_1505_),
    .A2(_1545_));
 sg13g2_nand3_1 _3987_ (.B(_1509_),
    .C(_1546_),
    .A(net1490),
    .Y(_1547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3988_ (.B1(_1547_),
    .VDD(VPWR),
    .Y(_1548_),
    .VSS(VGND),
    .A1(net1490),
    .A2(net618));
 sg13g2_inv_1 _3989_ (.VDD(VPWR),
    .Y(_0154_),
    .A(_1548_),
    .VSS(VGND));
 sg13g2_nor2_1 _3990_ (.A(net1013),
    .B(_2842_),
    .Y(_1549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3991_ (.B1(net1184),
    .VDD(VPWR),
    .Y(_1550_),
    .VSS(VGND),
    .A1(_1495_),
    .A2(_1549_));
 sg13g2_nand3b_1 _3992_ (.B(_1550_),
    .C(net1491),
    .Y(_1551_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1498_));
 sg13g2_o21ai_1 _3993_ (.B1(_1551_),
    .VDD(VPWR),
    .Y(_1552_),
    .VSS(VGND),
    .A1(net1491),
    .A2(net697));
 sg13g2_inv_1 _3994_ (.VDD(VPWR),
    .Y(_0155_),
    .A(_1552_),
    .VSS(VGND));
 sg13g2_nor2_1 _3995_ (.A(_2746_),
    .B(_2841_),
    .Y(_1553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3996_ (.B1(net1184),
    .VDD(VPWR),
    .Y(_1554_),
    .VSS(VGND),
    .A1(_1488_),
    .A2(_1553_));
 sg13g2_nor2_1 _3997_ (.A(net1387),
    .B(_1491_),
    .Y(_1555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3998_ (.Y(_0156_),
    .B1(_1554_),
    .B2(_1555_),
    .A2(_2834_),
    .A1(net1387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3999_ (.B1(net1137),
    .VDD(VPWR),
    .Y(_1556_),
    .VSS(VGND),
    .A1(net1396),
    .A2(net1129));
 sg13g2_nor2_1 _4000_ (.A(net1396),
    .B(_2747_),
    .Y(_1557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4001_ (.A(_1556_),
    .B(_1557_),
    .Y(_1558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4002_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1013),
    .A2(_1446_),
    .Y(_1559_),
    .B1(_1558_));
 sg13g2_o21ai_1 _4003_ (.B1(_1558_),
    .VDD(VPWR),
    .Y(_1560_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[9] [0]),
    .A2(net1134));
 sg13g2_nor2_1 _4004_ (.A(net1129),
    .B(_1556_),
    .Y(_1561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4005_ (.B1(net1014),
    .VDD(VPWR),
    .Y(_1562_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[9] [0]),
    .A2(net1174));
 sg13g2_nand2_1 _4006_ (.Y(_1563_),
    .A(_1560_),
    .B(_1562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4007_ (.B1(net1491),
    .VDD(VPWR),
    .Y(_1564_),
    .VSS(VGND),
    .A1(_1561_),
    .A2(_1563_));
 sg13g2_a21oi_1 _4008_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2733_),
    .A2(_1559_),
    .Y(_0157_),
    .B1(_1564_));
 sg13g2_and2_1 _4009_ (.A(net1491),
    .B(_1559_),
    .X(_0158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4010_ (.A0(net1170),
    .A1(net1458),
    .S(net1391),
    .X(_0159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4011_ (.A0(net1166),
    .A1(net1450),
    .S(net1390),
    .X(_0160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4012_ (.A(net1390),
    .B(net1162),
    .Y(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4013_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1390),
    .A2(net1334),
    .Y(_0161_),
    .B1(_1565_));
 sg13g2_nand2_1 _4014_ (.Y(_1566_),
    .A(net1391),
    .B(net1435),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4015_ (.B1(_1566_),
    .VDD(VPWR),
    .Y(_0162_),
    .VSS(VGND),
    .A1(net1391),
    .A2(net993));
 sg13g2_nor2_1 _4016_ (.A(net1390),
    .B(net1156),
    .Y(_1567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4017_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1390),
    .A2(_2768_),
    .Y(_0163_),
    .B1(_1567_));
 sg13g2_mux2_1 _4018_ (.A0(net1151),
    .A1(net1416),
    .S(net1390),
    .X(_0164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4019_ (.A0(net1147),
    .A1(net1407),
    .S(net1390),
    .X(_0165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4020_ (.A0(net1142),
    .A1(net1398),
    .S(net1391),
    .X(_0166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4021_ (.Y(_1568_),
    .A(net1131),
    .B(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4022_ (.A0(\s0.data_out[10][1] ),
    .A1(\s0.data_out[9][1] ),
    .S(net1133),
    .X(_1569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4023_ (.A(net1124),
    .B_N(net1168),
    .Y(_1570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4024_ (.A2(_1569_),
    .A1(net1124),
    .B1(_1570_),
    .X(_1571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4025_ (.Y(_1572_),
    .B(\s0.data_out[9][1] ),
    .A_N(net1174),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4026_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1462_),
    .A2(_1572_),
    .Y(_1573_),
    .B1(net1135));
 sg13g2_a21oi_1 _4027_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1136),
    .A2(_1571_),
    .Y(_1574_),
    .B1(_1573_));
 sg13g2_mux2_1 _4028_ (.A0(\s0.data_out[9][0] ),
    .A1(\s0.data_out[10][0] ),
    .S(net1174),
    .X(_1575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4029_ (.Y(_1576_),
    .A(net1014),
    .B(_1575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4030_ (.A(net1124),
    .B_N(net1171),
    .Y(_1577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4031_ (.Y(_1578_),
    .A(net1131),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4032_ (.A0(\s0.data_out[10][0] ),
    .A1(\s0.data_out[9][0] ),
    .S(net1131),
    .X(_1579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4033_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1124),
    .A2(_1579_),
    .Y(_1580_),
    .B1(_1577_));
 sg13g2_nand2b_1 _4034_ (.Y(_1581_),
    .B(net1135),
    .A_N(_1580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4035_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1581_),
    .C1(net1459),
    .B1(_1576_),
    .A1(net1455),
    .Y(_1582_),
    .A2(_1574_));
 sg13g2_nand2_1 _4036_ (.Y(_1583_),
    .A(net1131),
    .B(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4037_ (.A0(\s0.data_out[10][2] ),
    .A1(\s0.data_out[9][2] ),
    .S(net1133),
    .X(_1584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4038_ (.A(net1124),
    .B_N(net1164),
    .Y(_1585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4039_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1124),
    .A2(_1584_),
    .Y(_1586_),
    .B1(_1585_));
 sg13g2_mux2_1 _4040_ (.A0(\s0.data_out[9][2] ),
    .A1(\s0.data_out[10][2] ),
    .S(net1174),
    .X(_1587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4041_ (.Y(_1588_),
    .A(net1014),
    .B(_1587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4042_ (.B1(_1588_),
    .VDD(VPWR),
    .Y(_1589_),
    .VSS(VGND),
    .A1(net1014),
    .A2(_1586_));
 sg13g2_or2_1 _4043_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1590_),
    .B(_1589_),
    .A(net1335));
 sg13g2_xnor2_1 _4044_ (.Y(_1591_),
    .A(net1335),
    .B(_1589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4045_ (.Y(_1592_),
    .A(net1131),
    .B(net589),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4046_ (.A0(\s0.data_out[10][3] ),
    .A1(\s0.data_out[9][3] ),
    .S(net1133),
    .X(_1593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4047_ (.A(net1130),
    .B_N(\s0.data_new_delayed[3] ),
    .Y(_1594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4048_ (.A2(_1593_),
    .A1(net1130),
    .B1(_1594_),
    .X(_1595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4049_ (.Y(_1596_),
    .B(\s0.data_out[9][3] ),
    .A_N(net1177),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4050_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1477_),
    .A2(_1596_),
    .Y(_1597_),
    .B1(net1137));
 sg13g2_a21oi_1 _4051_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1137),
    .A2(_1595_),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_nor2_1 _4052_ (.A(net1441),
    .B(_1598_),
    .Y(_1599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4053_ (.A(net1455),
    .B(_1574_),
    .Y(_1600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _4054_ (.A(_1582_),
    .B(_1591_),
    .C(_1599_),
    .D(_1600_),
    .Y(_1601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4055_ (.Y(_1602_),
    .A(net1442),
    .B(_1598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4056_ (.B1(_1602_),
    .VDD(VPWR),
    .Y(_1603_),
    .VSS(VGND),
    .A1(_1590_),
    .A2(_1599_));
 sg13g2_nor2_1 _4057_ (.A(_1601_),
    .B(_1603_),
    .Y(_1604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4058_ (.Y(_1605_),
    .A(net1132),
    .B(\s0.data_out[9][7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4059_ (.A0(\s0.data_out[10][7] ),
    .A1(\s0.data_out[9][7] ),
    .S(net1134),
    .X(_1606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4060_ (.A(net1128),
    .B_N(net1144),
    .Y(_1607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4061_ (.A2(_1606_),
    .A1(net1128),
    .B1(_1607_),
    .X(_1608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4062_ (.Y(_1609_),
    .B(net505),
    .A_N(net1175),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4063_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1486_),
    .A2(_1609_),
    .Y(_1610_),
    .B1(net1138));
 sg13g2_a21oi_1 _4064_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1139),
    .A2(_1608_),
    .Y(_1611_),
    .B1(_1610_));
 sg13g2_nand2_1 _4065_ (.Y(_1612_),
    .A(net1132),
    .B(net509),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4066_ (.A0(\s0.data_out[10][6] ),
    .A1(\s0.data_out[9][6] ),
    .S(net1134),
    .X(_1613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4067_ (.A(net1129),
    .B_N(net1149),
    .Y(_1614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4068_ (.A2(_1613_),
    .A1(net1128),
    .B1(_1614_),
    .X(_1615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4069_ (.Y(_1616_),
    .B(net509),
    .A_N(net1175),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4070_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1493_),
    .A2(_1616_),
    .Y(_1617_),
    .B1(net1138));
 sg13g2_a21oi_1 _4071_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1139),
    .A2(_1615_),
    .Y(_1618_),
    .B1(_1617_));
 sg13g2_a22oi_1 _4072_ (.Y(_1619_),
    .B1(_1618_),
    .B2(net1414),
    .A2(_1611_),
    .A1(net1405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4073_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1620_),
    .B(_1618_),
    .A(net1414));
 sg13g2_nor2_1 _4074_ (.A(net1405),
    .B(_1611_),
    .Y(_1621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _4075_ (.B(_1619_),
    .C(_1620_),
    .Y(_1622_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1621_));
 sg13g2_nor2b_1 _4076_ (.A(net1130),
    .B_N(net1159),
    .Y(_1623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4077_ (.Y(_1624_),
    .A(net1132),
    .B(\s0.data_out[9][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4078_ (.A0(\s0.data_out[10][4] ),
    .A1(\s0.data_out[9][4] ),
    .S(net1134),
    .X(_1625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4079_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1130),
    .A2(_1625_),
    .Y(_1626_),
    .B1(_1623_));
 sg13g2_nand2b_1 _4080_ (.Y(_1627_),
    .B(net1141),
    .A_N(_1626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4081_ (.A0(\s0.data_out[9][4] ),
    .A1(\s0.data_out[10][4] ),
    .S(net1175),
    .X(_1628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4082_ (.Y(_1629_),
    .A(net1013),
    .B(_1628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4083_ (.B(_1627_),
    .C(_1629_),
    .A(net1433),
    .Y(_1630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4084_ (.Y(_1631_),
    .A(net1132),
    .B(\s0.data_out[9][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4085_ (.A0(\s0.data_out[10][5] ),
    .A1(\s0.data_out[9][5] ),
    .S(net1134),
    .X(_1632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4086_ (.A(net1128),
    .B_N(net1153),
    .Y(_1633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4087_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1128),
    .A2(_1632_),
    .Y(_1634_),
    .B1(_1633_));
 sg13g2_nand2b_1 _4088_ (.Y(_1635_),
    .B(net1138),
    .A_N(_1634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4089_ (.A0(\s0.data_out[9][5] ),
    .A1(\s0.data_out[10][5] ),
    .S(net1175),
    .X(_1636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4090_ (.Y(_1637_),
    .A(net1013),
    .B(_1636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4091_ (.B(_1635_),
    .C(_1637_),
    .A(net1424),
    .Y(_1638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4092_ (.Y(_1639_),
    .A(_1630_),
    .B(_1638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4093_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1627_),
    .A2(_1629_),
    .Y(_1640_),
    .B1(net1433));
 sg13g2_a21oi_1 _4094_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1635_),
    .A2(_1637_),
    .Y(_1641_),
    .B1(net1424));
 sg13g2_or2_1 _4095_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1642_),
    .B(_1641_),
    .A(_1640_));
 sg13g2_or4_1 _4096_ (.A(_1604_),
    .B(_1622_),
    .C(_1639_),
    .D(_1642_),
    .X(_1643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4097_ (.B1(_1638_),
    .VDD(VPWR),
    .Y(_1644_),
    .VSS(VGND),
    .A1(_1630_),
    .A2(_1641_));
 sg13g2_nor2b_1 _4098_ (.A(_1622_),
    .B_N(_1644_),
    .Y(_1645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4099_ (.B1(_1559_),
    .VDD(VPWR),
    .Y(_1646_),
    .VSS(VGND),
    .A1(_1619_),
    .A2(_1621_));
 sg13g2_nor2_1 _4100_ (.A(_1645_),
    .B(_1646_),
    .Y(_1647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4101_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1648_),
    .B(net1331),
    .A(net329));
 sg13g2_a21oi_1 _4102_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1643_),
    .A2(_1647_),
    .Y(_0167_),
    .B1(_1648_));
 sg13g2_and2_1 _4103_ (.A(net1123),
    .B(\s0.data_out[9][0] ),
    .X(_1649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4104_ (.B1(net1135),
    .VDD(VPWR),
    .Y(_1650_),
    .VSS(VGND),
    .A1(_1577_),
    .A2(_1649_));
 sg13g2_nand3_1 _4105_ (.B(_1576_),
    .C(_1650_),
    .A(net1488),
    .Y(_1651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4106_ (.B1(_1651_),
    .VDD(VPWR),
    .Y(_1652_),
    .VSS(VGND),
    .A1(net1488),
    .A2(net626));
 sg13g2_inv_1 _4107_ (.VDD(VPWR),
    .Y(_0168_),
    .A(_1652_),
    .VSS(VGND));
 sg13g2_and2_1 _4108_ (.A(net1124),
    .B(\s0.data_out[9][1] ),
    .X(_1653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4109_ (.B1(net1135),
    .VDD(VPWR),
    .Y(_1654_),
    .VSS(VGND),
    .A1(_1570_),
    .A2(_1653_));
 sg13g2_nor2_1 _4110_ (.A(net1385),
    .B(_1573_),
    .Y(_1655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4111_ (.Y(_0169_),
    .B1(_1654_),
    .B2(_1655_),
    .A2(_2839_),
    .A1(net1385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4112_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1124),
    .A2(net465),
    .Y(_1656_),
    .B1(_1585_));
 sg13g2_a21oi_1 _4113_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1014),
    .A2(_1587_),
    .Y(_1657_),
    .B1(net1385));
 sg13g2_o21ai_1 _4114_ (.B1(_1657_),
    .VDD(VPWR),
    .Y(_1658_),
    .VSS(VGND),
    .A1(net1014),
    .A2(_1656_));
 sg13g2_o21ai_1 _4115_ (.B1(_1658_),
    .VDD(VPWR),
    .Y(_1659_),
    .VSS(VGND),
    .A1(net1488),
    .A2(net674));
 sg13g2_inv_1 _4116_ (.VDD(VPWR),
    .Y(_0170_),
    .A(_1659_),
    .VSS(VGND));
 sg13g2_and2_1 _4117_ (.A(net1127),
    .B(\s0.data_out[9][3] ),
    .X(_1660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4118_ (.B1(net1137),
    .VDD(VPWR),
    .Y(_1661_),
    .VSS(VGND),
    .A1(_1594_),
    .A2(_1660_));
 sg13g2_nor2_1 _4119_ (.A(net1384),
    .B(_1597_),
    .Y(_1662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4120_ (.Y(_0171_),
    .B1(_1661_),
    .B2(_1662_),
    .A2(_2840_),
    .A1(net1388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4121_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1130),
    .A2(net675),
    .Y(_1663_),
    .B1(_1623_));
 sg13g2_a21oi_1 _4122_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1013),
    .A2(_1628_),
    .Y(_1664_),
    .B1(net1387));
 sg13g2_o21ai_1 _4123_ (.B1(_1664_),
    .VDD(VPWR),
    .Y(_1665_),
    .VSS(VGND),
    .A1(net1013),
    .A2(_1663_));
 sg13g2_o21ai_1 _4124_ (.B1(_1665_),
    .VDD(VPWR),
    .Y(_1666_),
    .VSS(VGND),
    .A1(net1490),
    .A2(net610));
 sg13g2_inv_1 _4125_ (.VDD(VPWR),
    .Y(_0172_),
    .A(_1666_),
    .VSS(VGND));
 sg13g2_a21oi_1 _4126_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1128),
    .A2(\s0.data_out[9][5] ),
    .Y(_1667_),
    .B1(_1633_));
 sg13g2_a21oi_1 _4127_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1013),
    .A2(_1636_),
    .Y(_1668_),
    .B1(net1387));
 sg13g2_o21ai_1 _4128_ (.B1(_1668_),
    .VDD(VPWR),
    .Y(_1669_),
    .VSS(VGND),
    .A1(net1013),
    .A2(_1667_));
 sg13g2_o21ai_1 _4129_ (.B1(_1669_),
    .VDD(VPWR),
    .Y(_1670_),
    .VSS(VGND),
    .A1(net1491),
    .A2(net613));
 sg13g2_inv_1 _4130_ (.VDD(VPWR),
    .Y(_0173_),
    .A(net614),
    .VSS(VGND));
 sg13g2_and2_1 _4131_ (.A(net1128),
    .B(net509),
    .X(_1671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4132_ (.B1(net1139),
    .VDD(VPWR),
    .Y(_1672_),
    .VSS(VGND),
    .A1(_1614_),
    .A2(_1671_));
 sg13g2_nor2_1 _4133_ (.A(net1386),
    .B(_1617_),
    .Y(_1673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4134_ (.Y(_0174_),
    .B1(_1672_),
    .B2(_1673_),
    .A2(_2842_),
    .A1(net1386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4135_ (.A(net1128),
    .B(net505),
    .X(_1674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4136_ (.B1(net1139),
    .VDD(VPWR),
    .Y(_1675_),
    .VSS(VGND),
    .A1(_1607_),
    .A2(_1674_));
 sg13g2_nor2_1 _4137_ (.A(net1386),
    .B(_1610_),
    .Y(_1676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4138_ (.Y(_0175_),
    .B1(_1675_),
    .B2(_1676_),
    .A2(_2841_),
    .A1(net1387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4139_ (.B1(net1126),
    .VDD(VPWR),
    .Y(_1677_),
    .VSS(VGND),
    .A1(net1396),
    .A2(net1117));
 sg13g2_nand2_1 _4140_ (.Y(_1678_),
    .A(net1338),
    .B(net1121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4141_ (.Y(_1679_),
    .B(_1678_),
    .A_N(_1677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4142_ (.B1(_1679_),
    .VDD(VPWR),
    .Y(_1680_),
    .VSS(VGND),
    .A1(net1126),
    .A2(_1557_));
 sg13g2_nor2_1 _4143_ (.A(net358),
    .B(net1121),
    .Y(_1681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4144_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1682_),
    .B(_1681_),
    .A(_1679_));
 sg13g2_nor2_1 _4145_ (.A(net1116),
    .B(_1677_),
    .Y(_1683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4146_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2732_),
    .A2(_2747_),
    .Y(_1684_),
    .B1(net1125));
 sg13g2_nor2_1 _4147_ (.A(_1683_),
    .B(_1684_),
    .Y(_1685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4148_ (.B1(net1488),
    .VDD(VPWR),
    .Y(_1686_),
    .VSS(VGND),
    .A1(net666),
    .A2(_1680_));
 sg13g2_a21oi_1 _4149_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1682_),
    .A2(_1685_),
    .Y(_0176_),
    .B1(_1686_));
 sg13g2_nor2_1 _4150_ (.A(net1384),
    .B(_1680_),
    .Y(_0177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4151_ (.A(net1482),
    .B(net324),
    .X(_0178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4152_ (.Y(_1687_),
    .A(net1118),
    .B(net518),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4153_ (.A0(\s0.data_out[9][2] ),
    .A1(\s0.data_out[8][2] ),
    .S(net1119),
    .X(_1688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4154_ (.A(net1113),
    .B_N(net1164),
    .Y(_1689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4155_ (.A2(_1688_),
    .A1(net1113),
    .B1(_1689_),
    .X(_1690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4156_ (.Y(_1691_),
    .B(\s0.data_out[8][2] ),
    .A_N(net1131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4157_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1583_),
    .A2(_1691_),
    .Y(_1692_),
    .B1(net1122));
 sg13g2_a21oi_1 _4158_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1122),
    .A2(_1690_),
    .Y(_1693_),
    .B1(_1692_));
 sg13g2_or2_1 _4159_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1694_),
    .B(_1693_),
    .A(net1446));
 sg13g2_nor2b_1 _4160_ (.A(net1111),
    .B_N(net1168),
    .Y(_1695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4161_ (.Y(_1696_),
    .A(net1118),
    .B(net673),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4162_ (.B1(_1696_),
    .VDD(VPWR),
    .Y(_1697_),
    .VSS(VGND),
    .A1(net1118),
    .A2(_2843_));
 sg13g2_a21o_1 _4163_ (.A2(_1697_),
    .A1(net1111),
    .B1(_1695_),
    .X(_1698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4164_ (.Y(_1699_),
    .A(_2747_),
    .B(\s0.data_out[8][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4165_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1568_),
    .A2(_1699_),
    .Y(_1700_),
    .B1(net1122));
 sg13g2_a21oi_1 _4166_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1122),
    .A2(_1698_),
    .Y(_1701_),
    .B1(_1700_));
 sg13g2_mux2_1 _4167_ (.A0(\s0.data_out[9][0] ),
    .A1(\s0.data_out[8][0] ),
    .S(net1118),
    .X(_1702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4168_ (.A(net1111),
    .B_N(net1171),
    .Y(_1703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4169_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1111),
    .A2(_1702_),
    .Y(_1704_),
    .B1(_1703_));
 sg13g2_nand2b_1 _4170_ (.Y(_1705_),
    .B(net1122),
    .A_N(_1704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4171_ (.B1(_1578_),
    .VDD(VPWR),
    .Y(_1706_),
    .VSS(VGND),
    .A1(net1131),
    .A2(_2854_));
 sg13g2_nand2b_1 _4172_ (.Y(_1707_),
    .B(_1706_),
    .A_N(net1122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4173_ (.B1(_1694_),
    .VDD(VPWR),
    .Y(_1708_),
    .VSS(VGND),
    .A1(net1455),
    .A2(_1701_));
 sg13g2_a221oi_1 _4174_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1707_),
    .C1(net1459),
    .B1(_1705_),
    .A1(net1455),
    .Y(_1709_),
    .A2(_1701_));
 sg13g2_nand2_1 _4175_ (.Y(_1710_),
    .A(net1119),
    .B(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4176_ (.B1(_1710_),
    .VDD(VPWR),
    .Y(_1711_),
    .VSS(VGND),
    .A1(net1119),
    .A2(_2844_));
 sg13g2_nor2_1 _4177_ (.A(net1112),
    .B(net994),
    .Y(_1712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4178_ (.A2(_1711_),
    .A1(net1113),
    .B1(_1712_),
    .X(_1713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4179_ (.Y(_1714_),
    .A(_2747_),
    .B(\s0.data_out[8][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4180_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1592_),
    .A2(_1714_),
    .Y(_1715_),
    .B1(net1123));
 sg13g2_a21oi_1 _4181_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1123),
    .A2(_1713_),
    .Y(_1716_),
    .B1(_1715_));
 sg13g2_a22oi_1 _4182_ (.Y(_1717_),
    .B1(_1716_),
    .B2(net1442),
    .A2(_1693_),
    .A1(net1446),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4183_ (.B1(_1717_),
    .VDD(VPWR),
    .Y(_1718_),
    .VSS(VGND),
    .A1(_1708_),
    .A2(_1709_));
 sg13g2_nand2_1 _4184_ (.Y(_1719_),
    .A(net1120),
    .B(net654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4185_ (.A0(\s0.data_out[9][6] ),
    .A1(\s0.data_out[8][6] ),
    .S(net1121),
    .X(_1720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4186_ (.A(net1116),
    .B_N(net1149),
    .Y(_1721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4187_ (.A2(_1720_),
    .A1(net1116),
    .B1(_1721_),
    .X(_1722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4188_ (.Y(_1723_),
    .B(\s0.data_out[8][6] ),
    .A_N(net1132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4189_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1612_),
    .A2(_1723_),
    .Y(_1724_),
    .B1(net1126));
 sg13g2_a21oi_1 _4190_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1126),
    .A2(_1722_),
    .Y(_1725_),
    .B1(_1724_));
 sg13g2_nand2_1 _4191_ (.Y(_1726_),
    .A(net1120),
    .B(net371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4192_ (.A0(\s0.data_out[9][7] ),
    .A1(\s0.data_out[8][7] ),
    .S(net1121),
    .X(_1727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4193_ (.A(net1116),
    .B_N(net1145),
    .Y(_1728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4194_ (.A2(_1727_),
    .A1(net1117),
    .B1(_1728_),
    .X(_1729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4195_ (.Y(_1730_),
    .B(net371),
    .A_N(net1132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4196_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1605_),
    .A2(_1730_),
    .Y(_1731_),
    .B1(net1126));
 sg13g2_a21oi_1 _4197_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1126),
    .A2(_1729_),
    .Y(_1732_),
    .B1(_1731_));
 sg13g2_a22oi_1 _4198_ (.Y(_1733_),
    .B1(_1732_),
    .B2(net1405),
    .A2(_1725_),
    .A1(net1414),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4199_ (.A(net1414),
    .B(_1725_),
    .Y(_1734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4200_ (.A(net1405),
    .B(_1732_),
    .Y(_1735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4201_ (.A(_1734_),
    .B(_1735_),
    .Y(_1736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4202_ (.Y(_1737_),
    .A(net1120),
    .B(net687),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4203_ (.A0(\s0.data_out[9][5] ),
    .A1(\s0.data_out[8][5] ),
    .S(net1121),
    .X(_1738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4204_ (.A(net1116),
    .B_N(net1154),
    .Y(_1739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4205_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1116),
    .A2(_1738_),
    .Y(_1740_),
    .B1(_1739_));
 sg13g2_nand2b_1 _4206_ (.Y(_1741_),
    .B(net1125),
    .A_N(_1740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4207_ (.B1(_1631_),
    .VDD(VPWR),
    .Y(_1742_),
    .VSS(VGND),
    .A1(net1132),
    .A2(_2849_));
 sg13g2_nand2b_1 _4208_ (.Y(_1743_),
    .B(_1742_),
    .A_N(net1125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4209_ (.B(_1741_),
    .C(_1743_),
    .A(net1424),
    .Y(_1744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4210_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1741_),
    .A2(_1743_),
    .Y(_1745_),
    .B1(net1424));
 sg13g2_nand2_1 _4211_ (.Y(_1746_),
    .A(net1120),
    .B(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4212_ (.A0(\s0.data_out[9][4] ),
    .A1(\s0.data_out[8][4] ),
    .S(net1121),
    .X(_1747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4213_ (.A(net1116),
    .B_N(net1159),
    .Y(_1748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4214_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1116),
    .A2(_1747_),
    .Y(_1749_),
    .B1(_1748_));
 sg13g2_nand2b_1 _4215_ (.Y(_1750_),
    .B(net1125),
    .A_N(_1749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4216_ (.B1(_1624_),
    .VDD(VPWR),
    .Y(_1751_),
    .VSS(VGND),
    .A1(net1132),
    .A2(_2850_));
 sg13g2_nand2b_1 _4217_ (.Y(_1752_),
    .B(_1751_),
    .A_N(net1125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4218_ (.B(_1750_),
    .C(_1752_),
    .A(net1433),
    .Y(_1753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4219_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1750_),
    .A2(_1752_),
    .Y(_1754_),
    .B1(net1433));
 sg13g2_o21ai_1 _4220_ (.B1(_1744_),
    .VDD(VPWR),
    .Y(_1755_),
    .VSS(VGND),
    .A1(net1442),
    .A2(_1716_));
 sg13g2_nand2b_1 _4221_ (.Y(_1756_),
    .B(_1753_),
    .A_N(_1745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4222_ (.A(_1754_),
    .B(_1755_),
    .C(_1756_),
    .Y(_1757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4223_ (.B(_1733_),
    .C(_1736_),
    .A(_1718_),
    .Y(_1758_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1757_));
 sg13g2_o21ai_1 _4224_ (.B1(_1744_),
    .VDD(VPWR),
    .Y(_1759_),
    .VSS(VGND),
    .A1(_1745_),
    .A2(_1753_));
 sg13g2_and3_1 _4225_ (.X(_1760_),
    .A(_1733_),
    .B(_1736_),
    .C(_1759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4226_ (.A(_1733_),
    .B(_1735_),
    .Y(_1761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4227_ (.A(_1680_),
    .B(_1760_),
    .C(_1761_),
    .Y(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4228_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1763_),
    .B(net1332),
    .A(net336));
 sg13g2_a21oi_1 _4229_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1758_),
    .A2(_1762_),
    .Y(_0179_),
    .B1(_1763_));
 sg13g2_nor2_1 _4230_ (.A(net1000),
    .B(_2854_),
    .Y(_1764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4231_ (.B1(net1122),
    .VDD(VPWR),
    .Y(_1765_),
    .VSS(VGND),
    .A1(_1703_),
    .A2(_1764_));
 sg13g2_nand3_1 _4232_ (.B(_1707_),
    .C(_1765_),
    .A(net1481),
    .Y(_1766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4233_ (.B1(_1766_),
    .VDD(VPWR),
    .Y(_1767_),
    .VSS(VGND),
    .A1(net1481),
    .A2(net596));
 sg13g2_inv_1 _4234_ (.VDD(VPWR),
    .Y(_0180_),
    .A(_1767_),
    .VSS(VGND));
 sg13g2_nor2_1 _4235_ (.A(net1000),
    .B(_2853_),
    .Y(_1768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4236_ (.B1(net1122),
    .VDD(VPWR),
    .Y(_1769_),
    .VSS(VGND),
    .A1(_1695_),
    .A2(_1768_));
 sg13g2_nor2_1 _4237_ (.A(net1374),
    .B(_1700_),
    .Y(_1770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4238_ (.Y(_0181_),
    .B1(_1769_),
    .B2(_1770_),
    .A2(_2843_),
    .A1(net1374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4239_ (.A(net1000),
    .B(_2852_),
    .Y(_1771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4240_ (.B1(net1123),
    .VDD(VPWR),
    .Y(_1772_),
    .VSS(VGND),
    .A1(_1689_),
    .A2(_1771_));
 sg13g2_nor2_1 _4241_ (.A(net1376),
    .B(_1692_),
    .Y(_1773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4242_ (.Y(_0182_),
    .B1(_1772_),
    .B2(_1773_),
    .A2(_2845_),
    .A1(net1376),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4243_ (.A(net1000),
    .B(_2851_),
    .Y(_1774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4244_ (.B1(net1123),
    .VDD(VPWR),
    .Y(_1775_),
    .VSS(VGND),
    .A1(_1712_),
    .A2(_1774_));
 sg13g2_nor2_1 _4245_ (.A(net1375),
    .B(_1715_),
    .Y(_1776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4246_ (.Y(_0183_),
    .B1(_1775_),
    .B2(_1776_),
    .A2(_2844_),
    .A1(net1375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4247_ (.A(net1000),
    .B(_2850_),
    .Y(_1777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4248_ (.B1(net1125),
    .VDD(VPWR),
    .Y(_1778_),
    .VSS(VGND),
    .A1(_1748_),
    .A2(_1777_));
 sg13g2_nand3_1 _4249_ (.B(_1752_),
    .C(_1778_),
    .A(net1488),
    .Y(_1779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4250_ (.B1(_1779_),
    .VDD(VPWR),
    .Y(_1780_),
    .VSS(VGND),
    .A1(net1489),
    .A2(net675));
 sg13g2_inv_1 _4251_ (.VDD(VPWR),
    .Y(_0184_),
    .A(_1780_),
    .VSS(VGND));
 sg13g2_nor2_1 _4252_ (.A(net1000),
    .B(_2849_),
    .Y(_1781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4253_ (.B1(net1125),
    .VDD(VPWR),
    .Y(_1782_),
    .VSS(VGND),
    .A1(_1739_),
    .A2(_1781_));
 sg13g2_nand3_1 _4254_ (.B(_1743_),
    .C(_1782_),
    .A(net1489),
    .Y(_1783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4255_ (.B1(_1783_),
    .VDD(VPWR),
    .Y(_1784_),
    .VSS(VGND),
    .A1(net1489),
    .A2(net680));
 sg13g2_inv_1 _4256_ (.VDD(VPWR),
    .Y(_0185_),
    .A(_1784_),
    .VSS(VGND));
 sg13g2_and2_1 _4257_ (.A(net1117),
    .B(\s0.data_out[8][6] ),
    .X(_1785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4258_ (.B1(net1126),
    .VDD(VPWR),
    .Y(_1786_),
    .VSS(VGND),
    .A1(_1721_),
    .A2(_1785_));
 sg13g2_nor2_1 _4259_ (.A(net1384),
    .B(_1724_),
    .Y(_1787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4260_ (.Y(_0186_),
    .B1(_1786_),
    .B2(_1787_),
    .A2(_2847_),
    .A1(net1384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4261_ (.A(net1000),
    .B(_2848_),
    .Y(_1788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4262_ (.B1(net1125),
    .VDD(VPWR),
    .Y(_1789_),
    .VSS(VGND),
    .A1(_1728_),
    .A2(_1788_));
 sg13g2_nor2_1 _4263_ (.A(net1384),
    .B(net372),
    .Y(_1790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4264_ (.Y(_0187_),
    .B1(_1789_),
    .B2(_1790_),
    .A2(_2846_),
    .A1(net1384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4265_ (.B1(net1114),
    .VDD(VPWR),
    .Y(_1791_),
    .VSS(VGND),
    .A1(net1394),
    .A2(net1103));
 sg13g2_nor2_1 _4266_ (.A(net1394),
    .B(_2760_),
    .Y(_1792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4267_ (.A(_1791_),
    .B(_1792_),
    .Y(_1793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4268_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2759_),
    .A2(_1678_),
    .Y(_1794_),
    .B1(_1793_));
 sg13g2_o21ai_1 _4269_ (.B1(_1793_),
    .VDD(VPWR),
    .Y(_1795_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[7] [0]),
    .A2(net1107));
 sg13g2_nor2_1 _4270_ (.A(net1103),
    .B(_1791_),
    .Y(_1796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4271_ (.B1(_2759_),
    .VDD(VPWR),
    .Y(_1797_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[7] [0]),
    .A2(net1120));
 sg13g2_nand2_1 _4272_ (.Y(_1798_),
    .A(_1795_),
    .B(_1797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4273_ (.B1(net1481),
    .VDD(VPWR),
    .Y(_1799_),
    .VSS(VGND),
    .A1(_1796_),
    .A2(_1798_));
 sg13g2_a21oi_1 _4274_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2732_),
    .A2(_1794_),
    .Y(_0188_),
    .B1(_1799_));
 sg13g2_and2_1 _4275_ (.A(net1481),
    .B(_1794_),
    .X(_0189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4276_ (.A(net1480),
    .B(net344),
    .X(_0190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4277_ (.Y(_1800_),
    .A(net1105),
    .B(net453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4278_ (.A0(\s0.data_out[8][2] ),
    .A1(\s0.data_out[7][2] ),
    .S(net1105),
    .X(_1801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4279_ (.A(net1098),
    .B_N(net1164),
    .Y(_1802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4280_ (.A2(_1801_),
    .A1(net1099),
    .B1(_1802_),
    .X(_1803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4281_ (.Y(_1804_),
    .B(net453),
    .A_N(net1118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4282_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1687_),
    .A2(_1804_),
    .Y(_1805_),
    .B1(net1110));
 sg13g2_a21oi_1 _4283_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1110),
    .A2(_1803_),
    .Y(_1806_),
    .B1(_1805_));
 sg13g2_or2_1 _4284_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1807_),
    .B(_1806_),
    .A(net1446));
 sg13g2_nand2_1 _4285_ (.Y(_1808_),
    .A(net1105),
    .B(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4286_ (.B1(_1808_),
    .VDD(VPWR),
    .Y(_1809_),
    .VSS(VGND),
    .A1(net1105),
    .A2(_2853_));
 sg13g2_nor2b_1 _4287_ (.A(net1098),
    .B_N(net1168),
    .Y(_1810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4288_ (.A2(_1809_),
    .A1(net1098),
    .B1(_1810_),
    .X(_1811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4289_ (.Y(_1812_),
    .B(net408),
    .A_N(net1118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4290_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1696_),
    .A2(_1812_),
    .Y(_1813_),
    .B1(net1110));
 sg13g2_a21oi_1 _4291_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1110),
    .A2(_1811_),
    .Y(_1814_),
    .B1(_1813_));
 sg13g2_nand2_1 _4292_ (.Y(_1815_),
    .A(net1106),
    .B(\s0.data_out[7][0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4293_ (.B1(_1815_),
    .VDD(VPWR),
    .Y(_1816_),
    .VSS(VGND),
    .A1(net1106),
    .A2(_2854_));
 sg13g2_nor2b_1 _4294_ (.A(net1098),
    .B_N(net1171),
    .Y(_1817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4295_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1098),
    .A2(_1816_),
    .Y(_1818_),
    .B1(_1817_));
 sg13g2_nand2b_1 _4296_ (.Y(_1819_),
    .B(net1110),
    .A_N(_1818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4297_ (.A0(\s0.data_out[7][0] ),
    .A1(\s0.data_out[8][0] ),
    .S(net1118),
    .X(_1820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4298_ (.Y(_1821_),
    .A(net1000),
    .B(_1820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4299_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1821_),
    .C1(net1459),
    .B1(_1819_),
    .A1(net1456),
    .Y(_1822_),
    .A2(_1814_));
 sg13g2_o21ai_1 _4300_ (.B1(_1807_),
    .VDD(VPWR),
    .Y(_1823_),
    .VSS(VGND),
    .A1(net1456),
    .A2(_1814_));
 sg13g2_nand2_1 _4301_ (.Y(_1824_),
    .A(net1106),
    .B(\s0.data_out[7][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4302_ (.B1(_1824_),
    .VDD(VPWR),
    .Y(_1825_),
    .VSS(VGND),
    .A1(net1106),
    .A2(_2851_));
 sg13g2_nor2_1 _4303_ (.A(net1099),
    .B(net994),
    .Y(_1826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4304_ (.A2(_1825_),
    .A1(net1099),
    .B1(_1826_),
    .X(_1827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4305_ (.Y(_1828_),
    .B(net632),
    .A_N(net1118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4306_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1710_),
    .A2(_1828_),
    .Y(_1829_),
    .B1(net1112));
 sg13g2_a21oi_1 _4307_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1112),
    .A2(_1827_),
    .Y(_1830_),
    .B1(_1829_));
 sg13g2_a22oi_1 _4308_ (.Y(_1831_),
    .B1(_1830_),
    .B2(net1441),
    .A2(_1806_),
    .A1(net1446),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4309_ (.B1(_1831_),
    .VDD(VPWR),
    .Y(_1832_),
    .VSS(VGND),
    .A1(_1822_),
    .A2(_1823_));
 sg13g2_nand2_1 _4310_ (.Y(_1833_),
    .A(net1107),
    .B(net627),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4311_ (.A0(\s0.data_out[8][6] ),
    .A1(\s0.data_out[7][6] ),
    .S(net1108),
    .X(_1834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4312_ (.A(net1103),
    .B_N(net1149),
    .Y(_1835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4313_ (.A2(_1834_),
    .A1(net1102),
    .B1(_1835_),
    .X(_1836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4314_ (.Y(_1837_),
    .B(net627),
    .A_N(net1120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4315_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1719_),
    .A2(_1837_),
    .Y(_1838_),
    .B1(net1115));
 sg13g2_a21oi_1 _4316_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1114),
    .A2(_1836_),
    .Y(_1839_),
    .B1(_1838_));
 sg13g2_nand2_1 _4317_ (.Y(_1840_),
    .A(net1107),
    .B(net555),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4318_ (.A0(\s0.data_out[8][7] ),
    .A1(\s0.data_out[7][7] ),
    .S(net1108),
    .X(_1841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4319_ (.A(net1102),
    .B_N(net1144),
    .Y(_1842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4320_ (.A2(_1841_),
    .A1(net1103),
    .B1(_1842_),
    .X(_1843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4321_ (.Y(_1844_),
    .B(net555),
    .A_N(net1120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4322_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1726_),
    .A2(_1844_),
    .Y(_1845_),
    .B1(net1115));
 sg13g2_a21oi_1 _4323_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1115),
    .A2(_1843_),
    .Y(_1846_),
    .B1(_1845_));
 sg13g2_a22oi_1 _4324_ (.Y(_1847_),
    .B1(_1846_),
    .B2(net1403),
    .A2(_1839_),
    .A1(net1412),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4325_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1848_),
    .B(_1839_),
    .A(net1412));
 sg13g2_or2_1 _4326_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1849_),
    .B(_1846_),
    .A(net1403));
 sg13g2_inv_1 _4327_ (.VDD(VPWR),
    .Y(_1850_),
    .A(_1849_),
    .VSS(VGND));
 sg13g2_and3_1 _4328_ (.X(_1851_),
    .A(_1847_),
    .B(_1848_),
    .C(_1849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4329_ (.B(_1848_),
    .C(_1849_),
    .A(_1847_),
    .Y(_1852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4330_ (.Y(_1853_),
    .A(net1107),
    .B(net470),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4331_ (.A0(\s0.data_out[8][5] ),
    .A1(\s0.data_out[7][5] ),
    .S(net1108),
    .X(_1854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4332_ (.A(net1102),
    .B_N(net1153),
    .Y(_1855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4333_ (.A2(_1854_),
    .A1(net1102),
    .B1(_1855_),
    .X(_1856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4334_ (.Y(_1857_),
    .B(net470),
    .A_N(net1120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4335_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1737_),
    .A2(_1857_),
    .Y(_1858_),
    .B1(net1114));
 sg13g2_a21oi_1 _4336_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1114),
    .A2(_1856_),
    .Y(_1859_),
    .B1(_1858_));
 sg13g2_nand2_1 _4337_ (.Y(_1860_),
    .A(net1422),
    .B(_1859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4338_ (.A0(\s0.data_out[8][4] ),
    .A1(\s0.data_out[7][4] ),
    .S(net1108),
    .X(_1861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4339_ (.A(net1102),
    .B_N(net1158),
    .Y(_1862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4340_ (.A2(_1861_),
    .A1(net1102),
    .B1(_1862_),
    .X(_1863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4341_ (.Y(_1864_),
    .B(net639),
    .A_N(net1119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4342_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1746_),
    .A2(_1864_),
    .Y(_1865_),
    .B1(net1114));
 sg13g2_a21oi_1 _4343_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1114),
    .A2(_1863_),
    .Y(_1866_),
    .B1(_1865_));
 sg13g2_nand2_1 _4344_ (.Y(_1867_),
    .A(net1431),
    .B(_1866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4345_ (.A(net1422),
    .B(_1859_),
    .Y(_1868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4346_ (.B1(_1860_),
    .VDD(VPWR),
    .Y(_1869_),
    .VSS(VGND),
    .A1(net1431),
    .A2(_1866_));
 sg13g2_o21ai_1 _4347_ (.B1(_1867_),
    .VDD(VPWR),
    .Y(_1870_),
    .VSS(VGND),
    .A1(net1441),
    .A2(_1830_));
 sg13g2_nor4_1 _4348_ (.A(_1852_),
    .B(_1868_),
    .C(_1869_),
    .D(_1870_),
    .Y(_1871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4349_ (.B1(_1860_),
    .VDD(VPWR),
    .Y(_1872_),
    .VSS(VGND),
    .A1(_1867_),
    .A2(_1868_));
 sg13g2_o21ai_1 _4350_ (.B1(_1794_),
    .VDD(VPWR),
    .Y(_1873_),
    .VSS(VGND),
    .A1(_1847_),
    .A2(_1850_));
 sg13g2_a221oi_1 _4351_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1851_),
    .C1(_1873_),
    .B1(_1872_),
    .A1(_1832_),
    .Y(_1874_),
    .A2(_1871_));
 sg13g2_nor3_1 _4352_ (.A(net324),
    .B(net1331),
    .C(_1874_),
    .Y(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4353_ (.A(net1098),
    .B(\s0.data_out[7][0] ),
    .X(_1875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4354_ (.B1(net1110),
    .VDD(VPWR),
    .Y(_1876_),
    .VSS(VGND),
    .A1(_1817_),
    .A2(_1875_));
 sg13g2_nand3_1 _4355_ (.B(_1821_),
    .C(_1876_),
    .A(net1481),
    .Y(_1877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4356_ (.B1(_1877_),
    .VDD(VPWR),
    .Y(_1878_),
    .VSS(VGND),
    .A1(net1481),
    .A2(net537));
 sg13g2_inv_1 _4357_ (.VDD(VPWR),
    .Y(_0192_),
    .A(net538),
    .VSS(VGND));
 sg13g2_and2_1 _4358_ (.A(net1098),
    .B(net408),
    .X(_1879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4359_ (.B1(net1110),
    .VDD(VPWR),
    .Y(_1880_),
    .VSS(VGND),
    .A1(_1810_),
    .A2(_1879_));
 sg13g2_nor2_1 _4360_ (.A(net1374),
    .B(_1813_),
    .Y(_1881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4361_ (.Y(_0193_),
    .B1(_1880_),
    .B2(_1881_),
    .A2(_2853_),
    .A1(net1374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4362_ (.A(net1098),
    .B(net453),
    .X(_1882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4363_ (.B1(net1110),
    .VDD(VPWR),
    .Y(_1883_),
    .VSS(VGND),
    .A1(_1802_),
    .A2(_1882_));
 sg13g2_nor2_1 _4364_ (.A(net1374),
    .B(_1805_),
    .Y(_1884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4365_ (.Y(_0194_),
    .B1(_1883_),
    .B2(_1884_),
    .A2(_2852_),
    .A1(net1374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4366_ (.A(net1099),
    .B(net632),
    .X(_1885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4367_ (.B1(net1112),
    .VDD(VPWR),
    .Y(_1886_),
    .VSS(VGND),
    .A1(_1826_),
    .A2(_1885_));
 sg13g2_nor2_1 _4368_ (.A(net1374),
    .B(_1829_),
    .Y(_1887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4369_ (.Y(_0195_),
    .B1(_1886_),
    .B2(_1887_),
    .A2(_2851_),
    .A1(net1374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4370_ (.A(net1102),
    .B(net639),
    .X(_1888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4371_ (.B1(net1114),
    .VDD(VPWR),
    .Y(_1889_),
    .VSS(VGND),
    .A1(_1862_),
    .A2(_1888_));
 sg13g2_nor2_1 _4372_ (.A(net1376),
    .B(_1865_),
    .Y(_1890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4373_ (.Y(_0196_),
    .B1(_1889_),
    .B2(_1890_),
    .A2(_2850_),
    .A1(net1375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4374_ (.A(net1102),
    .B(net470),
    .X(_1891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4375_ (.B1(net1114),
    .VDD(VPWR),
    .Y(_1892_),
    .VSS(VGND),
    .A1(_1855_),
    .A2(_1891_));
 sg13g2_nor2_1 _4376_ (.A(net1375),
    .B(_1858_),
    .Y(_1893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4377_ (.Y(_0197_),
    .B1(_1892_),
    .B2(_1893_),
    .A2(_2849_),
    .A1(net1375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4378_ (.A(net1103),
    .B(\s0.data_out[7][6] ),
    .X(_1894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4379_ (.B1(net1115),
    .VDD(VPWR),
    .Y(_1895_),
    .VSS(VGND),
    .A1(_1835_),
    .A2(_1894_));
 sg13g2_nand3b_1 _4380_ (.B(_1895_),
    .C(net1481),
    .Y(_1896_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1838_));
 sg13g2_o21ai_1 _4381_ (.B1(_1896_),
    .VDD(VPWR),
    .Y(_1897_),
    .VSS(VGND),
    .A1(net1481),
    .A2(net654));
 sg13g2_inv_1 _4382_ (.VDD(VPWR),
    .Y(_0198_),
    .A(net655),
    .VSS(VGND));
 sg13g2_and2_1 _4383_ (.A(net1103),
    .B(net555),
    .X(_1898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4384_ (.B1(net1115),
    .VDD(VPWR),
    .Y(_1899_),
    .VSS(VGND),
    .A1(_1842_),
    .A2(_1898_));
 sg13g2_nor2_1 _4385_ (.A(net1375),
    .B(_1845_),
    .Y(_1900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4386_ (.Y(_0199_),
    .B1(net556),
    .B2(_1900_),
    .A2(_2848_),
    .A1(net1375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4387_ (.B1(net1100),
    .VDD(VPWR),
    .Y(_1901_),
    .VSS(VGND),
    .A1(net1394),
    .A2(net1089));
 sg13g2_nand2_1 _4388_ (.Y(_1902_),
    .A(net1337),
    .B(net1094),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4389_ (.Y(_1903_),
    .B(_1902_),
    .A_N(_1901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4390_ (.B1(_1903_),
    .VDD(VPWR),
    .Y(_1904_),
    .VSS(VGND),
    .A1(net1101),
    .A2(_1792_));
 sg13g2_nor2_1 _4391_ (.A(net364),
    .B(net1094),
    .Y(_1905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4392_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1906_),
    .B(_1905_),
    .A(_1903_));
 sg13g2_nor2_1 _4393_ (.A(net1089),
    .B(_1901_),
    .Y(_1907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4394_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2731_),
    .A2(_2760_),
    .Y(_1908_),
    .B1(net1100));
 sg13g2_nor2_1 _4395_ (.A(_1907_),
    .B(_1908_),
    .Y(_1909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4396_ (.B1(net1482),
    .VDD(VPWR),
    .Y(_1910_),
    .VSS(VGND),
    .A1(net552),
    .A2(_1904_));
 sg13g2_a21oi_1 _4397_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1906_),
    .A2(_1909_),
    .Y(_0200_),
    .B1(_1910_));
 sg13g2_nor2_1 _4398_ (.A(net1375),
    .B(_1904_),
    .Y(_0201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4399_ (.A(net1475),
    .B(net339),
    .X(_0202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4400_ (.A0(\s0.data_out[7][2] ),
    .A1(\s0.data_out[6][2] ),
    .S(net1092),
    .X(_1911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4401_ (.A(net1085),
    .B_N(net1165),
    .Y(_1912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4402_ (.A2(_1911_),
    .A1(net1086),
    .B1(_1912_),
    .X(_1913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4403_ (.Y(_1914_),
    .B(\s0.data_out[6][2] ),
    .A_N(net1105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4404_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1800_),
    .A2(_1914_),
    .Y(_1915_),
    .B1(net1096));
 sg13g2_a21oi_1 _4405_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1097),
    .A2(_1913_),
    .Y(_1916_),
    .B1(_1915_));
 sg13g2_nor2_1 _4406_ (.A(net1447),
    .B(_1916_),
    .Y(_1917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4407_ (.Y(_1918_),
    .A(net1092),
    .B(net501),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4408_ (.A0(\s0.data_out[7][1] ),
    .A1(\s0.data_out[6][1] ),
    .S(net1092),
    .X(_1919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4409_ (.A(net1085),
    .B_N(net1169),
    .Y(_1920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4410_ (.A2(_1919_),
    .A1(net1085),
    .B1(_1920_),
    .X(_1921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4411_ (.Y(_1922_),
    .B(\s0.data_out[6][1] ),
    .A_N(net1105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4412_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1808_),
    .A2(_1922_),
    .Y(_1923_),
    .B1(net1096));
 sg13g2_a21oi_1 _4413_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1096),
    .A2(_1921_),
    .Y(_1924_),
    .B1(_1923_));
 sg13g2_mux2_1 _4414_ (.A0(\s0.data_out[7][0] ),
    .A1(\s0.data_out[6][0] ),
    .S(net1092),
    .X(_1925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4415_ (.A(net1086),
    .B_N(net1172),
    .Y(_1926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4416_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1086),
    .A2(_1925_),
    .Y(_1927_),
    .B1(_1926_));
 sg13g2_nand2b_1 _4417_ (.Y(_1928_),
    .B(net1096),
    .A_N(_1927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4418_ (.B1(_1815_),
    .VDD(VPWR),
    .Y(_1929_),
    .VSS(VGND),
    .A1(net1105),
    .A2(_2864_));
 sg13g2_nand2b_1 _4419_ (.Y(_1930_),
    .B(_1929_),
    .A_N(net1096),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4420_ (.A(net1453),
    .B(_1924_),
    .Y(_1931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4421_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1930_),
    .C1(net1460),
    .B1(_1928_),
    .A1(net1453),
    .Y(_1932_),
    .A2(_1924_));
 sg13g2_nor3_1 _4422_ (.A(_1917_),
    .B(_1931_),
    .C(_1932_),
    .Y(_1933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4423_ (.Y(_1934_),
    .A(net1093),
    .B(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4424_ (.B1(_1934_),
    .VDD(VPWR),
    .Y(_1935_),
    .VSS(VGND),
    .A1(net1093),
    .A2(_2857_));
 sg13g2_nor2_1 _4425_ (.A(net1087),
    .B(net994),
    .Y(_1936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4426_ (.A2(_1935_),
    .A1(net1087),
    .B1(_1936_),
    .X(_1937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4427_ (.Y(_1938_),
    .A(_2760_),
    .B(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4428_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1824_),
    .A2(_1938_),
    .Y(_1939_),
    .B1(net1097));
 sg13g2_a21oi_1 _4429_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1097),
    .A2(_1937_),
    .Y(_1940_),
    .B1(_1939_));
 sg13g2_a221oi_1 _4430_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net1442),
    .C1(_1933_),
    .B1(_1940_),
    .A1(net1447),
    .Y(_1941_),
    .A2(_1916_));
 sg13g2_nand2_1 _4431_ (.Y(_1942_),
    .A(net1094),
    .B(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4432_ (.A0(\s0.data_out[7][6] ),
    .A1(\s0.data_out[6][6] ),
    .S(net1094),
    .X(_1943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4433_ (.A(net1089),
    .B_N(net1149),
    .Y(_1944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4434_ (.A2(_1943_),
    .A1(net1089),
    .B1(_1944_),
    .X(_1945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4435_ (.Y(_1946_),
    .B(net578),
    .A_N(net1107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4436_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1833_),
    .A2(_1946_),
    .Y(_1947_),
    .B1(net1100));
 sg13g2_a21oi_1 _4437_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1100),
    .A2(_1945_),
    .Y(_1948_),
    .B1(_1947_));
 sg13g2_nand2_1 _4438_ (.Y(_1949_),
    .A(net1094),
    .B(net404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4439_ (.A0(\s0.data_out[7][7] ),
    .A1(\s0.data_out[6][7] ),
    .S(net1095),
    .X(_1950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4440_ (.A(net1089),
    .B_N(net1144),
    .Y(_1951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4441_ (.A2(_1950_),
    .A1(net1089),
    .B1(_1951_),
    .X(_1952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4442_ (.Y(_1953_),
    .B(net404),
    .A_N(net1107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4443_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1840_),
    .A2(_1953_),
    .Y(_1954_),
    .B1(net1100));
 sg13g2_a21oi_1 _4444_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1100),
    .A2(_1952_),
    .Y(_1955_),
    .B1(_1954_));
 sg13g2_a22oi_1 _4445_ (.Y(_1956_),
    .B1(_1955_),
    .B2(net1402),
    .A2(_1948_),
    .A1(net1411),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4446_ (.A(net1411),
    .B(_1948_),
    .Y(_1957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4447_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1958_),
    .B(_1955_),
    .A(net1402));
 sg13g2_nand3b_1 _4448_ (.B(_1958_),
    .C(_1956_),
    .Y(_1959_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1957_));
 sg13g2_mux2_1 _4449_ (.A0(\s0.data_out[7][5] ),
    .A1(\s0.data_out[6][5] ),
    .S(net1095),
    .X(_1960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4450_ (.A(net1090),
    .B_N(net1153),
    .Y(_1961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4451_ (.A2(_1960_),
    .A1(net1090),
    .B1(_1961_),
    .X(_1962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4452_ (.Y(_1963_),
    .B(\s0.data_out[6][5] ),
    .A_N(net1107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4453_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1853_),
    .A2(_1963_),
    .Y(_1964_),
    .B1(net1101));
 sg13g2_a21oi_1 _4454_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1101),
    .A2(_1962_),
    .Y(_1965_),
    .B1(_1964_));
 sg13g2_nand2_1 _4455_ (.Y(_1966_),
    .A(net1421),
    .B(_1965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4456_ (.A(net1087),
    .B_N(net1158),
    .Y(_1967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4457_ (.A0(\s0.data_out[7][4] ),
    .A1(\s0.data_out[6][4] ),
    .S(net1092),
    .X(_1968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4458_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1087),
    .A2(_1968_),
    .Y(_1969_),
    .B1(_1967_));
 sg13g2_nand2b_1 _4459_ (.Y(_1970_),
    .B(net1097),
    .A_N(_1969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4460_ (.A0(\s0.data_out[6][4] ),
    .A1(\s0.data_out[7][4] ),
    .S(net1105),
    .X(_1971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4461_ (.Y(_1972_),
    .B(_1971_),
    .A_N(net1097),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4462_ (.B(_1970_),
    .C(_1972_),
    .A(net1431),
    .Y(_1973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4463_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1970_),
    .A2(_1972_),
    .Y(_1974_),
    .B1(net1431));
 sg13g2_nor2_1 _4464_ (.A(net1421),
    .B(_1965_),
    .Y(_1975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4465_ (.B1(_1966_),
    .VDD(VPWR),
    .Y(_1976_),
    .VSS(VGND),
    .A1(net1442),
    .A2(_1940_));
 sg13g2_nor2_1 _4466_ (.A(_1974_),
    .B(_1975_),
    .Y(_1977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4467_ (.Y(_1978_),
    .A(_1973_),
    .B(_1977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _4468_ (.A(_1941_),
    .B(_1959_),
    .C(_1976_),
    .D(_1978_),
    .X(_1979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4469_ (.B1(_1966_),
    .VDD(VPWR),
    .Y(_1980_),
    .VSS(VGND),
    .A1(_1973_),
    .A2(_1975_));
 sg13g2_nor2b_1 _4470_ (.A(_1959_),
    .B_N(_1980_),
    .Y(_1981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4471_ (.A(_1956_),
    .B_N(_1958_),
    .Y(_1982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4472_ (.A(_1904_),
    .B(_1981_),
    .C(_1982_),
    .Y(_1983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4473_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1984_),
    .B(net1331),
    .A(net344));
 sg13g2_a21oi_1 _4474_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1979_),
    .A2(_1983_),
    .Y(_0203_),
    .B1(_1984_));
 sg13g2_nor2_1 _4475_ (.A(net997),
    .B(_2864_),
    .Y(_1985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4476_ (.B1(net1096),
    .VDD(VPWR),
    .Y(_1986_),
    .VSS(VGND),
    .A1(_1926_),
    .A2(_1985_));
 sg13g2_nand3_1 _4477_ (.B(_1930_),
    .C(_1986_),
    .A(net1479),
    .Y(_1987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4478_ (.B1(_1987_),
    .VDD(VPWR),
    .Y(_1988_),
    .VSS(VGND),
    .A1(net1479),
    .A2(net521));
 sg13g2_inv_1 _4479_ (.VDD(VPWR),
    .Y(_0204_),
    .A(_1988_),
    .VSS(VGND));
 sg13g2_nor2_1 _4480_ (.A(net997),
    .B(_2863_),
    .Y(_1989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4481_ (.B1(net1096),
    .VDD(VPWR),
    .Y(_1990_),
    .VSS(VGND),
    .A1(_1920_),
    .A2(_1989_));
 sg13g2_nor2_1 _4482_ (.A(net1371),
    .B(_1923_),
    .Y(_1991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4483_ (.Y(_0205_),
    .B1(_1990_),
    .B2(_1991_),
    .A2(_2859_),
    .A1(net1371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4484_ (.A(net1086),
    .B(\s0.data_out[6][2] ),
    .X(_1992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4485_ (.B1(net1096),
    .VDD(VPWR),
    .Y(_1993_),
    .VSS(VGND),
    .A1(_1912_),
    .A2(_1992_));
 sg13g2_nor2_1 _4486_ (.A(net1371),
    .B(_1915_),
    .Y(_1994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4487_ (.Y(_0206_),
    .B1(_1993_),
    .B2(_1994_),
    .A2(_2858_),
    .A1(net1371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4488_ (.A(net998),
    .B(_2862_),
    .Y(_1995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4489_ (.B1(net1097),
    .VDD(VPWR),
    .Y(_1996_),
    .VSS(VGND),
    .A1(_1936_),
    .A2(_1995_));
 sg13g2_nor2_1 _4490_ (.A(net1371),
    .B(net390),
    .Y(_1997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4491_ (.Y(_0207_),
    .B1(_1996_),
    .B2(_1997_),
    .A2(_2857_),
    .A1(net1371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4492_ (.A(net1087),
    .B(\s0.data_out[6][4] ),
    .X(_1998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4493_ (.B1(net1097),
    .VDD(VPWR),
    .Y(_1999_),
    .VSS(VGND),
    .A1(_1967_),
    .A2(_1998_));
 sg13g2_nand3_1 _4494_ (.B(_1972_),
    .C(_1999_),
    .A(net1479),
    .Y(_2000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4495_ (.B1(_2000_),
    .VDD(VPWR),
    .Y(_2001_),
    .VSS(VGND),
    .A1(net1479),
    .A2(net639));
 sg13g2_inv_1 _4496_ (.VDD(VPWR),
    .Y(_0208_),
    .A(_2001_),
    .VSS(VGND));
 sg13g2_and2_1 _4497_ (.A(net1090),
    .B(\s0.data_out[6][5] ),
    .X(_2002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4498_ (.B1(net1101),
    .VDD(VPWR),
    .Y(_2003_),
    .VSS(VGND),
    .A1(_1961_),
    .A2(_2002_));
 sg13g2_nor2_1 _4499_ (.A(net1372),
    .B(_1964_),
    .Y(_2004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4500_ (.Y(_0209_),
    .B1(_2003_),
    .B2(_2004_),
    .A2(_2856_),
    .A1(net1372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4501_ (.A(net998),
    .B(_2861_),
    .Y(_2005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4502_ (.B1(net1100),
    .VDD(VPWR),
    .Y(_2006_),
    .VSS(VGND),
    .A1(_1944_),
    .A2(_2005_));
 sg13g2_nand3b_1 _4503_ (.B(_2006_),
    .C(net1480),
    .Y(_2007_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1947_));
 sg13g2_o21ai_1 _4504_ (.B1(_2007_),
    .VDD(VPWR),
    .Y(_2008_),
    .VSS(VGND),
    .A1(net1480),
    .A2(net627));
 sg13g2_inv_1 _4505_ (.VDD(VPWR),
    .Y(_0210_),
    .A(_2008_),
    .VSS(VGND));
 sg13g2_nor2_1 _4506_ (.A(net998),
    .B(_2860_),
    .Y(_2009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4507_ (.B1(net1100),
    .VDD(VPWR),
    .Y(_2010_),
    .VSS(VGND),
    .A1(_1951_),
    .A2(_2009_));
 sg13g2_nor2_1 _4508_ (.A(net1372),
    .B(_1954_),
    .Y(_2011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4509_ (.Y(_0211_),
    .B1(_2010_),
    .B2(_2011_),
    .A2(_2855_),
    .A1(net1373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4510_ (.B1(net1088),
    .VDD(VPWR),
    .Y(_2012_),
    .VSS(VGND),
    .A1(net1396),
    .A2(net1078));
 sg13g2_a21oi_1 _4511_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1337),
    .A2(net1082),
    .Y(_2013_),
    .B1(_2012_));
 sg13g2_a21oi_1 _4512_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net998),
    .A2(_1902_),
    .Y(_2014_),
    .B1(_2013_));
 sg13g2_o21ai_1 _4513_ (.B1(_2013_),
    .VDD(VPWR),
    .Y(_2015_),
    .VSS(VGND),
    .A1(net345),
    .A2(net1083));
 sg13g2_nor2_1 _4514_ (.A(net1078),
    .B(_2012_),
    .Y(_2016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4515_ (.B1(net998),
    .VDD(VPWR),
    .Y(_2017_),
    .VSS(VGND),
    .A1(net345),
    .A2(net1094));
 sg13g2_nand2_1 _4516_ (.Y(_2018_),
    .A(_2015_),
    .B(_2017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4517_ (.B1(net1479),
    .VDD(VPWR),
    .Y(_2019_),
    .VSS(VGND),
    .A1(_2016_),
    .A2(_2018_));
 sg13g2_a21oi_1 _4518_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2731_),
    .A2(_2014_),
    .Y(_0212_),
    .B1(_2019_));
 sg13g2_and2_1 _4519_ (.A(net1479),
    .B(_2014_),
    .X(_0213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4520_ (.A(net1474),
    .B(net331),
    .X(_0214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4521_ (.Y(_2020_),
    .A(net1080),
    .B(net656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4522_ (.A0(\s0.data_out[6][1] ),
    .A1(\s0.data_out[5][1] ),
    .S(net1081),
    .X(_2021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4523_ (.A(net1074),
    .B_N(net1169),
    .Y(_2022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4524_ (.A2(_2021_),
    .A1(net1074),
    .B1(_2022_),
    .X(_2023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4525_ (.Y(_2024_),
    .B(\s0.data_out[5][1] ),
    .A_N(net1092),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4526_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1918_),
    .A2(_2024_),
    .Y(_2025_),
    .B1(net1085));
 sg13g2_a21oi_1 _4527_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1085),
    .A2(_2023_),
    .Y(_2026_),
    .B1(_2025_));
 sg13g2_mux2_1 _4528_ (.A0(net571),
    .A1(net692),
    .S(net1092),
    .X(_2027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4529_ (.Y(_2028_),
    .A(net997),
    .B(_2027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4530_ (.A(net1074),
    .B_N(net1172),
    .Y(_2029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4531_ (.A0(\s0.data_out[6][0] ),
    .A1(\s0.data_out[5][0] ),
    .S(net1081),
    .X(_2030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4532_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1075),
    .A2(_2030_),
    .Y(_2031_),
    .B1(_2029_));
 sg13g2_nand2b_1 _4533_ (.Y(_2032_),
    .B(net1085),
    .A_N(_2031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4534_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2032_),
    .C1(net1460),
    .B1(_2028_),
    .A1(net1452),
    .Y(_2033_),
    .A2(_2026_));
 sg13g2_nor2_1 _4535_ (.A(net1452),
    .B(_2026_),
    .Y(_2034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4536_ (.Y(_2035_),
    .A(net1080),
    .B(net549),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4537_ (.A0(\s0.data_out[6][3] ),
    .A1(\s0.data_out[5][3] ),
    .S(net1081),
    .X(_2036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4538_ (.A(net1075),
    .B_N(net1161),
    .Y(_2037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4539_ (.A2(_2036_),
    .A1(net1075),
    .B1(_2037_),
    .X(_2038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4540_ (.Y(_2039_),
    .B(\s0.data_out[5][3] ),
    .A_N(net1093),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4541_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1934_),
    .A2(_2039_),
    .Y(_2040_),
    .B1(net1091));
 sg13g2_a21oi_1 _4542_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1087),
    .A2(_2038_),
    .Y(_2041_),
    .B1(_2040_));
 sg13g2_nor2_1 _4543_ (.A(net1439),
    .B(_2041_),
    .Y(_2042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4544_ (.Y(_2043_),
    .A(net1080),
    .B(\s0.data_out[5][2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4545_ (.A0(\s0.data_out[6][2] ),
    .A1(\s0.data_out[5][2] ),
    .S(net1081),
    .X(_2044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4546_ (.A(net1074),
    .B_N(net1165),
    .Y(_2045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4547_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1074),
    .A2(_2044_),
    .Y(_2046_),
    .B1(_2045_));
 sg13g2_mux2_1 _4548_ (.A0(\s0.data_out[5][2] ),
    .A1(\s0.data_out[6][2] ),
    .S(net1092),
    .X(_2047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4549_ (.Y(_2048_),
    .A(net997),
    .B(_2047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4550_ (.B1(_2048_),
    .VDD(VPWR),
    .Y(_2049_),
    .VSS(VGND),
    .A1(net997),
    .A2(_2046_));
 sg13g2_or2_1 _4551_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2050_),
    .B(_2049_),
    .A(net1335));
 sg13g2_xnor2_1 _4552_ (.Y(_2051_),
    .A(net1335),
    .B(_2049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _4553_ (.A(_2033_),
    .B(_2034_),
    .C(_2042_),
    .D(_2051_),
    .Y(_2052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4554_ (.Y(_2053_),
    .A(net1439),
    .B(_2041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4555_ (.B1(_2053_),
    .VDD(VPWR),
    .Y(_2054_),
    .VSS(VGND),
    .A1(_2042_),
    .A2(_2050_));
 sg13g2_nor2_1 _4556_ (.A(_2052_),
    .B(_2054_),
    .Y(_2055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4557_ (.Y(_2056_),
    .A(net1082),
    .B(net488),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4558_ (.A0(\s0.data_out[6][7] ),
    .A1(\s0.data_out[5][7] ),
    .S(net1083),
    .X(_2057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4559_ (.A(net1078),
    .B_N(net1144),
    .Y(_2058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4560_ (.A2(_2057_),
    .A1(net1078),
    .B1(_2058_),
    .X(_2059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4561_ (.Y(_2060_),
    .B(\s0.data_out[5][7] ),
    .A_N(net1094),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4562_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1949_),
    .A2(_2060_),
    .Y(_2061_),
    .B1(net1088));
 sg13g2_a21oi_1 _4563_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1088),
    .A2(_2059_),
    .Y(_2062_),
    .B1(_2061_));
 sg13g2_nand2_1 _4564_ (.Y(_2063_),
    .A(net1082),
    .B(net449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4565_ (.A0(\s0.data_out[6][6] ),
    .A1(\s0.data_out[5][6] ),
    .S(net1083),
    .X(_2064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4566_ (.A(net1078),
    .B_N(net1148),
    .Y(_2065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4567_ (.A2(_2064_),
    .A1(net1079),
    .B1(_2065_),
    .X(_2066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4568_ (.Y(_2067_),
    .B(net449),
    .A_N(net1094),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4569_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1942_),
    .A2(_2067_),
    .Y(_2068_),
    .B1(net1088));
 sg13g2_a21oi_1 _4570_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1088),
    .A2(_2066_),
    .Y(_2069_),
    .B1(_2068_));
 sg13g2_a22oi_1 _4571_ (.Y(_2070_),
    .B1(_2069_),
    .B2(net1412),
    .A2(_2062_),
    .A1(net1403),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4572_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2071_),
    .B(_2069_),
    .A(net1412));
 sg13g2_nor2_1 _4573_ (.A(net1403),
    .B(_2062_),
    .Y(_2072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _4574_ (.B(_2070_),
    .C(_2071_),
    .Y(_2073_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2072_));
 sg13g2_nor2b_1 _4575_ (.A(net1075),
    .B_N(net1158),
    .Y(_2074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4576_ (.A0(\s0.data_out[6][4] ),
    .A1(\s0.data_out[5][4] ),
    .S(net1081),
    .X(_2075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4577_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1075),
    .A2(_2075_),
    .Y(_2076_),
    .B1(_2074_));
 sg13g2_nand2b_1 _4578_ (.Y(_2077_),
    .B(net1090),
    .A_N(_2076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4579_ (.A0(\s0.data_out[5][4] ),
    .A1(\s0.data_out[6][4] ),
    .S(net1093),
    .X(_2078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4580_ (.Y(_2079_),
    .A(net999),
    .B(_2078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4581_ (.B(_2077_),
    .C(_2079_),
    .A(net1430),
    .Y(_2080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4582_ (.A0(\s0.data_out[6][5] ),
    .A1(\s0.data_out[5][5] ),
    .S(net1083),
    .X(_2081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4583_ (.A(net1078),
    .B_N(net1153),
    .Y(_2082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4584_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1078),
    .A2(_2081_),
    .Y(_2083_),
    .B1(_2082_));
 sg13g2_nand2b_1 _4585_ (.Y(_2084_),
    .B(net1090),
    .A_N(_2083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4586_ (.A0(\s0.data_out[5][5] ),
    .A1(\s0.data_out[6][5] ),
    .S(net1095),
    .X(_2085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4587_ (.Y(_2086_),
    .A(net999),
    .B(_2085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4588_ (.B(_2084_),
    .C(_2086_),
    .A(net1422),
    .Y(_2087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4589_ (.Y(_2088_),
    .A(_2080_),
    .B(_2087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4590_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2077_),
    .A2(_2079_),
    .Y(_2089_),
    .B1(net1430));
 sg13g2_a21oi_1 _4591_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2084_),
    .A2(_2086_),
    .Y(_2090_),
    .B1(net1422));
 sg13g2_or2_1 _4592_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2091_),
    .B(_2090_),
    .A(_2089_));
 sg13g2_or4_1 _4593_ (.A(_2055_),
    .B(_2073_),
    .C(_2088_),
    .D(_2091_),
    .X(_2092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4594_ (.B1(_2087_),
    .VDD(VPWR),
    .Y(_2093_),
    .VSS(VGND),
    .A1(_2080_),
    .A2(_2090_));
 sg13g2_nand2b_1 _4595_ (.Y(_2094_),
    .B(_2093_),
    .A_N(_2073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4596_ (.B1(_2014_),
    .VDD(VPWR),
    .Y(_2095_),
    .VSS(VGND),
    .A1(_2070_),
    .A2(_2072_));
 sg13g2_nor2b_1 _4597_ (.A(_2095_),
    .B_N(_2094_),
    .Y(_2096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4598_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2097_),
    .B(net1331),
    .A(net339));
 sg13g2_a21oi_1 _4599_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2092_),
    .A2(_2096_),
    .Y(_0215_),
    .B1(_2097_));
 sg13g2_and2_1 _4600_ (.A(net1074),
    .B(net571),
    .X(_2098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4601_ (.B1(net1085),
    .VDD(VPWR),
    .Y(_2099_),
    .VSS(VGND),
    .A1(_2029_),
    .A2(_2098_));
 sg13g2_a21oi_1 _4602_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net997),
    .A2(_2027_),
    .Y(_2100_),
    .B1(net1370));
 sg13g2_a22oi_1 _4603_ (.Y(_0216_),
    .B1(_2099_),
    .B2(_2100_),
    .A2(_2864_),
    .A1(net1370),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4604_ (.A(net1074),
    .B(\s0.data_out[5][1] ),
    .X(_2101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4605_ (.B1(net1085),
    .VDD(VPWR),
    .Y(_2102_),
    .VSS(VGND),
    .A1(_2022_),
    .A2(_2101_));
 sg13g2_nor2_1 _4606_ (.A(net1370),
    .B(_2025_),
    .Y(_2103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4607_ (.Y(_0217_),
    .B1(_2102_),
    .B2(_2103_),
    .A2(_2863_),
    .A1(net1370),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4608_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1074),
    .A2(net606),
    .Y(_2104_),
    .B1(_2045_));
 sg13g2_a21oi_1 _4609_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net997),
    .A2(_2047_),
    .Y(_2105_),
    .B1(net1370));
 sg13g2_o21ai_1 _4610_ (.B1(_2105_),
    .VDD(VPWR),
    .Y(_2106_),
    .VSS(VGND),
    .A1(net997),
    .A2(_2104_));
 sg13g2_o21ai_1 _4611_ (.B1(_2106_),
    .VDD(VPWR),
    .Y(_2107_),
    .VSS(VGND),
    .A1(net1479),
    .A2(net682));
 sg13g2_inv_1 _4612_ (.VDD(VPWR),
    .Y(_0218_),
    .A(_2107_),
    .VSS(VGND));
 sg13g2_and2_1 _4613_ (.A(net1075),
    .B(\s0.data_out[5][3] ),
    .X(_2108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4614_ (.B1(net1091),
    .VDD(VPWR),
    .Y(_2109_),
    .VSS(VGND),
    .A1(_2037_),
    .A2(_2108_));
 sg13g2_nor2_1 _4615_ (.A(net1370),
    .B(_2040_),
    .Y(_2110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4616_ (.Y(_0219_),
    .B1(net447),
    .B2(_2110_),
    .A2(_2862_),
    .A1(net1370),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4617_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1075),
    .A2(net570),
    .Y(_2111_),
    .B1(_2074_));
 sg13g2_a21oi_1 _4618_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net998),
    .A2(_2078_),
    .Y(_2112_),
    .B1(net1370));
 sg13g2_o21ai_1 _4619_ (.B1(_2112_),
    .VDD(VPWR),
    .Y(_2113_),
    .VSS(VGND),
    .A1(net998),
    .A2(_2111_));
 sg13g2_o21ai_1 _4620_ (.B1(_2113_),
    .VDD(VPWR),
    .Y(_2114_),
    .VSS(VGND),
    .A1(net1479),
    .A2(net669));
 sg13g2_inv_1 _4621_ (.VDD(VPWR),
    .Y(_0220_),
    .A(_2114_),
    .VSS(VGND));
 sg13g2_a21oi_1 _4622_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1078),
    .A2(net568),
    .Y(_2115_),
    .B1(_2082_));
 sg13g2_a21oi_1 _4623_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net999),
    .A2(_2085_),
    .Y(_2116_),
    .B1(net1372));
 sg13g2_o21ai_1 _4624_ (.B1(_2116_),
    .VDD(VPWR),
    .Y(_2117_),
    .VSS(VGND),
    .A1(net999),
    .A2(_2115_));
 sg13g2_o21ai_1 _4625_ (.B1(_2117_),
    .VDD(VPWR),
    .Y(_2118_),
    .VSS(VGND),
    .A1(net1480),
    .A2(net630));
 sg13g2_inv_1 _4626_ (.VDD(VPWR),
    .Y(_0221_),
    .A(_2118_),
    .VSS(VGND));
 sg13g2_and2_1 _4627_ (.A(net1079),
    .B(net449),
    .X(_2119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4628_ (.B1(net1088),
    .VDD(VPWR),
    .Y(_2120_),
    .VSS(VGND),
    .A1(_2065_),
    .A2(_2119_));
 sg13g2_nor2_1 _4629_ (.A(net1372),
    .B(_2068_),
    .Y(_2121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4630_ (.Y(_0222_),
    .B1(_2120_),
    .B2(_2121_),
    .A2(_2861_),
    .A1(net1372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4631_ (.A(net1079),
    .B(net488),
    .X(_2122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4632_ (.B1(net1088),
    .VDD(VPWR),
    .Y(_2123_),
    .VSS(VGND),
    .A1(_2058_),
    .A2(_2122_));
 sg13g2_nor2_1 _4633_ (.A(net1372),
    .B(net405),
    .Y(_2124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4634_ (.Y(_0223_),
    .B1(_2123_),
    .B2(_2124_),
    .A2(_2860_),
    .A1(net1372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4635_ (.B1(net1076),
    .VDD(VPWR),
    .Y(_2125_),
    .VSS(VGND),
    .A1(net1393),
    .A2(net1065));
 sg13g2_a21oi_1 _4636_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1336),
    .A2(net1070),
    .Y(_2126_),
    .B1(_2125_));
 sg13g2_a21oi_1 _4637_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1336),
    .A2(net1082),
    .Y(_2127_),
    .B1(net1076));
 sg13g2_nor2_1 _4638_ (.A(_2126_),
    .B(_2127_),
    .Y(_2128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4639_ (.B1(_2126_),
    .VDD(VPWR),
    .Y(_2129_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[4] [0]),
    .A2(net1070));
 sg13g2_nor2_1 _4640_ (.A(net1065),
    .B(_2125_),
    .Y(_2130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4641_ (.A(\s0.was_valid_out[4] [0]),
    .B(net1082),
    .Y(_2131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4642_ (.B1(_2129_),
    .VDD(VPWR),
    .Y(_2132_),
    .VSS(VGND),
    .A1(net1077),
    .A2(_2131_));
 sg13g2_o21ai_1 _4643_ (.B1(net1474),
    .VDD(VPWR),
    .Y(_2133_),
    .VSS(VGND),
    .A1(_2130_),
    .A2(_2132_));
 sg13g2_a21oi_1 _4644_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2730_),
    .A2(_2128_),
    .Y(_0224_),
    .B1(_2133_));
 sg13g2_nor3_1 _4645_ (.A(net1363),
    .B(_2126_),
    .C(_2127_),
    .Y(_0225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4646_ (.A(net1475),
    .B(net321),
    .X(_0226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4647_ (.Y(_2134_),
    .A(net1067),
    .B(net642),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4648_ (.B1(_2134_),
    .VDD(VPWR),
    .Y(_2135_),
    .VSS(VGND),
    .A1(net1068),
    .A2(_2865_));
 sg13g2_nor2b_1 _4649_ (.A(net1061),
    .B_N(net1167),
    .Y(_2136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4650_ (.A2(_2135_),
    .A1(net1061),
    .B1(_2136_),
    .X(_2137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4651_ (.Y(_2138_),
    .B(net642),
    .A_N(net1080),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4652_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2020_),
    .A2(_2138_),
    .Y(_2139_),
    .B1(net1072));
 sg13g2_a21oi_1 _4653_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1072),
    .A2(_2137_),
    .Y(_2140_),
    .B1(_2139_));
 sg13g2_mux2_1 _4654_ (.A0(\s0.data_out[4][0] ),
    .A1(\s0.data_out[5][0] ),
    .S(net1080),
    .X(_2141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4655_ (.Y(_2142_),
    .B(_2141_),
    .A_N(net1072),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4656_ (.A(net1061),
    .B_N(net1172),
    .Y(_2143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4657_ (.A0(\s0.data_out[5][0] ),
    .A1(\s0.data_out[4][0] ),
    .S(net1068),
    .X(_2144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4658_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1061),
    .A2(_2144_),
    .Y(_2145_),
    .B1(_2143_));
 sg13g2_nand2b_1 _4659_ (.Y(_2146_),
    .B(net1072),
    .A_N(_2145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4660_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2146_),
    .C1(net1460),
    .B1(_2142_),
    .A1(net1452),
    .Y(_2147_),
    .A2(_2140_));
 sg13g2_nand2_1 _4661_ (.Y(_2148_),
    .A(net1067),
    .B(net676),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4662_ (.A0(\s0.data_out[5][2] ),
    .A1(\s0.data_out[4][2] ),
    .S(net1068),
    .X(_2149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4663_ (.A(net1061),
    .B_N(net1163),
    .Y(_2150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4664_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1061),
    .A2(_2149_),
    .Y(_2151_),
    .B1(_2150_));
 sg13g2_nand2b_1 _4665_ (.Y(_2152_),
    .B(net1072),
    .A_N(_2151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4666_ (.B1(_2043_),
    .VDD(VPWR),
    .Y(_2153_),
    .VSS(VGND),
    .A1(net1080),
    .A2(_2872_));
 sg13g2_nand2b_1 _4667_ (.Y(_2154_),
    .B(_2153_),
    .A_N(net1072),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4668_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2152_),
    .A2(_2154_),
    .Y(_2155_),
    .B1(net1447));
 sg13g2_nand2_1 _4669_ (.Y(_2156_),
    .A(net1068),
    .B(net444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4670_ (.B1(_2156_),
    .VDD(VPWR),
    .Y(_2157_),
    .VSS(VGND),
    .A1(net1068),
    .A2(_2866_));
 sg13g2_nor2_1 _4671_ (.A(net1062),
    .B(net993),
    .Y(_2158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4672_ (.A2(_2157_),
    .A1(net1062),
    .B1(_2158_),
    .X(_2159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4673_ (.Y(_2160_),
    .B(net444),
    .A_N(net1080),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4674_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2035_),
    .A2(_2160_),
    .Y(_2161_),
    .B1(net1073));
 sg13g2_a21oi_1 _4675_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1073),
    .A2(_2159_),
    .Y(_2162_),
    .B1(_2161_));
 sg13g2_nor2_1 _4676_ (.A(net1439),
    .B(_2162_),
    .Y(_2163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4677_ (.B(_2152_),
    .C(_2154_),
    .A(net1447),
    .Y(_2164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4678_ (.B1(_2164_),
    .VDD(VPWR),
    .Y(_2165_),
    .VSS(VGND),
    .A1(net1452),
    .A2(_2140_));
 sg13g2_nor4_1 _4679_ (.A(_2147_),
    .B(_2155_),
    .C(_2163_),
    .D(_2165_),
    .Y(_2166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4680_ (.Y(_2167_),
    .A(net1439),
    .B(_2162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4681_ (.B1(_2167_),
    .VDD(VPWR),
    .Y(_2168_),
    .VSS(VGND),
    .A1(_2163_),
    .A2(_2164_));
 sg13g2_nand2_1 _4682_ (.Y(_2169_),
    .A(net1069),
    .B(net507),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4683_ (.A0(\s0.data_out[5][6] ),
    .A1(\s0.data_out[4][6] ),
    .S(net1070),
    .X(_2170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4684_ (.A(net1065),
    .B_N(net1148),
    .Y(_2171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4685_ (.A2(_2170_),
    .A1(net1065),
    .B1(_2171_),
    .X(_2172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4686_ (.Y(_2173_),
    .B(\s0.data_out[4][6] ),
    .A_N(net1082),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4687_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2063_),
    .A2(_2173_),
    .Y(_2174_),
    .B1(net1076));
 sg13g2_a21oi_1 _4688_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1076),
    .A2(_2172_),
    .Y(_2175_),
    .B1(_2174_));
 sg13g2_nand2_1 _4689_ (.Y(_2176_),
    .A(net1069),
    .B(net492),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4690_ (.A0(\s0.data_out[5][7] ),
    .A1(\s0.data_out[4][7] ),
    .S(net1070),
    .X(_2177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4691_ (.A(net1065),
    .B_N(net1143),
    .Y(_2178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4692_ (.A2(_2177_),
    .A1(net1066),
    .B1(_2178_),
    .X(_2179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4693_ (.Y(_2180_),
    .B(net492),
    .A_N(net1082),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4694_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2056_),
    .A2(_2180_),
    .Y(_2181_),
    .B1(net1076));
 sg13g2_a21oi_1 _4695_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1076),
    .A2(_2179_),
    .Y(_2182_),
    .B1(_2181_));
 sg13g2_a22oi_1 _4696_ (.Y(_2183_),
    .B1(_2182_),
    .B2(net1400),
    .A2(_2175_),
    .A1(net1409),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4697_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2184_),
    .B(_2175_),
    .A(net1410));
 sg13g2_nor2_1 _4698_ (.A(net1400),
    .B(_2182_),
    .Y(_2185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _4699_ (.B(_2183_),
    .C(_2184_),
    .Y(_2186_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2185_));
 sg13g2_nor2b_1 _4700_ (.A(net1062),
    .B_N(net1157),
    .Y(_2187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4701_ (.Y(_2188_),
    .A(net1067),
    .B(\s0.data_out[4][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4702_ (.A0(\s0.data_out[5][4] ),
    .A1(\s0.data_out[4][4] ),
    .S(net1068),
    .X(_2189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4703_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1062),
    .A2(_2189_),
    .Y(_2190_),
    .B1(_2187_));
 sg13g2_nand2b_1 _4704_ (.Y(_2191_),
    .B(net1073),
    .A_N(_2190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4705_ (.A0(\s0.data_out[4][4] ),
    .A1(\s0.data_out[5][4] ),
    .S(net1080),
    .X(_2192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4706_ (.Y(_2193_),
    .B(_2192_),
    .A_N(net1073),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4707_ (.B(_2191_),
    .C(_2193_),
    .A(net1427),
    .Y(_2194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4708_ (.Y(_2195_),
    .A(net1069),
    .B(\s0.data_out[4][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4709_ (.A0(\s0.data_out[5][5] ),
    .A1(\s0.data_out[4][5] ),
    .S(net1070),
    .X(_2196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4710_ (.A(net1065),
    .B_N(net1151),
    .Y(_2197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4711_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1065),
    .A2(_2196_),
    .Y(_2198_),
    .B1(_2197_));
 sg13g2_nand2b_1 _4712_ (.Y(_2199_),
    .B(net1077),
    .A_N(_2198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4713_ (.A0(\s0.data_out[4][5] ),
    .A1(\s0.data_out[5][5] ),
    .S(net1082),
    .X(_2200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4714_ (.Y(_2201_),
    .B(_2200_),
    .A_N(net1077),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4715_ (.B(_2199_),
    .C(_2201_),
    .A(net1418),
    .Y(_2202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4716_ (.Y(_2203_),
    .A(_2194_),
    .B(_2202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4717_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2191_),
    .A2(_2193_),
    .Y(_2204_),
    .B1(net1427));
 sg13g2_a21oi_1 _4718_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2199_),
    .A2(_2201_),
    .Y(_2205_),
    .B1(net1418));
 sg13g2_nor4_1 _4719_ (.A(_2186_),
    .B(_2203_),
    .C(_2204_),
    .D(_2205_),
    .Y(_2206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4720_ (.B1(_2206_),
    .VDD(VPWR),
    .Y(_2207_),
    .VSS(VGND),
    .A1(_2166_),
    .A2(_2168_));
 sg13g2_o21ai_1 _4721_ (.B1(_2202_),
    .VDD(VPWR),
    .Y(_2208_),
    .VSS(VGND),
    .A1(_2194_),
    .A2(_2205_));
 sg13g2_nor2b_1 _4722_ (.A(_2186_),
    .B_N(_2208_),
    .Y(_2209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4723_ (.B1(_2128_),
    .VDD(VPWR),
    .Y(_2210_),
    .VSS(VGND),
    .A1(_2183_),
    .A2(_2185_));
 sg13g2_nor2_1 _4724_ (.A(_2209_),
    .B(_2210_),
    .Y(_2211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4725_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2212_),
    .B(net1329),
    .A(net331));
 sg13g2_a21oi_1 _4726_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2207_),
    .A2(_2211_),
    .Y(_0227_),
    .B1(_2212_));
 sg13g2_and2_1 _4727_ (.A(net1061),
    .B(\s0.data_out[4][0] ),
    .X(_2213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4728_ (.B1(net1073),
    .VDD(VPWR),
    .Y(_2214_),
    .VSS(VGND),
    .A1(_2143_),
    .A2(_2213_));
 sg13g2_nand3_1 _4729_ (.B(_2142_),
    .C(_2214_),
    .A(net1474),
    .Y(_2215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4730_ (.B1(_2215_),
    .VDD(VPWR),
    .Y(_2216_),
    .VSS(VGND),
    .A1(net1474),
    .A2(net571));
 sg13g2_inv_1 _4731_ (.VDD(VPWR),
    .Y(_0228_),
    .A(_2216_),
    .VSS(VGND));
 sg13g2_nor2_1 _4732_ (.A(net995),
    .B(_2873_),
    .Y(_2217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4733_ (.B1(net1072),
    .VDD(VPWR),
    .Y(_2218_),
    .VSS(VGND),
    .A1(_2136_),
    .A2(_2217_));
 sg13g2_nor2_1 _4734_ (.A(net1363),
    .B(_2139_),
    .Y(_2219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4735_ (.Y(_0229_),
    .B1(_2218_),
    .B2(_2219_),
    .A2(_2865_),
    .A1(net1363),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4736_ (.A(net995),
    .B(_2872_),
    .Y(_2220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4737_ (.B1(net1072),
    .VDD(VPWR),
    .Y(_2221_),
    .VSS(VGND),
    .A1(_2150_),
    .A2(_2220_));
 sg13g2_nand3_1 _4738_ (.B(_2154_),
    .C(_2221_),
    .A(net1474),
    .Y(_2222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4739_ (.B1(_2222_),
    .VDD(VPWR),
    .Y(_2223_),
    .VSS(VGND),
    .A1(net1474),
    .A2(net606));
 sg13g2_inv_1 _4740_ (.VDD(VPWR),
    .Y(_0230_),
    .A(_2223_),
    .VSS(VGND));
 sg13g2_nor2_1 _4741_ (.A(net995),
    .B(_2871_),
    .Y(_2224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4742_ (.B1(net1073),
    .VDD(VPWR),
    .Y(_2225_),
    .VSS(VGND),
    .A1(_2158_),
    .A2(_2224_));
 sg13g2_nor2_1 _4743_ (.A(net1363),
    .B(_2161_),
    .Y(_2226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4744_ (.Y(_0231_),
    .B1(_2225_),
    .B2(_2226_),
    .A2(_2866_),
    .A1(net1363),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4745_ (.A(net1061),
    .B(\s0.data_out[4][4] ),
    .X(_2227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4746_ (.B1(net1073),
    .VDD(VPWR),
    .Y(_2228_),
    .VSS(VGND),
    .A1(_2187_),
    .A2(_2227_));
 sg13g2_nand3_1 _4747_ (.B(_2193_),
    .C(_2228_),
    .A(net1474),
    .Y(_2229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4748_ (.B1(_2229_),
    .VDD(VPWR),
    .Y(_2230_),
    .VSS(VGND),
    .A1(net1474),
    .A2(net570));
 sg13g2_inv_1 _4749_ (.VDD(VPWR),
    .Y(_0232_),
    .A(_2230_),
    .VSS(VGND));
 sg13g2_and2_1 _4750_ (.A(net1065),
    .B(\s0.data_out[4][5] ),
    .X(_2231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4751_ (.B1(net1077),
    .VDD(VPWR),
    .Y(_2232_),
    .VSS(VGND),
    .A1(_2197_),
    .A2(_2231_));
 sg13g2_nand3_1 _4752_ (.B(_2201_),
    .C(_2232_),
    .A(net1475),
    .Y(_2233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4753_ (.B1(_2233_),
    .VDD(VPWR),
    .Y(_2234_),
    .VSS(VGND),
    .A1(net1475),
    .A2(net568));
 sg13g2_inv_1 _4754_ (.VDD(VPWR),
    .Y(_0233_),
    .A(_2234_),
    .VSS(VGND));
 sg13g2_nor2_1 _4755_ (.A(net996),
    .B(_2870_),
    .Y(_2235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4756_ (.B1(net1076),
    .VDD(VPWR),
    .Y(_2236_),
    .VSS(VGND),
    .A1(_2171_),
    .A2(_2235_));
 sg13g2_nor2_1 _4757_ (.A(net1363),
    .B(_2174_),
    .Y(_2237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4758_ (.Y(_0234_),
    .B1(_2236_),
    .B2(_2237_),
    .A2(_2868_),
    .A1(net1363),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4759_ (.A(net996),
    .B(_2869_),
    .Y(_2238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4760_ (.B1(net1076),
    .VDD(VPWR),
    .Y(_2239_),
    .VSS(VGND),
    .A1(_2178_),
    .A2(_2238_));
 sg13g2_nor2_1 _4761_ (.A(net1363),
    .B(_2181_),
    .Y(_2240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4762_ (.Y(_0235_),
    .B1(_2239_),
    .B2(_2240_),
    .A2(_2867_),
    .A1(net1364),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4763_ (.B1(net1064),
    .VDD(VPWR),
    .Y(_2241_),
    .VSS(VGND),
    .A1(net1393),
    .A2(net1054));
 sg13g2_nor2_1 _4764_ (.A(net1397),
    .B(_2748_),
    .Y(_2242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4765_ (.A(_2241_),
    .B(_2242_),
    .Y(_2243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4766_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1338),
    .A2(net1069),
    .Y(_2244_),
    .B1(net1064));
 sg13g2_nor2_1 _4767_ (.A(_2243_),
    .B(_2244_),
    .Y(_2245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4768_ (.Y(_2246_),
    .B(_2245_),
    .A_N(net699),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4769_ (.B1(_2243_),
    .VDD(VPWR),
    .Y(_2247_),
    .VSS(VGND),
    .A1(net524),
    .A2(net1059));
 sg13g2_or2_1 _4770_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2248_),
    .B(_2241_),
    .A(net1054));
 sg13g2_o21ai_1 _4771_ (.B1(net996),
    .VDD(VPWR),
    .Y(_2249_),
    .VSS(VGND),
    .A1(net524),
    .A2(net1069));
 sg13g2_nand3_1 _4772_ (.B(_2248_),
    .C(_2249_),
    .A(_2247_),
    .Y(_2250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4773_ (.X(_0236_),
    .A(net1473),
    .B(_2246_),
    .C(_2250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4774_ (.A(net1361),
    .B(_2243_),
    .C(_2244_),
    .Y(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4775_ (.A(net1473),
    .B(net340),
    .X(_0238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4776_ (.Y(_2251_),
    .A(net1056),
    .B(net434),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4777_ (.A0(\s0.data_out[4][2] ),
    .A1(\s0.data_out[3][2] ),
    .S(net1057),
    .X(_2252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4778_ (.A(net1049),
    .B_N(net1163),
    .Y(_2253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4779_ (.A2(_2252_),
    .A1(net1049),
    .B1(_2253_),
    .X(_2254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4780_ (.Y(_2255_),
    .B(net434),
    .A_N(net1067),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4781_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2148_),
    .A2(_2255_),
    .Y(_2256_),
    .B1(net1060));
 sg13g2_a21oi_1 _4782_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1060),
    .A2(_2254_),
    .Y(_2257_),
    .B1(_2256_));
 sg13g2_or2_1 _4783_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2258_),
    .B(_2257_),
    .A(net1444));
 sg13g2_nand2_1 _4784_ (.Y(_2259_),
    .A(net1056),
    .B(net400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4785_ (.B1(_2259_),
    .VDD(VPWR),
    .Y(_2260_),
    .VSS(VGND),
    .A1(net1057),
    .A2(_2873_));
 sg13g2_nor2b_1 _4786_ (.A(net1049),
    .B_N(net1167),
    .Y(_2261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4787_ (.A2(_2260_),
    .A1(net1049),
    .B1(_2261_),
    .X(_2262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4788_ (.Y(_2263_),
    .B(net400),
    .A_N(net1067),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4789_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2134_),
    .A2(_2263_),
    .Y(_2264_),
    .B1(net1060));
 sg13g2_a21oi_1 _4790_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1060),
    .A2(_2262_),
    .Y(_2265_),
    .B1(_2264_));
 sg13g2_mux2_1 _4791_ (.A0(\s0.data_out[4][0] ),
    .A1(\s0.data_out[3][0] ),
    .S(net1057),
    .X(_2266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4792_ (.A(net1050),
    .B_N(net1170),
    .Y(_2267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4793_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1049),
    .A2(_2266_),
    .Y(_2268_),
    .B1(_2267_));
 sg13g2_nand2b_1 _4794_ (.Y(_2269_),
    .B(net1060),
    .A_N(_2268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4795_ (.A0(\s0.data_out[3][0] ),
    .A1(\s0.data_out[4][0] ),
    .S(net1067),
    .X(_2270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4796_ (.Y(_2271_),
    .A(net995),
    .B(_2270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4797_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2271_),
    .C1(net1458),
    .B1(_2269_),
    .A1(net1451),
    .Y(_2272_),
    .A2(_2265_));
 sg13g2_o21ai_1 _4798_ (.B1(_2258_),
    .VDD(VPWR),
    .Y(_2273_),
    .VSS(VGND),
    .A1(net1451),
    .A2(_2265_));
 sg13g2_nand2_1 _4799_ (.Y(_2274_),
    .A(net1056),
    .B(net574),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4800_ (.A0(\s0.data_out[4][3] ),
    .A1(\s0.data_out[3][3] ),
    .S(net1057),
    .X(_2275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4801_ (.A(net1050),
    .B_N(net1161),
    .Y(_2276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4802_ (.A2(_2275_),
    .A1(net1050),
    .B1(_2276_),
    .X(_2277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4803_ (.Y(_2278_),
    .B(\s0.data_out[3][3] ),
    .A_N(net1067),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4804_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2156_),
    .A2(_2278_),
    .Y(_2279_),
    .B1(net1060));
 sg13g2_a21oi_1 _4805_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1063),
    .A2(_2277_),
    .Y(_2280_),
    .B1(_2279_));
 sg13g2_a22oi_1 _4806_ (.Y(_2281_),
    .B1(_2280_),
    .B2(net1437),
    .A2(_2257_),
    .A1(net1444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4807_ (.B1(_2281_),
    .VDD(VPWR),
    .Y(_2282_),
    .VSS(VGND),
    .A1(_2272_),
    .A2(_2273_));
 sg13g2_nand2_1 _4808_ (.Y(_2283_),
    .A(net1058),
    .B(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4809_ (.A0(\s0.data_out[4][7] ),
    .A1(\s0.data_out[3][7] ),
    .S(net1059),
    .X(_2284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4810_ (.A(net1053),
    .B_N(net1143),
    .Y(_2285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4811_ (.A2(_2284_),
    .A1(net1053),
    .B1(_2285_),
    .X(_2286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4812_ (.Y(_2287_),
    .B(net484),
    .A_N(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4813_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2176_),
    .A2(_2287_),
    .Y(_2288_),
    .B1(net1064));
 sg13g2_a21oi_1 _4814_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1064),
    .A2(_2286_),
    .Y(_2289_),
    .B1(_2288_));
 sg13g2_nand2_1 _4815_ (.Y(_2290_),
    .A(net1058),
    .B(net678),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4816_ (.A0(\s0.data_out[4][6] ),
    .A1(\s0.data_out[3][6] ),
    .S(net1058),
    .X(_2291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4817_ (.A(net1053),
    .B_N(net1148),
    .Y(_2292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4818_ (.A2(_2291_),
    .A1(net1053),
    .B1(_2292_),
    .X(_2293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4819_ (.Y(_2294_),
    .B(\s0.data_out[3][6] ),
    .A_N(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4820_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2169_),
    .A2(_2294_),
    .Y(_2295_),
    .B1(net1064));
 sg13g2_a21oi_1 _4821_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1064),
    .A2(_2293_),
    .Y(_2296_),
    .B1(_2295_));
 sg13g2_a22oi_1 _4822_ (.Y(_2297_),
    .B1(_2296_),
    .B2(net1410),
    .A2(_2289_),
    .A1(net1401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4823_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2298_),
    .B(_2296_),
    .A(net1409));
 sg13g2_nor2_1 _4824_ (.A(net1401),
    .B(_2289_),
    .Y(_2299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4825_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2300_),
    .B(_2289_),
    .A(net1401));
 sg13g2_and3_1 _4826_ (.X(_2301_),
    .A(_2297_),
    .B(_2298_),
    .C(_2300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4827_ (.A(net1050),
    .B_N(net1157),
    .Y(_2302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4828_ (.Y(_2303_),
    .A(net1056),
    .B(net387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4829_ (.A0(\s0.data_out[4][4] ),
    .A1(\s0.data_out[3][4] ),
    .S(net1057),
    .X(_2304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4830_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1050),
    .A2(_2304_),
    .Y(_2305_),
    .B1(_2302_));
 sg13g2_nand2b_1 _4831_ (.Y(_2306_),
    .B(net1063),
    .A_N(_2305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4832_ (.B1(_2188_),
    .VDD(VPWR),
    .Y(_2307_),
    .VSS(VGND),
    .A1(net1067),
    .A2(_2876_));
 sg13g2_nand2_1 _4833_ (.Y(_2308_),
    .A(net996),
    .B(_2307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4834_ (.B(_2306_),
    .C(_2308_),
    .A(net1428),
    .Y(_2309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4835_ (.A(net1437),
    .B(_2280_),
    .Y(_2310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4836_ (.Y(_2311_),
    .A(net1058),
    .B(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4837_ (.A0(\s0.data_out[4][5] ),
    .A1(\s0.data_out[3][5] ),
    .S(net1059),
    .X(_2312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4838_ (.A(net1053),
    .B_N(net1152),
    .Y(_2313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4839_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1053),
    .A2(_2312_),
    .Y(_2314_),
    .B1(_2313_));
 sg13g2_nand2b_1 _4840_ (.Y(_2315_),
    .B(net1064),
    .A_N(_2314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4841_ (.B1(_2195_),
    .VDD(VPWR),
    .Y(_2316_),
    .VSS(VGND),
    .A1(net1069),
    .A2(_2875_));
 sg13g2_nand2_1 _4842_ (.Y(_2317_),
    .A(net996),
    .B(_2316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4843_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2315_),
    .A2(_2317_),
    .Y(_2318_),
    .B1(net1419));
 sg13g2_nand3_1 _4844_ (.B(_2315_),
    .C(_2317_),
    .A(net1419),
    .Y(_2319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4845_ (.A(_2318_),
    .B_N(_2319_),
    .Y(_2320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4846_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2306_),
    .A2(_2308_),
    .Y(_2321_),
    .B1(net1428));
 sg13g2_nor2_1 _4847_ (.A(_2310_),
    .B(_2321_),
    .Y(_2322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4848_ (.A(_2301_),
    .B(_2309_),
    .C(_2320_),
    .D(_2322_),
    .X(_2323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4849_ (.B1(_2319_),
    .VDD(VPWR),
    .Y(_2324_),
    .VSS(VGND),
    .A1(_2309_),
    .A2(_2318_));
 sg13g2_o21ai_1 _4850_ (.B1(_2245_),
    .VDD(VPWR),
    .Y(_2325_),
    .VSS(VGND),
    .A1(_2297_),
    .A2(_2299_));
 sg13g2_a221oi_1 _4851_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2301_),
    .C1(_2325_),
    .B1(_2324_),
    .A1(_2282_),
    .Y(_2326_),
    .A2(_2323_));
 sg13g2_nor3_1 _4852_ (.A(net321),
    .B(net1330),
    .C(_2326_),
    .Y(_0239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4853_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1049),
    .A2(net540),
    .Y(_2327_),
    .B1(_2267_));
 sg13g2_a21oi_1 _4854_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net995),
    .A2(_2270_),
    .Y(_2328_),
    .B1(net1358));
 sg13g2_o21ai_1 _4855_ (.B1(_2328_),
    .VDD(VPWR),
    .Y(_2329_),
    .VSS(VGND),
    .A1(net995),
    .A2(_2327_));
 sg13g2_o21ai_1 _4856_ (.B1(_2329_),
    .VDD(VPWR),
    .Y(_2330_),
    .VSS(VGND),
    .A1(net1473),
    .A2(net600));
 sg13g2_inv_1 _4857_ (.VDD(VPWR),
    .Y(_0240_),
    .A(_2330_),
    .VSS(VGND));
 sg13g2_and2_1 _4858_ (.A(net1049),
    .B(net400),
    .X(_2331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4859_ (.B1(net1060),
    .VDD(VPWR),
    .Y(_2332_),
    .VSS(VGND),
    .A1(_2261_),
    .A2(_2331_));
 sg13g2_nor2_1 _4860_ (.A(net1358),
    .B(_2264_),
    .Y(_2333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4861_ (.Y(_0241_),
    .B1(_2332_),
    .B2(_2333_),
    .A2(_2873_),
    .A1(net1359),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4862_ (.A(net1049),
    .B(net434),
    .X(_2334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4863_ (.B1(net1060),
    .VDD(VPWR),
    .Y(_2335_),
    .VSS(VGND),
    .A1(_2253_),
    .A2(_2334_));
 sg13g2_nor2_1 _4864_ (.A(net1359),
    .B(_2256_),
    .Y(_2336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4865_ (.Y(_0242_),
    .B1(_2335_),
    .B2(_2336_),
    .A2(_2872_),
    .A1(net1359),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4866_ (.A(net1050),
    .B(\s0.data_out[3][3] ),
    .X(_2337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4867_ (.B1(net1063),
    .VDD(VPWR),
    .Y(_2338_),
    .VSS(VGND),
    .A1(_2276_),
    .A2(_2337_));
 sg13g2_nor2_1 _4868_ (.A(net1358),
    .B(_2279_),
    .Y(_2339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4869_ (.Y(_0243_),
    .B1(_2338_),
    .B2(_2339_),
    .A2(_2871_),
    .A1(net1358),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4870_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1050),
    .A2(net387),
    .Y(_2340_),
    .B1(_2302_));
 sg13g2_a21oi_1 _4871_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net995),
    .A2(_2307_),
    .Y(_2341_),
    .B1(net1359));
 sg13g2_o21ai_1 _4872_ (.B1(_2341_),
    .VDD(VPWR),
    .Y(_2342_),
    .VSS(VGND),
    .A1(net995),
    .A2(_2340_));
 sg13g2_o21ai_1 _4873_ (.B1(_2342_),
    .VDD(VPWR),
    .Y(_2343_),
    .VSS(VGND),
    .A1(net1473),
    .A2(net569));
 sg13g2_inv_1 _4874_ (.VDD(VPWR),
    .Y(_0244_),
    .A(_2343_),
    .VSS(VGND));
 sg13g2_a21oi_1 _4875_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1053),
    .A2(net601),
    .Y(_2344_),
    .B1(_2313_));
 sg13g2_a21oi_1 _4876_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net996),
    .A2(_2316_),
    .Y(_2345_),
    .B1(net1361));
 sg13g2_o21ai_1 _4877_ (.B1(_2345_),
    .VDD(VPWR),
    .Y(_2346_),
    .VSS(VGND),
    .A1(net996),
    .A2(_2344_));
 sg13g2_o21ai_1 _4878_ (.B1(_2346_),
    .VDD(VPWR),
    .Y(_2347_),
    .VSS(VGND),
    .A1(net1473),
    .A2(net681));
 sg13g2_inv_1 _4879_ (.VDD(VPWR),
    .Y(_0245_),
    .A(_2347_),
    .VSS(VGND));
 sg13g2_and2_1 _4880_ (.A(net1054),
    .B(\s0.data_out[3][6] ),
    .X(_2348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4881_ (.B1(net1064),
    .VDD(VPWR),
    .Y(_2349_),
    .VSS(VGND),
    .A1(_2292_),
    .A2(_2348_));
 sg13g2_nor2_1 _4882_ (.A(net1361),
    .B(_2295_),
    .Y(_2350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4883_ (.Y(_0246_),
    .B1(_2349_),
    .B2(_2350_),
    .A2(_2870_),
    .A1(net1360),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4884_ (.A(net1053),
    .B(net484),
    .X(_2351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4885_ (.B1(net1066),
    .VDD(VPWR),
    .Y(_2352_),
    .VSS(VGND),
    .A1(_2285_),
    .A2(_2351_));
 sg13g2_nor2_1 _4886_ (.A(net1360),
    .B(_2288_),
    .Y(_2353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4887_ (.Y(_0247_),
    .B1(_2352_),
    .B2(_2353_),
    .A2(_2869_),
    .A1(net1361),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4888_ (.B1(net1052),
    .VDD(VPWR),
    .Y(_2354_),
    .VSS(VGND),
    .A1(net1397),
    .A2(net1040));
 sg13g2_nand2_1 _4889_ (.Y(_2355_),
    .A(net1336),
    .B(net1046),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4890_ (.Y(_2356_),
    .B(_2355_),
    .A_N(_2354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4891_ (.B1(_2356_),
    .VDD(VPWR),
    .Y(_2357_),
    .VSS(VGND),
    .A1(net1051),
    .A2(_2242_));
 sg13g2_nor2_1 _4892_ (.A(net356),
    .B(net1045),
    .Y(_2358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4893_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2359_),
    .B(_2358_),
    .A(_2356_));
 sg13g2_nor2_1 _4894_ (.A(net1040),
    .B(_2354_),
    .Y(_2360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4895_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2729_),
    .A2(_2748_),
    .Y(_2361_),
    .B1(net1051));
 sg13g2_nor2_1 _4896_ (.A(_2360_),
    .B(_2361_),
    .Y(_2362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4897_ (.B1(net1473),
    .VDD(VPWR),
    .Y(_2363_),
    .VSS(VGND),
    .A1(net524),
    .A2(_2357_));
 sg13g2_a21oi_1 _4898_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2359_),
    .A2(_2362_),
    .Y(_0248_),
    .B1(_2363_));
 sg13g2_nor2_1 _4899_ (.A(net1360),
    .B(_2357_),
    .Y(_0249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4900_ (.A(net1468),
    .B(net334),
    .X(_0250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4901_ (.A0(\s0.data_out[3][2] ),
    .A1(\s0.data_out[2][2] ),
    .S(net1043),
    .X(_2364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4902_ (.A(net1036),
    .B_N(net1163),
    .Y(_2365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4903_ (.A2(_2364_),
    .A1(net1036),
    .B1(_2365_),
    .X(_2366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4904_ (.Y(_2367_),
    .B(\s0.data_out[2][2] ),
    .A_N(net1056),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4905_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2251_),
    .A2(_2367_),
    .Y(_2368_),
    .B1(net1047));
 sg13g2_a21oi_1 _4906_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1048),
    .A2(_2366_),
    .Y(_2369_),
    .B1(_2368_));
 sg13g2_nor2_1 _4907_ (.A(net1444),
    .B(_2369_),
    .Y(_2370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4908_ (.Y(_2371_),
    .A(net1043),
    .B(net514),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4909_ (.A0(\s0.data_out[3][1] ),
    .A1(\s0.data_out[2][1] ),
    .S(net1044),
    .X(_2372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4910_ (.A(net1036),
    .B_N(net1167),
    .Y(_2373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4911_ (.A2(_2372_),
    .A1(net1036),
    .B1(_2373_),
    .X(_2374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4912_ (.Y(_2375_),
    .B(\s0.data_out[2][1] ),
    .A_N(net1056),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4913_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2259_),
    .A2(_2375_),
    .Y(_2376_),
    .B1(net1047));
 sg13g2_a21oi_1 _4914_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1047),
    .A2(_2374_),
    .Y(_2377_),
    .B1(_2376_));
 sg13g2_mux2_1 _4915_ (.A0(\s0.data_out[3][0] ),
    .A1(\s0.data_out[2][0] ),
    .S(net1043),
    .X(_2378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4916_ (.A(net1036),
    .B_N(net1173),
    .Y(_2379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4917_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1036),
    .A2(_2378_),
    .Y(_2380_),
    .B1(_2379_));
 sg13g2_nand2b_1 _4918_ (.Y(_2381_),
    .B(net1047),
    .A_N(_2380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4919_ (.A0(\s0.data_out[2][0] ),
    .A1(\s0.data_out[3][0] ),
    .S(net1056),
    .X(_2382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4920_ (.Y(_2383_),
    .B(_2382_),
    .A_N(net1047),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4921_ (.A(net1457),
    .B(_2377_),
    .Y(_2384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4922_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2383_),
    .C1(net1461),
    .B1(_2381_),
    .A1(net1457),
    .Y(_2385_),
    .A2(_2377_));
 sg13g2_nor3_1 _4923_ (.A(_2370_),
    .B(_2384_),
    .C(_2385_),
    .Y(_2386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4924_ (.Y(_2387_),
    .A(net1044),
    .B(net463),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4925_ (.B1(_2387_),
    .VDD(VPWR),
    .Y(_2388_),
    .VSS(VGND),
    .A1(net1044),
    .A2(_2877_));
 sg13g2_nor2_1 _4926_ (.A(net1037),
    .B(net993),
    .Y(_2389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4927_ (.A2(_2388_),
    .A1(net1037),
    .B1(_2389_),
    .X(_2390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4928_ (.Y(_2391_),
    .A(_2748_),
    .B(net463),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4929_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2274_),
    .A2(_2391_),
    .Y(_2392_),
    .B1(net1048));
 sg13g2_a21oi_1 _4930_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1048),
    .A2(_2390_),
    .Y(_2393_),
    .B1(_2392_));
 sg13g2_a221oi_1 _4931_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net1438),
    .C1(_2386_),
    .B1(_2393_),
    .A1(net1444),
    .Y(_2394_),
    .A2(_2369_));
 sg13g2_nand2_1 _4932_ (.Y(_2395_),
    .A(net1045),
    .B(net512),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4933_ (.A0(\s0.data_out[3][7] ),
    .A1(\s0.data_out[2][7] ),
    .S(net1046),
    .X(_2396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4934_ (.A(net1040),
    .B_N(net1142),
    .Y(_2397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4935_ (.A2(_2396_),
    .A1(net1040),
    .B1(_2397_),
    .X(_2398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4936_ (.Y(_2399_),
    .B(\s0.data_out[2][7] ),
    .A_N(net1058),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4937_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2283_),
    .A2(_2399_),
    .Y(_2400_),
    .B1(net1051));
 sg13g2_a21oi_1 _4938_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1051),
    .A2(_2398_),
    .Y(_2401_),
    .B1(_2400_));
 sg13g2_nand2_1 _4939_ (.Y(_2402_),
    .A(net1045),
    .B(net580),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4940_ (.A0(\s0.data_out[3][6] ),
    .A1(\s0.data_out[2][6] ),
    .S(net1046),
    .X(_2403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4941_ (.A(net1040),
    .B_N(net1147),
    .Y(_2404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4942_ (.A2(_2403_),
    .A1(net1041),
    .B1(_2404_),
    .X(_2405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4943_ (.Y(_2406_),
    .B(net580),
    .A_N(net1058),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4944_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2290_),
    .A2(_2406_),
    .Y(_2407_),
    .B1(net1052));
 sg13g2_a21oi_1 _4945_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1052),
    .A2(_2405_),
    .Y(_2408_),
    .B1(_2407_));
 sg13g2_a22oi_1 _4946_ (.Y(_2409_),
    .B1(_2408_),
    .B2(net1409),
    .A2(_2401_),
    .A1(net1400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4947_ (.A(net1409),
    .B(_2408_),
    .Y(_2410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4948_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2411_),
    .B(_2401_),
    .A(net1400));
 sg13g2_nand3b_1 _4949_ (.B(_2411_),
    .C(_2409_),
    .Y(_2412_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2410_));
 sg13g2_mux2_1 _4950_ (.A0(\s0.data_out[3][5] ),
    .A1(\s0.data_out[2][5] ),
    .S(net1045),
    .X(_2413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4951_ (.A(net1040),
    .B_N(net1152),
    .Y(_2414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4952_ (.A2(_2413_),
    .A1(net1040),
    .B1(_2414_),
    .X(_2415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4953_ (.Y(_2416_),
    .B(net576),
    .A_N(net1058),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4954_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2311_),
    .A2(_2416_),
    .Y(_2417_),
    .B1(net1051));
 sg13g2_a21oi_1 _4955_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1051),
    .A2(_2415_),
    .Y(_2418_),
    .B1(_2417_));
 sg13g2_nand2_1 _4956_ (.Y(_2419_),
    .A(net1419),
    .B(_2418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4957_ (.B1(_2419_),
    .VDD(VPWR),
    .Y(_2420_),
    .VSS(VGND),
    .A1(net1438),
    .A2(_2393_));
 sg13g2_nor2_1 _4958_ (.A(net1419),
    .B(_2418_),
    .Y(_2421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4959_ (.A0(\s0.data_out[3][4] ),
    .A1(\s0.data_out[2][4] ),
    .S(net1044),
    .X(_2422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4960_ (.A(net1037),
    .B_N(net1157),
    .Y(_2423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4961_ (.A2(_2422_),
    .A1(net1037),
    .B1(_2423_),
    .X(_2424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4962_ (.Y(_2425_),
    .B(\s0.data_out[2][4] ),
    .A_N(net1056),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4963_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2303_),
    .A2(_2425_),
    .Y(_2426_),
    .B1(net1048));
 sg13g2_a21oi_1 _4964_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1051),
    .A2(_2424_),
    .Y(_2427_),
    .B1(_2426_));
 sg13g2_nand2_1 _4965_ (.Y(_2428_),
    .A(net1428),
    .B(_2427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4966_ (.A(_2421_),
    .B_N(_2428_),
    .Y(_2429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4967_ (.B1(_2429_),
    .VDD(VPWR),
    .Y(_2430_),
    .VSS(VGND),
    .A1(net1428),
    .A2(_2427_));
 sg13g2_or4_1 _4968_ (.A(_2394_),
    .B(_2412_),
    .C(_2420_),
    .D(_2430_),
    .X(_2431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4969_ (.B1(_2419_),
    .VDD(VPWR),
    .Y(_2432_),
    .VSS(VGND),
    .A1(_2421_),
    .A2(_2428_));
 sg13g2_nor2b_1 _4970_ (.A(_2412_),
    .B_N(_2432_),
    .Y(_2433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4971_ (.A(_2409_),
    .B_N(_2411_),
    .Y(_2434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4972_ (.A(_2357_),
    .B(_2433_),
    .C(_2434_),
    .Y(_2435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4973_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2436_),
    .B(net1330),
    .A(net340));
 sg13g2_a21oi_1 _4974_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2431_),
    .A2(_2435_),
    .Y(_0251_),
    .B1(_2436_));
 sg13g2_and2_1 _4975_ (.A(net1036),
    .B(\s0.data_out[2][0] ),
    .X(_2437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4976_ (.B1(net1047),
    .VDD(VPWR),
    .Y(_2438_),
    .VSS(VGND),
    .A1(_2379_),
    .A2(_2437_));
 sg13g2_nand3_1 _4977_ (.B(_2383_),
    .C(_2438_),
    .A(net1473),
    .Y(_2439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4978_ (.B1(_2439_),
    .VDD(VPWR),
    .Y(_2440_),
    .VSS(VGND),
    .A1(net1473),
    .A2(net540));
 sg13g2_inv_1 _4979_ (.VDD(VPWR),
    .Y(_0252_),
    .A(_2440_),
    .VSS(VGND));
 sg13g2_nor2_1 _4980_ (.A(net1009),
    .B(_2883_),
    .Y(_2441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4981_ (.B1(net1047),
    .VDD(VPWR),
    .Y(_2442_),
    .VSS(VGND),
    .A1(_2373_),
    .A2(_2441_));
 sg13g2_nor2_1 _4982_ (.A(net1358),
    .B(_2376_),
    .Y(_2443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4983_ (.Y(_0253_),
    .B1(_2442_),
    .B2(_2443_),
    .A2(_2879_),
    .A1(net1358),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4984_ (.A(net1036),
    .B(\s0.data_out[2][2] ),
    .X(_2444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4985_ (.B1(net1047),
    .VDD(VPWR),
    .Y(_2445_),
    .VSS(VGND),
    .A1(_2365_),
    .A2(_2444_));
 sg13g2_nor2_1 _4986_ (.A(net1358),
    .B(_2368_),
    .Y(_2446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4987_ (.Y(_0254_),
    .B1(_2445_),
    .B2(_2446_),
    .A2(_2878_),
    .A1(net1358),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4988_ (.A(net1009),
    .B(_2882_),
    .Y(_2447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4989_ (.B1(net1048),
    .VDD(VPWR),
    .Y(_2448_),
    .VSS(VGND),
    .A1(_2389_),
    .A2(_2447_));
 sg13g2_nor2_1 _4990_ (.A(net1348),
    .B(_2392_),
    .Y(_2449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4991_ (.Y(_0255_),
    .B1(_2448_),
    .B2(_2449_),
    .A2(_2877_),
    .A1(net1348),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4992_ (.A(net1037),
    .B(net583),
    .X(_2450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4993_ (.B1(net1048),
    .VDD(VPWR),
    .Y(_2451_),
    .VSS(VGND),
    .A1(_2423_),
    .A2(_2450_));
 sg13g2_nor2_1 _4994_ (.A(net1360),
    .B(net388),
    .Y(_2452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4995_ (.Y(_0256_),
    .B1(_2451_),
    .B2(_2452_),
    .A2(_2876_),
    .A1(net1360),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4996_ (.A(net1040),
    .B(net576),
    .X(_2453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4997_ (.B1(net1051),
    .VDD(VPWR),
    .Y(_2454_),
    .VSS(VGND),
    .A1(_2414_),
    .A2(_2453_));
 sg13g2_nor2_1 _4998_ (.A(net1360),
    .B(_2417_),
    .Y(_2455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4999_ (.Y(_0257_),
    .B1(_2454_),
    .B2(_2455_),
    .A2(_2875_),
    .A1(net1360),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5000_ (.A(net1010),
    .B(_2881_),
    .Y(_2456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5001_ (.B1(net1052),
    .VDD(VPWR),
    .Y(_2457_),
    .VSS(VGND),
    .A1(_2404_),
    .A2(_2456_));
 sg13g2_nand3b_1 _5002_ (.B(_2457_),
    .C(net1475),
    .Y(_2458_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2407_));
 sg13g2_o21ai_1 _5003_ (.B1(_2458_),
    .VDD(VPWR),
    .Y(_2459_),
    .VSS(VGND),
    .A1(net1475),
    .A2(net678));
 sg13g2_inv_1 _5004_ (.VDD(VPWR),
    .Y(_0258_),
    .A(_2459_),
    .VSS(VGND));
 sg13g2_nor2_1 _5005_ (.A(net1010),
    .B(_2880_),
    .Y(_2460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5006_ (.B1(net1052),
    .VDD(VPWR),
    .Y(_2461_),
    .VSS(VGND),
    .A1(_2397_),
    .A2(_2460_));
 sg13g2_nor2_1 _5007_ (.A(net1360),
    .B(_2400_),
    .Y(_2462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5008_ (.Y(_0259_),
    .B1(_2461_),
    .B2(_2462_),
    .A2(_2874_),
    .A1(net1348),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5009_ (.B1(net1039),
    .VDD(VPWR),
    .Y(_2463_),
    .VSS(VGND),
    .A1(net1392),
    .A2(net1030));
 sg13g2_nor2b_1 _5010_ (.A(net1392),
    .B_N(net1034),
    .Y(_2464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5011_ (.A(_2463_),
    .B(_2464_),
    .Y(_2465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5012_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1010),
    .A2(_2355_),
    .Y(_2466_),
    .B1(_2465_));
 sg13g2_o21ai_1 _5013_ (.B1(_2465_),
    .VDD(VPWR),
    .Y(_2467_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[1] [0]),
    .A2(net1034));
 sg13g2_nor2_1 _5014_ (.A(net1030),
    .B(_2463_),
    .Y(_2468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5015_ (.B1(net1010),
    .VDD(VPWR),
    .Y(_2469_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[1] [0]),
    .A2(net1045));
 sg13g2_nand2_1 _5016_ (.Y(_2470_),
    .A(_2467_),
    .B(_2469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5017_ (.B1(net1468),
    .VDD(VPWR),
    .Y(_2471_),
    .VSS(VGND),
    .A1(_2468_),
    .A2(_2470_));
 sg13g2_a21oi_1 _5018_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2729_),
    .A2(_2466_),
    .Y(_0260_),
    .B1(_2471_));
 sg13g2_and2_1 _5019_ (.A(net1469),
    .B(_2466_),
    .X(_0261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5020_ (.A(net1463),
    .B(net335),
    .X(_0262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5021_ (.Y(_2472_),
    .A(net1033),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5022_ (.A0(\s0.data_out[2][1] ),
    .A1(\s0.data_out[1][1] ),
    .S(net1033),
    .X(_2473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5023_ (.A(net1027),
    .B_N(net1166),
    .Y(_2474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5024_ (.A2(_2473_),
    .A1(net1027),
    .B1(_2474_),
    .X(_2475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5025_ (.Y(_2476_),
    .B(net494),
    .A_N(net1043),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5026_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2371_),
    .A2(_2476_),
    .Y(_2477_),
    .B1(net1038));
 sg13g2_a21oi_1 _5027_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1038),
    .A2(_2475_),
    .Y(_2478_),
    .B1(_2477_));
 sg13g2_mux2_1 _5028_ (.A0(\s0.data_out[1][0] ),
    .A1(\s0.data_out[2][0] ),
    .S(net1043),
    .X(_2479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5029_ (.Y(_2480_),
    .A(net1009),
    .B(_2479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5030_ (.A(net1027),
    .B_N(net1170),
    .Y(_2481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5031_ (.A0(\s0.data_out[2][0] ),
    .A1(\s0.data_out[1][0] ),
    .S(net1035),
    .X(_2482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5032_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1027),
    .A2(_2482_),
    .Y(_2483_),
    .B1(_2481_));
 sg13g2_nand2b_1 _5033_ (.Y(_2484_),
    .B(net1038),
    .A_N(_2483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5034_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2484_),
    .C1(net1458),
    .B1(_2480_),
    .A1(net1450),
    .Y(_2485_),
    .A2(_2478_));
 sg13g2_mux2_1 _5035_ (.A0(\s0.data_out[2][2] ),
    .A1(\s0.data_out[1][2] ),
    .S(net1033),
    .X(_2486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5036_ (.A(net1027),
    .B_N(net1162),
    .Y(_2487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5037_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1027),
    .A2(_2486_),
    .Y(_2488_),
    .B1(_2487_));
 sg13g2_mux2_1 _5038_ (.A0(\s0.data_out[1][2] ),
    .A1(\s0.data_out[2][2] ),
    .S(net1043),
    .X(_2489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5039_ (.Y(_2490_),
    .A(net1009),
    .B(_2489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5040_ (.B1(_2490_),
    .VDD(VPWR),
    .Y(_2491_),
    .VSS(VGND),
    .A1(net1009),
    .A2(_2488_));
 sg13g2_or2_1 _5041_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2492_),
    .B(_2491_),
    .A(net1334));
 sg13g2_xnor2_1 _5042_ (.Y(_2493_),
    .A(net1334),
    .B(_2491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5043_ (.A0(\s0.data_out[2][3] ),
    .A1(\s0.data_out[1][3] ),
    .S(net1035),
    .X(_2494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5044_ (.A(net1028),
    .B_N(net1161),
    .Y(_2495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5045_ (.A2(_2494_),
    .A1(net1028),
    .B1(_2495_),
    .X(_2496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5046_ (.Y(_2497_),
    .B(\s0.data_out[1][3] ),
    .A_N(net1043),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5047_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2387_),
    .A2(_2497_),
    .Y(_2498_),
    .B1(net1038));
 sg13g2_a21oi_1 _5048_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1038),
    .A2(_2496_),
    .Y(_2499_),
    .B1(_2498_));
 sg13g2_nor2_1 _5049_ (.A(net1435),
    .B(_2499_),
    .Y(_2500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5050_ (.A(net1450),
    .B(_2478_),
    .Y(_2501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _5051_ (.A(_2485_),
    .B(_2493_),
    .C(_2500_),
    .D(_2501_),
    .Y(_2502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5052_ (.Y(_2503_),
    .A(net1436),
    .B(_2499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5053_ (.B1(_2503_),
    .VDD(VPWR),
    .Y(_2504_),
    .VSS(VGND),
    .A1(_2492_),
    .A2(_2500_));
 sg13g2_nor2_1 _5054_ (.A(_2502_),
    .B(_2504_),
    .Y(_2505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5055_ (.A0(\s0.data_out[2][7] ),
    .A1(\s0.data_out[1][7] ),
    .S(net1034),
    .X(_2506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5056_ (.A(net1030),
    .B_N(net1142),
    .Y(_2507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5057_ (.A2(_2506_),
    .A1(net1030),
    .B1(_2507_),
    .X(_2508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5058_ (.Y(_2509_),
    .B(\s0.data_out[1][7] ),
    .A_N(net1045),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5059_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2395_),
    .A2(_2509_),
    .Y(_2510_),
    .B1(net1039));
 sg13g2_a21oi_1 _5060_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1039),
    .A2(_2508_),
    .Y(_2511_),
    .B1(_2510_));
 sg13g2_mux2_1 _5061_ (.A0(\s0.data_out[2][6] ),
    .A1(\s0.data_out[1][6] ),
    .S(net1034),
    .X(_2512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5062_ (.A(net1032),
    .B_N(net1147),
    .Y(_2513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5063_ (.A2(_2512_),
    .A1(net1030),
    .B1(_2513_),
    .X(_2514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5064_ (.Y(_2515_),
    .B(\s0.data_out[1][6] ),
    .A_N(net1045),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5065_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2402_),
    .A2(_2515_),
    .Y(_2516_),
    .B1(net1039));
 sg13g2_a21oi_1 _5066_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1039),
    .A2(_2514_),
    .Y(_2517_),
    .B1(_2516_));
 sg13g2_a22oi_1 _5067_ (.Y(_2518_),
    .B1(_2517_),
    .B2(net1408),
    .A2(_2511_),
    .A1(net1399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5068_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2519_),
    .B(_2517_),
    .A(net1408));
 sg13g2_nor2_1 _5069_ (.A(net1399),
    .B(_2511_),
    .Y(_2520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _5070_ (.B(_2518_),
    .C(_2519_),
    .Y(_2521_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2520_));
 sg13g2_nor2b_1 _5071_ (.A(net1028),
    .B_N(net1156),
    .Y(_2522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5072_ (.A0(\s0.data_out[2][4] ),
    .A1(\s0.data_out[1][4] ),
    .S(net1035),
    .X(_2523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5073_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1028),
    .A2(_2523_),
    .Y(_2524_),
    .B1(_2522_));
 sg13g2_nand2b_1 _5074_ (.Y(_2525_),
    .B(net1039),
    .A_N(_2524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5075_ (.A0(\s0.data_out[1][4] ),
    .A1(\s0.data_out[2][4] ),
    .S(net1043),
    .X(_2526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5076_ (.Y(_2527_),
    .A(_2751_),
    .B(_2526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5077_ (.B(_2525_),
    .C(_2527_),
    .A(net1426),
    .Y(_2528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5078_ (.A0(\s0.data_out[2][5] ),
    .A1(\s0.data_out[1][5] ),
    .S(net1035),
    .X(_2529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5079_ (.A(net1030),
    .B_N(net1151),
    .Y(_2530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5080_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1030),
    .A2(_2529_),
    .Y(_2531_),
    .B1(_2530_));
 sg13g2_nand2b_1 _5081_ (.Y(_2532_),
    .B(net1039),
    .A_N(_2531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5082_ (.A0(\s0.data_out[1][5] ),
    .A1(\s0.data_out[2][5] ),
    .S(net1045),
    .X(_2533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5083_ (.Y(_2534_),
    .A(_2751_),
    .B(_2533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5084_ (.B(_2532_),
    .C(_2534_),
    .A(net1417),
    .Y(_2535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5085_ (.Y(_2536_),
    .A(_2528_),
    .B(_2535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5086_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2525_),
    .A2(_2527_),
    .Y(_2537_),
    .B1(net1429));
 sg13g2_a21oi_1 _5087_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2532_),
    .A2(_2534_),
    .Y(_2538_),
    .B1(net1417));
 sg13g2_or2_1 _5088_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2539_),
    .B(_2538_),
    .A(_2537_));
 sg13g2_or4_1 _5089_ (.A(_2505_),
    .B(_2521_),
    .C(_2536_),
    .D(_2539_),
    .X(_2540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5090_ (.B1(_2535_),
    .VDD(VPWR),
    .Y(_2541_),
    .VSS(VGND),
    .A1(_2528_),
    .A2(_2538_));
 sg13g2_nor2b_1 _5091_ (.A(_2521_),
    .B_N(_2541_),
    .Y(_2542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5092_ (.B1(_2466_),
    .VDD(VPWR),
    .Y(_2543_),
    .VSS(VGND),
    .A1(_2518_),
    .A2(_2520_));
 sg13g2_nor2_1 _5093_ (.A(_2542_),
    .B(_2543_),
    .Y(_2544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5094_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2545_),
    .B(net1329),
    .A(net334));
 sg13g2_a21oi_1 _5095_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2540_),
    .A2(_2544_),
    .Y(_0263_),
    .B1(_2545_));
 sg13g2_a21oi_1 _5096_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1027),
    .A2(net652),
    .Y(_2546_),
    .B1(_2481_));
 sg13g2_a21oi_1 _5097_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1009),
    .A2(_2479_),
    .Y(_2547_),
    .B1(net1348));
 sg13g2_o21ai_1 _5098_ (.B1(_2547_),
    .VDD(VPWR),
    .Y(_2548_),
    .VSS(VGND),
    .A1(net1009),
    .A2(_2546_));
 sg13g2_o21ai_1 _5099_ (.B1(_2548_),
    .VDD(VPWR),
    .Y(_2549_),
    .VSS(VGND),
    .A1(net1468),
    .A2(net663));
 sg13g2_inv_1 _5100_ (.VDD(VPWR),
    .Y(_0264_),
    .A(_2549_),
    .VSS(VGND));
 sg13g2_nor2_1 _5101_ (.A(net1004),
    .B(_2884_),
    .Y(_2550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5102_ (.B1(net1038),
    .VDD(VPWR),
    .Y(_2551_),
    .VSS(VGND),
    .A1(_2474_),
    .A2(_2550_));
 sg13g2_nor2_1 _5103_ (.A(net1348),
    .B(_2477_),
    .Y(_2552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5104_ (.Y(_0265_),
    .B1(_2551_),
    .B2(_2552_),
    .A2(_2883_),
    .A1(net1348),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5105_ (.A(net1027),
    .B(\s0.data_out[1][2] ),
    .X(_2553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5106_ (.B1(net1038),
    .VDD(VPWR),
    .Y(_2554_),
    .VSS(VGND),
    .A1(_2487_),
    .A2(_2553_));
 sg13g2_nand3_1 _5107_ (.B(_2490_),
    .C(_2554_),
    .A(net1468),
    .Y(_2555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5108_ (.B1(_2555_),
    .VDD(VPWR),
    .Y(_2556_),
    .VSS(VGND),
    .A1(net1468),
    .A2(net582));
 sg13g2_inv_1 _5109_ (.VDD(VPWR),
    .Y(_0266_),
    .A(_2556_),
    .VSS(VGND));
 sg13g2_and2_1 _5110_ (.A(net1028),
    .B(\s0.data_out[1][3] ),
    .X(_2557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5111_ (.B1(net1038),
    .VDD(VPWR),
    .Y(_2558_),
    .VSS(VGND),
    .A1(_2495_),
    .A2(_2557_));
 sg13g2_nor2_1 _5112_ (.A(net1348),
    .B(_2498_),
    .Y(_2559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5113_ (.Y(_0267_),
    .B1(_2558_),
    .B2(_2559_),
    .A2(_2882_),
    .A1(net1348),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5114_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1028),
    .A2(\s0.data_out[1][4] ),
    .Y(_2560_),
    .B1(_2522_));
 sg13g2_a21oi_1 _5115_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1009),
    .A2(_2526_),
    .Y(_2561_),
    .B1(net1349));
 sg13g2_o21ai_1 _5116_ (.B1(_2561_),
    .VDD(VPWR),
    .Y(_2562_),
    .VSS(VGND),
    .A1(net1010),
    .A2(_2560_));
 sg13g2_o21ai_1 _5117_ (.B1(_2562_),
    .VDD(VPWR),
    .Y(_2563_),
    .VSS(VGND),
    .A1(net1468),
    .A2(net583));
 sg13g2_inv_1 _5118_ (.VDD(VPWR),
    .Y(_0268_),
    .A(net584),
    .VSS(VGND));
 sg13g2_a21oi_1 _5119_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1030),
    .A2(\s0.data_out[1][5] ),
    .Y(_2564_),
    .B1(_2530_));
 sg13g2_a21oi_1 _5120_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1010),
    .A2(_2533_),
    .Y(_2565_),
    .B1(net1349));
 sg13g2_o21ai_1 _5121_ (.B1(_2565_),
    .VDD(VPWR),
    .Y(_2566_),
    .VSS(VGND),
    .A1(net1010),
    .A2(_2564_));
 sg13g2_o21ai_1 _5122_ (.B1(_2566_),
    .VDD(VPWR),
    .Y(_2567_),
    .VSS(VGND),
    .A1(net1468),
    .A2(net576));
 sg13g2_inv_1 _5123_ (.VDD(VPWR),
    .Y(_0269_),
    .A(net577),
    .VSS(VGND));
 sg13g2_and2_1 _5124_ (.A(net1032),
    .B(\s0.data_out[1][6] ),
    .X(_2568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5125_ (.B1(net1041),
    .VDD(VPWR),
    .Y(_2569_),
    .VSS(VGND),
    .A1(_2513_),
    .A2(_2568_));
 sg13g2_nor2_1 _5126_ (.A(net1349),
    .B(_2516_),
    .Y(_2570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5127_ (.Y(_0270_),
    .B1(_2569_),
    .B2(_2570_),
    .A2(_2881_),
    .A1(net1349),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5128_ (.A(net1032),
    .B(\s0.data_out[1][7] ),
    .X(_2571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5129_ (.B1(net1041),
    .VDD(VPWR),
    .Y(_2572_),
    .VSS(VGND),
    .A1(_2507_),
    .A2(_2571_));
 sg13g2_nor2_1 _5130_ (.A(net1349),
    .B(_2510_),
    .Y(_2573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5131_ (.Y(_0271_),
    .B1(_2572_),
    .B2(_2573_),
    .A2(_2880_),
    .A1(net1349),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5132_ (.B1(net1031),
    .VDD(VPWR),
    .Y(_2574_),
    .VSS(VGND),
    .A1(net1392),
    .A2(net1022));
 sg13g2_a21oi_1 _5133_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1336),
    .A2(net1025),
    .Y(_2575_),
    .B1(_2574_));
 sg13g2_inv_1 _5134_ (.VDD(VPWR),
    .Y(_2576_),
    .A(_2575_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5135_ (.B1(_2576_),
    .VDD(VPWR),
    .Y(_2577_),
    .VSS(VGND),
    .A1(net1031),
    .A2(_2464_));
 sg13g2_or2_1 _5136_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2578_),
    .B(net1026),
    .A(net427));
 sg13g2_o21ai_1 _5137_ (.B1(net1006),
    .VDD(VPWR),
    .Y(_2579_),
    .VSS(VGND),
    .A1(net427),
    .A2(net1034));
 sg13g2_o21ai_1 _5138_ (.B1(_2579_),
    .VDD(VPWR),
    .Y(_2580_),
    .VSS(VGND),
    .A1(net1022),
    .A2(_2574_));
 sg13g2_a21oi_1 _5139_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2575_),
    .A2(_2578_),
    .Y(_2581_),
    .B1(_2580_));
 sg13g2_o21ai_1 _5140_ (.B1(net1468),
    .VDD(VPWR),
    .Y(_2582_),
    .VSS(VGND),
    .A1(net516),
    .A2(_2577_));
 sg13g2_nor2_1 _5141_ (.A(_2581_),
    .B(_2582_),
    .Y(_0272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5142_ (.A(net1346),
    .B(_2577_),
    .Y(_0273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5143_ (.A(net1471),
    .B(net327),
    .X(_0274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5144_ (.A0(\s0.data_out[0][2] ),
    .A1(\s0.data_out[1][2] ),
    .S(net1033),
    .X(_2583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5145_ (.A0(\s0.data_out[1][2] ),
    .A1(\s0.data_out[0][2] ),
    .S(net1024),
    .X(_2584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5146_ (.A(net1019),
    .B_N(net1162),
    .Y(_2585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5147_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1020),
    .A2(_2584_),
    .Y(_2586_),
    .B1(_2585_));
 sg13g2_nor2_1 _5148_ (.A(net1004),
    .B(_2586_),
    .Y(_2587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5149_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1004),
    .A2(_2583_),
    .Y(_2588_),
    .B1(_2587_));
 sg13g2_nand2b_1 _5150_ (.Y(_2589_),
    .B(net375),
    .A_N(net1033),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5151_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2472_),
    .A2(_2589_),
    .Y(_2590_),
    .B1(net1029));
 sg13g2_mux2_1 _5152_ (.A0(\s0.data_out[1][1] ),
    .A1(\s0.data_out[0][1] ),
    .S(net1026),
    .X(_2591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5153_ (.A(net1020),
    .B_N(net1166),
    .Y(_2592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5154_ (.A2(_2591_),
    .A1(net1020),
    .B1(_2592_),
    .X(_2593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5155_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1029),
    .A2(_2593_),
    .Y(_2594_),
    .B1(_2590_));
 sg13g2_mux2_1 _5156_ (.A0(\s0.data_out[0][0] ),
    .A1(\s0.data_out[1][0] ),
    .S(net1033),
    .X(_2595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5157_ (.Y(_2596_),
    .A(net1004),
    .B(_2595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5158_ (.A0(\s0.data_out[1][0] ),
    .A1(\s0.data_out[0][0] ),
    .S(net1026),
    .X(_2597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5159_ (.A(net1020),
    .B_N(net1170),
    .Y(_2598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5160_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1020),
    .A2(_2597_),
    .Y(_2599_),
    .B1(_2598_));
 sg13g2_nand2b_1 _5161_ (.Y(_2600_),
    .B(net1029),
    .A_N(_2599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5162_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2601_),
    .B(_2594_),
    .A(net1450));
 sg13g2_a221oi_1 _5163_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2600_),
    .C1(net1458),
    .B1(_2596_),
    .A1(net1449),
    .Y(_2602_),
    .A2(_2594_));
 sg13g2_o21ai_1 _5164_ (.B1(_2601_),
    .VDD(VPWR),
    .Y(_2603_),
    .VSS(VGND),
    .A1(net1443),
    .A2(_2588_));
 sg13g2_mux2_1 _5165_ (.A0(\s0.data_out[0][3] ),
    .A1(\s0.data_out[1][3] ),
    .S(net1033),
    .X(_2604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5166_ (.A0(\s0.data_out[1][3] ),
    .A1(\s0.data_out[0][3] ),
    .S(net1024),
    .X(_2605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5167_ (.A(net1020),
    .B_N(net1161),
    .Y(_2606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5168_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1021),
    .A2(_2605_),
    .Y(_2607_),
    .B1(_2606_));
 sg13g2_nor2_1 _5169_ (.A(net1005),
    .B(_2607_),
    .Y(_2608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5170_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1005),
    .A2(_2604_),
    .Y(_2609_),
    .B1(_2608_));
 sg13g2_a22oi_1 _5171_ (.Y(_2610_),
    .B1(_2609_),
    .B2(net1436),
    .A2(_2588_),
    .A1(net1443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5172_ (.B1(_2610_),
    .VDD(VPWR),
    .Y(_2611_),
    .VSS(VGND),
    .A1(_2602_),
    .A2(_2603_));
 sg13g2_mux2_1 _5173_ (.A0(\s0.data_out[0][7] ),
    .A1(\s0.data_out[1][7] ),
    .S(net1034),
    .X(_2612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5174_ (.A0(\s0.data_out[1][7] ),
    .A1(\s0.data_out[0][7] ),
    .S(net1025),
    .X(_2613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5175_ (.A(net1022),
    .B_N(net1142),
    .Y(_2614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5176_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\s0.shift_out[0] [0]),
    .A2(_2613_),
    .Y(_2615_),
    .B1(_2614_));
 sg13g2_nor2_1 _5177_ (.A(net1031),
    .B(_2612_),
    .Y(_2616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5178_ (.A2(_2615_),
    .A1(net1031),
    .B1(_2616_),
    .X(_2617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5179_ (.A0(\s0.data_out[0][6] ),
    .A1(\s0.data_out[1][6] ),
    .S(net1034),
    .X(_2618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5180_ (.A0(\s0.data_out[1][6] ),
    .A1(\s0.data_out[0][6] ),
    .S(net1025),
    .X(_2619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5181_ (.A(net1022),
    .B_N(net1147),
    .Y(_2620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5182_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1022),
    .A2(_2619_),
    .Y(_2621_),
    .B1(_2620_));
 sg13g2_nor2_1 _5183_ (.A(net1031),
    .B(_2618_),
    .Y(_2622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5184_ (.A2(_2621_),
    .A1(net1031),
    .B1(_2622_),
    .X(_2623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5185_ (.Y(_2624_),
    .B1(_2623_),
    .B2(net1408),
    .A2(_2617_),
    .A1(net1399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5186_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2625_),
    .B(_2623_),
    .A(net1408));
 sg13g2_or2_1 _5187_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2626_),
    .B(_2617_),
    .A(net1399));
 sg13g2_and3_1 _5188_ (.X(_2627_),
    .A(_2624_),
    .B(_2625_),
    .C(_2626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5189_ (.B(_2625_),
    .C(_2626_),
    .A(_2624_),
    .Y(_2628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5190_ (.A0(\s0.data_out[0][4] ),
    .A1(\s0.data_out[1][4] ),
    .S(net1033),
    .X(_2629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5191_ (.Y(_2630_),
    .A(net1005),
    .B(_2629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5192_ (.Y(_2631_),
    .A(net1024),
    .B(\s0.data_out[0][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5193_ (.Y(_2632_),
    .B(\s0.data_out[1][4] ),
    .A_N(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5194_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2631_),
    .A2(_2632_),
    .Y(_2633_),
    .B1(net1001));
 sg13g2_nor2b_1 _5195_ (.A(net1019),
    .B_N(net1156),
    .Y(_2634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5196_ (.B1(net1029),
    .VDD(VPWR),
    .Y(_2635_),
    .VSS(VGND),
    .A1(_2633_),
    .A2(_2634_));
 sg13g2_a21oi_1 _5197_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2630_),
    .A2(_2635_),
    .Y(_2636_),
    .B1(net1426));
 sg13g2_mux2_1 _5198_ (.A0(\s0.data_out[0][5] ),
    .A1(\s0.data_out[1][5] ),
    .S(net1034),
    .X(_2637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5199_ (.Y(_2638_),
    .A(net1006),
    .B(_2637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5200_ (.A0(\s0.data_out[1][5] ),
    .A1(\s0.data_out[0][5] ),
    .S(net1025),
    .X(_2639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5201_ (.A(net1023),
    .B_N(net1151),
    .Y(_2640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5202_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1022),
    .A2(_2639_),
    .Y(_2641_),
    .B1(_2640_));
 sg13g2_nand2b_1 _5203_ (.Y(_2642_),
    .B(net1031),
    .A_N(_2641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5204_ (.B(_2638_),
    .C(_2642_),
    .A(net1417),
    .Y(_2643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5205_ (.B(_2630_),
    .C(_2635_),
    .A(net1426),
    .Y(_2644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5206_ (.A(net1436),
    .B(_2609_),
    .Y(_2645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5207_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2638_),
    .A2(_2642_),
    .Y(_2646_),
    .B1(net1417));
 sg13g2_a21o_1 _5208_ (.A2(_2642_),
    .A1(_2638_),
    .B1(net1417),
    .X(_2647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5209_ (.B(_2644_),
    .C(_2647_),
    .A(_2643_),
    .Y(_2648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _5210_ (.A(_2628_),
    .B(_2636_),
    .C(_2645_),
    .D(_2648_),
    .Y(_2649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5211_ (.B1(_2643_),
    .VDD(VPWR),
    .Y(_2650_),
    .VSS(VGND),
    .A1(_2644_),
    .A2(_2646_));
 sg13g2_nand2b_1 _5212_ (.Y(_2651_),
    .B(_2626_),
    .A_N(_2624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5213_ (.Y(_2652_),
    .B(_2651_),
    .A_N(_2577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5214_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2627_),
    .C1(_2652_),
    .B1(_2650_),
    .A1(_2611_),
    .Y(_2653_),
    .A2(_2649_));
 sg13g2_nor3_1 _5215_ (.A(net325),
    .B(net1329),
    .C(_2653_),
    .Y(_0275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5216_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1020),
    .A2(net547),
    .Y(_2654_),
    .B1(_2598_));
 sg13g2_a21oi_1 _5217_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1004),
    .A2(_2595_),
    .Y(_2655_),
    .B1(net1346));
 sg13g2_o21ai_1 _5218_ (.B1(_2655_),
    .VDD(VPWR),
    .Y(_2656_),
    .VSS(VGND),
    .A1(net1004),
    .A2(_2654_));
 sg13g2_o21ai_1 _5219_ (.B1(_2656_),
    .VDD(VPWR),
    .Y(_2657_),
    .VSS(VGND),
    .A1(net1465),
    .A2(net652));
 sg13g2_inv_1 _5220_ (.VDD(VPWR),
    .Y(_0276_),
    .A(_2657_),
    .VSS(VGND));
 sg13g2_and2_1 _5221_ (.A(net1020),
    .B(net375),
    .X(_2658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5222_ (.B1(net1029),
    .VDD(VPWR),
    .Y(_2659_),
    .VSS(VGND),
    .A1(_2592_),
    .A2(_2658_));
 sg13g2_nor2_1 _5223_ (.A(net1346),
    .B(_2590_),
    .Y(_2660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5224_ (.Y(_0277_),
    .B1(_2659_),
    .B2(_2660_),
    .A2(_2884_),
    .A1(net1346),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5225_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1019),
    .A2(net386),
    .Y(_2661_),
    .B1(_2585_));
 sg13g2_a21oi_1 _5226_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1004),
    .A2(_2583_),
    .Y(_2662_),
    .B1(net1346));
 sg13g2_o21ai_1 _5227_ (.B1(_2662_),
    .VDD(VPWR),
    .Y(_2663_),
    .VSS(VGND),
    .A1(net1004),
    .A2(_2661_));
 sg13g2_o21ai_1 _5228_ (.B1(_2663_),
    .VDD(VPWR),
    .Y(_2664_),
    .VSS(VGND),
    .A1(net1464),
    .A2(net683));
 sg13g2_inv_1 _5229_ (.VDD(VPWR),
    .Y(_0278_),
    .A(_2664_),
    .VSS(VGND));
 sg13g2_a21oi_1 _5230_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1021),
    .A2(net402),
    .Y(_2665_),
    .B1(_2606_));
 sg13g2_a21oi_1 _5231_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1005),
    .A2(_2604_),
    .Y(_2666_),
    .B1(net1346));
 sg13g2_o21ai_1 _5232_ (.B1(_2666_),
    .VDD(VPWR),
    .Y(_2667_),
    .VSS(VGND),
    .A1(net1005),
    .A2(_2665_));
 sg13g2_o21ai_1 _5233_ (.B1(_2667_),
    .VDD(VPWR),
    .Y(_2668_),
    .VSS(VGND),
    .A1(net1465),
    .A2(net541));
 sg13g2_inv_1 _5234_ (.VDD(VPWR),
    .Y(_0279_),
    .A(net542),
    .VSS(VGND));
 sg13g2_a21oi_1 _5235_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1021),
    .A2(net385),
    .Y(_2669_),
    .B1(_2634_));
 sg13g2_a21oi_1 _5236_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1005),
    .A2(_2629_),
    .Y(_2670_),
    .B1(net1347));
 sg13g2_o21ai_1 _5237_ (.B1(_2670_),
    .VDD(VPWR),
    .Y(_2671_),
    .VSS(VGND),
    .A1(net1005),
    .A2(_2669_));
 sg13g2_o21ai_1 _5238_ (.B1(_2671_),
    .VDD(VPWR),
    .Y(_2672_),
    .VSS(VGND),
    .A1(net1467),
    .A2(net677));
 sg13g2_inv_1 _5239_ (.VDD(VPWR),
    .Y(_0280_),
    .A(_2672_),
    .VSS(VGND));
 sg13g2_a21oi_1 _5240_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1023),
    .A2(net395),
    .Y(_2673_),
    .B1(_2640_));
 sg13g2_a21oi_1 _5241_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1006),
    .A2(_2637_),
    .Y(_2674_),
    .B1(net1347));
 sg13g2_o21ai_1 _5242_ (.B1(_2674_),
    .VDD(VPWR),
    .Y(_2675_),
    .VSS(VGND),
    .A1(net1006),
    .A2(_2673_));
 sg13g2_o21ai_1 _5243_ (.B1(_2675_),
    .VDD(VPWR),
    .Y(_2676_),
    .VSS(VGND),
    .A1(net1467),
    .A2(net579));
 sg13g2_inv_1 _5244_ (.VDD(VPWR),
    .Y(_0281_),
    .A(_2676_),
    .VSS(VGND));
 sg13g2_a21oi_1 _5245_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1022),
    .A2(net394),
    .Y(_2677_),
    .B1(_2620_));
 sg13g2_a21oi_1 _5246_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2754_),
    .A2(_2618_),
    .Y(_2678_),
    .B1(net1347));
 sg13g2_o21ai_1 _5247_ (.B1(_2678_),
    .VDD(VPWR),
    .Y(_2679_),
    .VSS(VGND),
    .A1(net1006),
    .A2(_2677_));
 sg13g2_o21ai_1 _5248_ (.B1(_2679_),
    .VDD(VPWR),
    .Y(_2680_),
    .VSS(VGND),
    .A1(net1467),
    .A2(net605));
 sg13g2_inv_1 _5249_ (.VDD(VPWR),
    .Y(_0282_),
    .A(_2680_),
    .VSS(VGND));
 sg13g2_a21oi_1 _5250_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1022),
    .A2(net361),
    .Y(_2681_),
    .B1(_2614_));
 sg13g2_a21oi_1 _5251_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2754_),
    .A2(_2612_),
    .Y(_2682_),
    .B1(net1347));
 sg13g2_o21ai_1 _5252_ (.B1(_2682_),
    .VDD(VPWR),
    .Y(_2683_),
    .VSS(VGND),
    .A1(net1006),
    .A2(_2681_));
 sg13g2_o21ai_1 _5253_ (.B1(_2683_),
    .VDD(VPWR),
    .Y(_2684_),
    .VSS(VGND),
    .A1(net1467),
    .A2(net625));
 sg13g2_inv_1 _5254_ (.VDD(VPWR),
    .Y(_0283_),
    .A(_2684_),
    .VSS(VGND));
 sg13g2_a21oi_1 _5255_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net427),
    .A2(net1001),
    .Y(_2685_),
    .B1(net1392));
 sg13g2_o21ai_1 _5256_ (.B1(net1466),
    .VDD(VPWR),
    .Y(_2686_),
    .VSS(VGND),
    .A1(net1025),
    .A2(net1023));
 sg13g2_nor2_1 _5257_ (.A(_2685_),
    .B(_2686_),
    .Y(_0284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5258_ (.A(net1392),
    .B(_2686_),
    .Y(_0285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5259_ (.A(net1489),
    .B(net336),
    .X(_0286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5260_ (.A2(net395),
    .A1(net1025),
    .B1(net1023),
    .X(_2687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5261_ (.B1(_2687_),
    .VDD(VPWR),
    .Y(_2688_),
    .VSS(VGND),
    .A1(net1001),
    .A2(net1151));
 sg13g2_or2_1 _5262_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2689_),
    .B(_2688_),
    .A(net1416));
 sg13g2_a21o_1 _5263_ (.A2(net375),
    .A1(net1024),
    .B1(net1019),
    .X(_2690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5264_ (.B1(_2690_),
    .VDD(VPWR),
    .Y(_2691_),
    .VSS(VGND),
    .A1(net1001),
    .A2(net1166));
 sg13g2_nand2_1 _5265_ (.Y(_2692_),
    .A(net1019),
    .B(net1170),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5266_ (.B(net1001),
    .C(net547),
    .A(net1024),
    .Y(_2693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5267_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2693_),
    .C1(net1458),
    .B1(_2692_),
    .A1(net1449),
    .Y(_2694_),
    .A2(_2691_));
 sg13g2_a21o_1 _5268_ (.A2(net386),
    .A1(net1024),
    .B1(net1019),
    .X(_2695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5269_ (.B1(_2695_),
    .VDD(VPWR),
    .Y(_2696_),
    .VSS(VGND),
    .A1(net1001),
    .A2(net1162));
 sg13g2_nor2_1 _5270_ (.A(net1443),
    .B(_2696_),
    .Y(_2697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5271_ (.A(net1449),
    .B(_2691_),
    .Y(_2698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5272_ (.A(_2694_),
    .B(_2697_),
    .C(_2698_),
    .X(_2699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5273_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1026),
    .A2(net402),
    .Y(_2700_),
    .B1(net1019));
 sg13g2_a21oi_1 _5274_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1019),
    .A2(net993),
    .Y(_2701_),
    .B1(_2700_));
 sg13g2_inv_1 _5275_ (.VDD(VPWR),
    .Y(_2702_),
    .A(_2701_),
    .VSS(VGND));
 sg13g2_a22oi_1 _5276_ (.Y(_2703_),
    .B1(_2702_),
    .B2(net1436),
    .A2(_2696_),
    .A1(net1443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5277_ (.A2(net385),
    .A1(net1024),
    .B1(net1021),
    .X(_2704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5278_ (.B1(_2704_),
    .VDD(VPWR),
    .Y(_2705_),
    .VSS(VGND),
    .A1(net1001),
    .A2(net1156));
 sg13g2_nand2b_1 _5279_ (.Y(_2706_),
    .B(_2768_),
    .A_N(_2705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5280_ (.B1(_2706_),
    .VDD(VPWR),
    .Y(_2707_),
    .VSS(VGND),
    .A1(net1435),
    .A2(_2702_));
 sg13g2_a21oi_1 _5281_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2699_),
    .A2(_2703_),
    .Y(_2708_),
    .B1(_2707_));
 sg13g2_and2_1 _5282_ (.A(net1429),
    .B(_2705_),
    .X(_2709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5283_ (.B1(_2689_),
    .VDD(VPWR),
    .Y(_2710_),
    .VSS(VGND),
    .A1(_2708_),
    .A2(_2709_));
 sg13g2_a21o_1 _5284_ (.A2(net394),
    .A1(net1025),
    .B1(net1023),
    .X(_2711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5285_ (.B1(_2711_),
    .VDD(VPWR),
    .Y(_2712_),
    .VSS(VGND),
    .A1(net1001),
    .A2(net1147));
 sg13g2_a22oi_1 _5286_ (.Y(_2713_),
    .B1(_2712_),
    .B2(net1408),
    .A2(_2688_),
    .A1(net1416),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5287_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2714_),
    .B(_2712_),
    .A(net1408));
 sg13g2_a21o_1 _5288_ (.A2(net361),
    .A1(net1025),
    .B1(net1023),
    .X(_2715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5289_ (.B1(_2715_),
    .VDD(VPWR),
    .Y(_2716_),
    .VSS(VGND),
    .A1(_2758_),
    .A2(net1142));
 sg13g2_o21ai_1 _5290_ (.B1(_2714_),
    .VDD(VPWR),
    .Y(_2717_),
    .VSS(VGND),
    .A1(net1399),
    .A2(_2716_));
 sg13g2_a21o_1 _5291_ (.A2(_2713_),
    .A1(_2710_),
    .B1(_2717_),
    .X(_2718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5292_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1399),
    .A2(_2716_),
    .Y(_2719_),
    .B1(net1393));
 sg13g2_or2_1 _5293_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2720_),
    .B(net1329),
    .A(net333));
 sg13g2_a21oi_1 _5294_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2718_),
    .A2(_2719_),
    .Y(_0287_),
    .B1(_2720_));
 sg13g2_a21oi_1 _5295_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2692_),
    .A2(_2693_),
    .Y(_2721_),
    .B1(net1346));
 sg13g2_a21o_1 _5296_ (.A2(net547),
    .A1(net1346),
    .B1(_2721_),
    .X(_0288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5297_ (.A(net1464),
    .B(net375),
    .Y(_2722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5298_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1464),
    .A2(_2691_),
    .Y(_0289_),
    .B1(_2722_));
 sg13g2_nor2_1 _5299_ (.A(net1465),
    .B(net386),
    .Y(_2723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5300_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1464),
    .A2(_2696_),
    .Y(_0290_),
    .B1(_2723_));
 sg13g2_nor2_1 _5301_ (.A(net1464),
    .B(net402),
    .Y(_2724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5302_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1464),
    .A2(_2702_),
    .Y(_0291_),
    .B1(_2724_));
 sg13g2_nor2_1 _5303_ (.A(net1464),
    .B(net385),
    .Y(_2725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5304_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1465),
    .A2(_2705_),
    .Y(_0292_),
    .B1(_2725_));
 sg13g2_nor2_1 _5305_ (.A(net1466),
    .B(net395),
    .Y(_2726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5306_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1466),
    .A2(_2688_),
    .Y(_0293_),
    .B1(_2726_));
 sg13g2_nor2_1 _5307_ (.A(net1466),
    .B(net394),
    .Y(_2727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5308_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1466),
    .A2(_2712_),
    .Y(_0294_),
    .B1(_2727_));
 sg13g2_nor2_1 _5309_ (.A(net1466),
    .B(net361),
    .Y(_2728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5310_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1467),
    .A2(_2716_),
    .Y(_0295_),
    .B1(_2728_));
 sg13g2_inv_1 _5311_ (.VDD(VPWR),
    .Y(_2729_),
    .A(net356),
    .VSS(VGND));
 sg13g2_inv_1 _5312_ (.VDD(VPWR),
    .Y(_2730_),
    .A(net345),
    .VSS(VGND));
 sg13g2_inv_1 _5313_ (.VDD(VPWR),
    .Y(_2731_),
    .A(net364),
    .VSS(VGND));
 sg13g2_inv_1 _5314_ (.VDD(VPWR),
    .Y(_2732_),
    .A(net358),
    .VSS(VGND));
 sg13g2_inv_1 _5315_ (.VDD(VPWR),
    .Y(_2733_),
    .A(net350),
    .VSS(VGND));
 sg13g2_inv_1 _5316_ (.VDD(VPWR),
    .Y(_2734_),
    .A(net348),
    .VSS(VGND));
 sg13g2_inv_1 _5317_ (.VDD(VPWR),
    .Y(_2735_),
    .A(net362),
    .VSS(VGND));
 sg13g2_inv_1 _5318_ (.VDD(VPWR),
    .Y(_2736_),
    .A(net370),
    .VSS(VGND));
 sg13g2_inv_1 _5319_ (.VDD(VPWR),
    .Y(_2737_),
    .A(net383),
    .VSS(VGND));
 sg13g2_inv_1 _5320_ (.VDD(VPWR),
    .Y(_2738_),
    .A(net366),
    .VSS(VGND));
 sg13g2_inv_1 _5321_ (.VDD(VPWR),
    .Y(_2739_),
    .A(net392),
    .VSS(VGND));
 sg13g2_inv_2 _5322_ (.Y(_2740_),
    .A(net1212),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5323_ (.Y(_2741_),
    .A(net1217),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5324_ (.VDD(VPWR),
    .Y(_2742_),
    .A(net1471),
    .VSS(VGND));
 sg13g2_inv_1 _5325_ (.VDD(VPWR),
    .Y(_2743_),
    .A(net1394),
    .VSS(VGND));
 sg13g2_inv_2 _5326_ (.Y(_2744_),
    .A(net1195),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5327_ (.Y(_2745_),
    .A(net1187),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5328_ (.Y(_2746_),
    .A(net1138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5329_ (.Y(_2747_),
    .A(net1131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5330_ (.Y(_2748_),
    .A(net1058),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5331_ (.Y(_2749_),
    .A(net1316),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5332_ (.Y(_2750_),
    .A(net1328),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5333_ (.Y(_2751_),
    .A(net1039),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5334_ (.VDD(VPWR),
    .Y(_2752_),
    .A(net1305),
    .VSS(VGND));
 sg13g2_inv_2 _5335_ (.Y(_2753_),
    .A(net1297),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5336_ (.Y(_2754_),
    .A(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5337_ (.Y(_2755_),
    .A(net1275),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5338_ (.VDD(VPWR),
    .Y(_2756_),
    .A(net1272),
    .VSS(VGND));
 sg13g2_inv_2 _5339_ (.Y(_2757_),
    .A(net1254),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5340_ (.VDD(VPWR),
    .Y(_2758_),
    .A(net1023),
    .VSS(VGND));
 sg13g2_inv_2 _5341_ (.Y(_2759_),
    .A(net1112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5342_ (.VDD(VPWR),
    .Y(_2760_),
    .A(net1107),
    .VSS(VGND));
 sg13g2_inv_1 _5343_ (.VDD(VPWR),
    .Y(_2761_),
    .A(net1088),
    .VSS(VGND));
 sg13g2_inv_2 _5344_ (.Y(_2762_),
    .A(net1066),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5345_ (.VDD(VPWR),
    .Y(_2763_),
    .A(net377),
    .VSS(VGND));
 sg13g2_inv_1 _5346_ (.VDD(VPWR),
    .Y(_2764_),
    .A(net438),
    .VSS(VGND));
 sg13g2_inv_1 _5347_ (.VDD(VPWR),
    .Y(_2765_),
    .A(net593),
    .VSS(VGND));
 sg13g2_inv_1 _5348_ (.VDD(VPWR),
    .Y(_2766_),
    .A(net455),
    .VSS(VGND));
 sg13g2_inv_1 _5349_ (.VDD(VPWR),
    .Y(_2767_),
    .A(net459),
    .VSS(VGND));
 sg13g2_inv_8 _5350_ (.Y(_2768_),
    .A(net1426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5351_ (.VDD(VPWR),
    .Y(_2769_),
    .A(net416),
    .VSS(VGND));
 sg13g2_inv_1 _5352_ (.VDD(VPWR),
    .Y(_2770_),
    .A(net586),
    .VSS(VGND));
 sg13g2_inv_2 _5353_ (.Y(_2771_),
    .A(net354),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5354_ (.Y(_2772_),
    .A(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5355_ (.VDD(VPWR),
    .Y(_2773_),
    .A(net412),
    .VSS(VGND));
 sg13g2_inv_2 _5356_ (.Y(_2774_),
    .A(net1443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5357_ (.VDD(VPWR),
    .Y(_2775_),
    .A(net640),
    .VSS(VGND));
 sg13g2_inv_2 _5358_ (.Y(_2776_),
    .A(net381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5359_ (.VDD(VPWR),
    .Y(_2777_),
    .A(net603),
    .VSS(VGND));
 sg13g2_inv_2 _5360_ (.Y(_2778_),
    .A(net379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5361_ (.VDD(VPWR),
    .Y(_2779_),
    .A(net527),
    .VSS(VGND));
 sg13g2_inv_1 _5362_ (.VDD(VPWR),
    .Y(_2780_),
    .A(net650),
    .VSS(VGND));
 sg13g2_inv_1 _5363_ (.VDD(VPWR),
    .Y(_2781_),
    .A(net519),
    .VSS(VGND));
 sg13g2_inv_1 _5364_ (.VDD(VPWR),
    .Y(_2782_),
    .A(net557),
    .VSS(VGND));
 sg13g2_inv_1 _5365_ (.VDD(VPWR),
    .Y(_2783_),
    .A(\s0.data_out[21][0] ),
    .VSS(VGND));
 sg13g2_inv_1 _5366_ (.VDD(VPWR),
    .Y(_2784_),
    .A(net473),
    .VSS(VGND));
 sg13g2_inv_1 _5367_ (.VDD(VPWR),
    .Y(_2785_),
    .A(net432),
    .VSS(VGND));
 sg13g2_inv_2 _5368_ (.Y(_2786_),
    .A(net468),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5369_ (.Y(_2787_),
    .A(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5370_ (.VDD(VPWR),
    .Y(_2788_),
    .A(net628),
    .VSS(VGND));
 sg13g2_inv_1 _5371_ (.VDD(VPWR),
    .Y(_2789_),
    .A(net424),
    .VSS(VGND));
 sg13g2_inv_1 _5372_ (.VDD(VPWR),
    .Y(_2790_),
    .A(net633),
    .VSS(VGND));
 sg13g2_inv_1 _5373_ (.VDD(VPWR),
    .Y(_2791_),
    .A(net506),
    .VSS(VGND));
 sg13g2_inv_1 _5374_ (.VDD(VPWR),
    .Y(_2792_),
    .A(net352),
    .VSS(VGND));
 sg13g2_inv_1 _5375_ (.VDD(VPWR),
    .Y(_2793_),
    .A(net486),
    .VSS(VGND));
 sg13g2_inv_1 _5376_ (.VDD(VPWR),
    .Y(_2794_),
    .A(net690),
    .VSS(VGND));
 sg13g2_inv_1 _5377_ (.VDD(VPWR),
    .Y(_2795_),
    .A(net657),
    .VSS(VGND));
 sg13g2_inv_1 _5378_ (.VDD(VPWR),
    .Y(_2796_),
    .A(net695),
    .VSS(VGND));
 sg13g2_inv_1 _5379_ (.VDD(VPWR),
    .Y(_2797_),
    .A(net499),
    .VSS(VGND));
 sg13g2_inv_1 _5380_ (.VDD(VPWR),
    .Y(_2798_),
    .A(net436),
    .VSS(VGND));
 sg13g2_inv_1 _5381_ (.VDD(VPWR),
    .Y(_2799_),
    .A(net440),
    .VSS(VGND));
 sg13g2_inv_1 _5382_ (.VDD(VPWR),
    .Y(_2800_),
    .A(net410),
    .VSS(VGND));
 sg13g2_inv_1 _5383_ (.VDD(VPWR),
    .Y(_2801_),
    .A(net428),
    .VSS(VGND));
 sg13g2_inv_1 _5384_ (.VDD(VPWR),
    .Y(_2802_),
    .A(net418),
    .VSS(VGND));
 sg13g2_inv_1 _5385_ (.VDD(VPWR),
    .Y(_2803_),
    .A(net560),
    .VSS(VGND));
 sg13g2_inv_1 _5386_ (.VDD(VPWR),
    .Y(_2804_),
    .A(net368),
    .VSS(VGND));
 sg13g2_inv_1 _5387_ (.VDD(VPWR),
    .Y(_2805_),
    .A(net689),
    .VSS(VGND));
 sg13g2_inv_1 _5388_ (.VDD(VPWR),
    .Y(_2806_),
    .A(net511),
    .VSS(VGND));
 sg13g2_inv_2 _5389_ (.Y(_2807_),
    .A(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5390_ (.VDD(VPWR),
    .Y(_2808_),
    .A(net503),
    .VSS(VGND));
 sg13g2_inv_1 _5391_ (.VDD(VPWR),
    .Y(_2809_),
    .A(net475),
    .VSS(VGND));
 sg13g2_inv_2 _5392_ (.Y(_2810_),
    .A(net525),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5393_ (.VDD(VPWR),
    .Y(_2811_),
    .A(net482),
    .VSS(VGND));
 sg13g2_inv_1 _5394_ (.VDD(VPWR),
    .Y(_2812_),
    .A(net426),
    .VSS(VGND));
 sg13g2_inv_1 _5395_ (.VDD(VPWR),
    .Y(_2813_),
    .A(net479),
    .VSS(VGND));
 sg13g2_inv_1 _5396_ (.VDD(VPWR),
    .Y(_2814_),
    .A(net561),
    .VSS(VGND));
 sg13g2_inv_1 _5397_ (.VDD(VPWR),
    .Y(_2815_),
    .A(net430),
    .VSS(VGND));
 sg13g2_inv_1 _5398_ (.VDD(VPWR),
    .Y(_2816_),
    .A(net553),
    .VSS(VGND));
 sg13g2_inv_1 _5399_ (.VDD(VPWR),
    .Y(_2817_),
    .A(net420),
    .VSS(VGND));
 sg13g2_inv_1 _5400_ (.VDD(VPWR),
    .Y(_2818_),
    .A(net530),
    .VSS(VGND));
 sg13g2_inv_2 _5401_ (.Y(_2819_),
    .A(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5402_ (.Y(_2820_),
    .A(net545),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _5403_ (.Y(_2821_),
    .A(\s0.data_out[14][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5404_ (.VDD(VPWR),
    .Y(_2822_),
    .A(net602),
    .VSS(VGND));
 sg13g2_inv_1 _5405_ (.VDD(VPWR),
    .Y(_2823_),
    .A(net548),
    .VSS(VGND));
 sg13g2_inv_1 _5406_ (.VDD(VPWR),
    .Y(_2824_),
    .A(net647),
    .VSS(VGND));
 sg13g2_inv_1 _5407_ (.VDD(VPWR),
    .Y(_2825_),
    .A(net406),
    .VSS(VGND));
 sg13g2_inv_1 _5408_ (.VDD(VPWR),
    .Y(_2826_),
    .A(net491),
    .VSS(VGND));
 sg13g2_inv_1 _5409_ (.VDD(VPWR),
    .Y(_2827_),
    .A(net532),
    .VSS(VGND));
 sg13g2_inv_1 _5410_ (.VDD(VPWR),
    .Y(_2828_),
    .A(net457),
    .VSS(VGND));
 sg13g2_inv_1 _5411_ (.VDD(VPWR),
    .Y(_2829_),
    .A(net481),
    .VSS(VGND));
 sg13g2_inv_1 _5412_ (.VDD(VPWR),
    .Y(_2830_),
    .A(net595),
    .VSS(VGND));
 sg13g2_inv_1 _5413_ (.VDD(VPWR),
    .Y(_2831_),
    .A(net619),
    .VSS(VGND));
 sg13g2_inv_1 _5414_ (.VDD(VPWR),
    .Y(_2832_),
    .A(net467),
    .VSS(VGND));
 sg13g2_inv_1 _5415_ (.VDD(VPWR),
    .Y(_2833_),
    .A(net442),
    .VSS(VGND));
 sg13g2_inv_1 _5416_ (.VDD(VPWR),
    .Y(_2834_),
    .A(net451),
    .VSS(VGND));
 sg13g2_inv_1 _5417_ (.VDD(VPWR),
    .Y(_2835_),
    .A(net373),
    .VSS(VGND));
 sg13g2_inv_1 _5418_ (.VDD(VPWR),
    .Y(_2836_),
    .A(net461),
    .VSS(VGND));
 sg13g2_inv_1 _5419_ (.VDD(VPWR),
    .Y(_2837_),
    .A(net422),
    .VSS(VGND));
 sg13g2_inv_1 _5420_ (.VDD(VPWR),
    .Y(_2838_),
    .A(net588),
    .VSS(VGND));
 sg13g2_inv_1 _5421_ (.VDD(VPWR),
    .Y(_2839_),
    .A(net489),
    .VSS(VGND));
 sg13g2_inv_1 _5422_ (.VDD(VPWR),
    .Y(_2840_),
    .A(net477),
    .VSS(VGND));
 sg13g2_inv_1 _5423_ (.VDD(VPWR),
    .Y(_2841_),
    .A(net536),
    .VSS(VGND));
 sg13g2_inv_1 _5424_ (.VDD(VPWR),
    .Y(_2842_),
    .A(net636),
    .VSS(VGND));
 sg13g2_inv_1 _5425_ (.VDD(VPWR),
    .Y(_2843_),
    .A(net572),
    .VSS(VGND));
 sg13g2_inv_1 _5426_ (.VDD(VPWR),
    .Y(_2844_),
    .A(net589),
    .VSS(VGND));
 sg13g2_inv_1 _5427_ (.VDD(VPWR),
    .Y(_2845_),
    .A(net465),
    .VSS(VGND));
 sg13g2_inv_1 _5428_ (.VDD(VPWR),
    .Y(_2846_),
    .A(net505),
    .VSS(VGND));
 sg13g2_inv_1 _5429_ (.VDD(VPWR),
    .Y(_2847_),
    .A(net509),
    .VSS(VGND));
 sg13g2_inv_1 _5430_ (.VDD(VPWR),
    .Y(_2848_),
    .A(net371),
    .VSS(VGND));
 sg13g2_inv_1 _5431_ (.VDD(VPWR),
    .Y(_2849_),
    .A(net687),
    .VSS(VGND));
 sg13g2_inv_1 _5432_ (.VDD(VPWR),
    .Y(_2850_),
    .A(net670),
    .VSS(VGND));
 sg13g2_inv_1 _5433_ (.VDD(VPWR),
    .Y(_2851_),
    .A(net637),
    .VSS(VGND));
 sg13g2_inv_1 _5434_ (.VDD(VPWR),
    .Y(_2852_),
    .A(net518),
    .VSS(VGND));
 sg13g2_inv_1 _5435_ (.VDD(VPWR),
    .Y(_2853_),
    .A(net673),
    .VSS(VGND));
 sg13g2_inv_2 _5436_ (.Y(_2854_),
    .A(net537),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5437_ (.VDD(VPWR),
    .Y(_2855_),
    .A(net555),
    .VSS(VGND));
 sg13g2_inv_1 _5438_ (.VDD(VPWR),
    .Y(_2856_),
    .A(net470),
    .VSS(VGND));
 sg13g2_inv_1 _5439_ (.VDD(VPWR),
    .Y(_2857_),
    .A(net632),
    .VSS(VGND));
 sg13g2_inv_1 _5440_ (.VDD(VPWR),
    .Y(_2858_),
    .A(net453),
    .VSS(VGND));
 sg13g2_inv_1 _5441_ (.VDD(VPWR),
    .Y(_2859_),
    .A(net408),
    .VSS(VGND));
 sg13g2_inv_1 _5442_ (.VDD(VPWR),
    .Y(_2860_),
    .A(net404),
    .VSS(VGND));
 sg13g2_inv_1 _5443_ (.VDD(VPWR),
    .Y(_2861_),
    .A(net578),
    .VSS(VGND));
 sg13g2_inv_1 _5444_ (.VDD(VPWR),
    .Y(_2862_),
    .A(net389),
    .VSS(VGND));
 sg13g2_inv_1 _5445_ (.VDD(VPWR),
    .Y(_2863_),
    .A(net501),
    .VSS(VGND));
 sg13g2_inv_1 _5446_ (.VDD(VPWR),
    .Y(_2864_),
    .A(net692),
    .VSS(VGND));
 sg13g2_inv_1 _5447_ (.VDD(VPWR),
    .Y(_2865_),
    .A(net656),
    .VSS(VGND));
 sg13g2_inv_1 _5448_ (.VDD(VPWR),
    .Y(_2866_),
    .A(net549),
    .VSS(VGND));
 sg13g2_inv_1 _5449_ (.VDD(VPWR),
    .Y(_2867_),
    .A(net488),
    .VSS(VGND));
 sg13g2_inv_1 _5450_ (.VDD(VPWR),
    .Y(_2868_),
    .A(net449),
    .VSS(VGND));
 sg13g2_inv_1 _5451_ (.VDD(VPWR),
    .Y(_2869_),
    .A(net492),
    .VSS(VGND));
 sg13g2_inv_1 _5452_ (.VDD(VPWR),
    .Y(_2870_),
    .A(net507),
    .VSS(VGND));
 sg13g2_inv_1 _5453_ (.VDD(VPWR),
    .Y(_2871_),
    .A(net444),
    .VSS(VGND));
 sg13g2_inv_1 _5454_ (.VDD(VPWR),
    .Y(_2872_),
    .A(net676),
    .VSS(VGND));
 sg13g2_inv_1 _5455_ (.VDD(VPWR),
    .Y(_2873_),
    .A(net642),
    .VSS(VGND));
 sg13g2_inv_1 _5456_ (.VDD(VPWR),
    .Y(_2874_),
    .A(net484),
    .VSS(VGND));
 sg13g2_inv_1 _5457_ (.VDD(VPWR),
    .Y(_2875_),
    .A(net601),
    .VSS(VGND));
 sg13g2_inv_1 _5458_ (.VDD(VPWR),
    .Y(_2876_),
    .A(net387),
    .VSS(VGND));
 sg13g2_inv_1 _5459_ (.VDD(VPWR),
    .Y(_2877_),
    .A(net574),
    .VSS(VGND));
 sg13g2_inv_1 _5460_ (.VDD(VPWR),
    .Y(_2878_),
    .A(net434),
    .VSS(VGND));
 sg13g2_inv_1 _5461_ (.VDD(VPWR),
    .Y(_2879_),
    .A(net400),
    .VSS(VGND));
 sg13g2_inv_1 _5462_ (.VDD(VPWR),
    .Y(_2880_),
    .A(net512),
    .VSS(VGND));
 sg13g2_inv_1 _5463_ (.VDD(VPWR),
    .Y(_2881_),
    .A(net580),
    .VSS(VGND));
 sg13g2_inv_1 _5464_ (.VDD(VPWR),
    .Y(_2882_),
    .A(net463),
    .VSS(VGND));
 sg13g2_inv_1 _5465_ (.VDD(VPWR),
    .Y(_2883_),
    .A(net514),
    .VSS(VGND));
 sg13g2_inv_1 _5466_ (.VDD(VPWR),
    .Y(_2884_),
    .A(net494),
    .VSS(VGND));
 sg13g2_nor2_1 _5467_ (.A(\s0.was_valid_out[23] [0]),
    .B(net1326),
    .Y(_2885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5468_ (.Y(_2886_),
    .A(net1458),
    .B(net992),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5469_ (.B1(_2886_),
    .VDD(VPWR),
    .Y(net2),
    .VSS(VGND),
    .A1(_2778_),
    .A2(net992));
 sg13g2_nand2_1 _5470_ (.Y(_2887_),
    .A(net1449),
    .B(_2885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5471_ (.B1(_2887_),
    .VDD(VPWR),
    .Y(net3),
    .VSS(VGND),
    .A1(_2776_),
    .A2(net992));
 sg13g2_nor2_1 _5472_ (.A(\s0.data_out[23][2] ),
    .B(net992),
    .Y(_2888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5473_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1334),
    .A2(net992),
    .Y(net4),
    .B1(_2888_));
 sg13g2_nand2_1 _5474_ (.Y(_2889_),
    .A(net1435),
    .B(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5475_ (.B1(_2889_),
    .VDD(VPWR),
    .Y(net5),
    .VSS(VGND),
    .A1(_2771_),
    .A2(net992));
 sg13g2_nor2_1 _5476_ (.A(\s0.data_out[23][4] ),
    .B(net991),
    .Y(_2890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5477_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2768_),
    .A2(net991),
    .Y(net6),
    .B1(_2890_));
 sg13g2_nand2_1 _5478_ (.Y(_2891_),
    .A(net1416),
    .B(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5479_ (.B1(_2891_),
    .VDD(VPWR),
    .Y(net7),
    .VSS(VGND),
    .A1(_2767_),
    .A2(net991));
 sg13g2_nand2_1 _5480_ (.Y(_2892_),
    .A(net1407),
    .B(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5481_ (.B1(_2892_),
    .VDD(VPWR),
    .Y(net8),
    .VSS(VGND),
    .A1(_2766_),
    .A2(net991));
 sg13g2_nand2_1 _5482_ (.Y(_2893_),
    .A(net1398),
    .B(net992),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5483_ (.B1(_2893_),
    .VDD(VPWR),
    .Y(net9),
    .VSS(VGND),
    .A1(_2764_),
    .A2(net991));
 sg13g2_and2_1 _5484_ (.A(net1466),
    .B(net333),
    .X(_0000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5485_ (.B1(net1324),
    .VDD(VPWR),
    .Y(_2894_),
    .VSS(VGND),
    .A1(net1392),
    .A2(net1312));
 sg13g2_nand2_1 _5486_ (.Y(_2895_),
    .A(net1336),
    .B(net1318),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5487_ (.Y(_2896_),
    .B(_2895_),
    .A_N(_2894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5488_ (.A(net1392),
    .B(_2750_),
    .Y(_2897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5489_ (.B1(_2896_),
    .VDD(VPWR),
    .Y(_2898_),
    .VSS(VGND),
    .A1(net1324),
    .A2(_2897_));
 sg13g2_nor2_1 _5490_ (.A(net392),
    .B(net1318),
    .Y(_2899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5491_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2900_),
    .B(_2899_),
    .A(_2896_));
 sg13g2_nor2_1 _5492_ (.A(net1312),
    .B(_2894_),
    .Y(_2901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5493_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2739_),
    .A2(_2750_),
    .Y(_2902_),
    .B1(net1324));
 sg13g2_nor2_1 _5494_ (.A(_2901_),
    .B(_2902_),
    .Y(_2903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5495_ (.B1(net1463),
    .VDD(VPWR),
    .Y(_2904_),
    .VSS(VGND),
    .A1(net559),
    .A2(_2898_));
 sg13g2_a21oi_1 _5496_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2900_),
    .A2(_2903_),
    .Y(_0001_),
    .B1(_2904_));
 sg13g2_nor2_1 _5497_ (.A(net1340),
    .B(_2898_),
    .Y(_0002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5498_ (.A(net1462),
    .B(net330),
    .X(_0003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5499_ (.A(net412),
    .B_N(net1328),
    .Y(_2905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5500_ (.A(net1328),
    .B(\s0.data_out[22][2] ),
    .Y(_2906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5501_ (.A(net1325),
    .B(_2905_),
    .C(_2906_),
    .Y(_2907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5502_ (.A0(\s0.data_out[23][2] ),
    .A1(\s0.data_out[22][2] ),
    .S(net1320),
    .X(_2908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5503_ (.A(net1315),
    .B_N(net1162),
    .Y(_2909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5504_ (.A2(_2908_),
    .A1(net1315),
    .B1(_2909_),
    .X(_2910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5505_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1325),
    .A2(_2910_),
    .Y(_2911_),
    .B1(_2907_));
 sg13g2_or2_1 _5506_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2912_),
    .B(_2911_),
    .A(net1443));
 sg13g2_a21o_1 _5507_ (.A2(_2775_),
    .A1(_2750_),
    .B1(net1325),
    .X(_2913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5508_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1328),
    .A2(_2776_),
    .Y(_2914_),
    .B1(_2913_));
 sg13g2_nand2_1 _5509_ (.Y(_2915_),
    .A(net1321),
    .B(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5510_ (.B1(_2915_),
    .VDD(VPWR),
    .Y(_2916_),
    .VSS(VGND),
    .A1(net1320),
    .A2(_2776_));
 sg13g2_nor2b_1 _5511_ (.A(net1315),
    .B_N(net1166),
    .Y(_2917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5512_ (.A2(_2916_),
    .A1(net1315),
    .B1(_2917_),
    .X(_2918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5513_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1325),
    .A2(_2918_),
    .Y(_2919_),
    .B1(_2914_));
 sg13g2_nand2_1 _5514_ (.Y(_2920_),
    .A(net1449),
    .B(_2919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5515_ (.A2(_2777_),
    .A1(_2750_),
    .B1(net1325),
    .X(_2921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5516_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1328),
    .A2(_2778_),
    .Y(_2922_),
    .B1(_2921_));
 sg13g2_nand2_1 _5517_ (.Y(_2923_),
    .A(net1321),
    .B(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5518_ (.B1(_2923_),
    .VDD(VPWR),
    .Y(_2924_),
    .VSS(VGND),
    .A1(net1320),
    .A2(_2778_));
 sg13g2_nor2b_1 _5519_ (.A(net1315),
    .B_N(net1170),
    .Y(_2925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5520_ (.A2(_2924_),
    .A1(net1315),
    .B1(_2925_),
    .X(_2926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5521_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1325),
    .A2(_2926_),
    .Y(_2927_),
    .B1(_2922_));
 sg13g2_nor2_1 _5522_ (.A(net1458),
    .B(_2927_),
    .Y(_2928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5523_ (.B1(_2912_),
    .VDD(VPWR),
    .Y(_2929_),
    .VSS(VGND),
    .A1(net1449),
    .A2(_2919_));
 sg13g2_a21oi_1 _5524_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2920_),
    .A2(_2928_),
    .Y(_2930_),
    .B1(_2929_));
 sg13g2_a21o_1 _5525_ (.A2(_2770_),
    .A1(_2750_),
    .B1(net1326),
    .X(_2931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5526_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1328),
    .A2(_2771_),
    .Y(_2932_),
    .B1(_2931_));
 sg13g2_nand2_1 _5527_ (.Y(_2933_),
    .A(net1320),
    .B(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5528_ (.B1(_2933_),
    .VDD(VPWR),
    .Y(_2934_),
    .VSS(VGND),
    .A1(net1320),
    .A2(_2771_));
 sg13g2_nor2_1 _5529_ (.A(net1315),
    .B(net993),
    .Y(_2935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5530_ (.A2(_2934_),
    .A1(net1315),
    .B1(_2935_),
    .X(_2936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5531_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1326),
    .A2(_2936_),
    .Y(_2937_),
    .B1(_2932_));
 sg13g2_a22oi_1 _5532_ (.Y(_2938_),
    .B1(_2937_),
    .B2(net1435),
    .A2(_2911_),
    .A1(net1443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5533_ (.VDD(VPWR),
    .Y(_2939_),
    .A(_2938_),
    .VSS(VGND));
 sg13g2_nor2b_1 _5534_ (.A(net438),
    .B_N(net1327),
    .Y(_2940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5535_ (.A(net1327),
    .B(net377),
    .Y(_2941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5536_ (.A(net1323),
    .B(_2940_),
    .C(_2941_),
    .Y(_2942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5537_ (.Y(_2943_),
    .A(net1319),
    .B(net377),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5538_ (.A0(\s0.data_out[23][7] ),
    .A1(\s0.data_out[22][7] ),
    .S(net1318),
    .X(_2944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5539_ (.A(net1311),
    .B_N(net1142),
    .Y(_2945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5540_ (.A2(_2944_),
    .A1(net1311),
    .B1(_2945_),
    .X(_2946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5541_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1323),
    .A2(_2946_),
    .Y(_2947_),
    .B1(_2942_));
 sg13g2_nor2b_1 _5542_ (.A(net455),
    .B_N(net1327),
    .Y(_2948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5543_ (.A(net1327),
    .B(\s0.data_out[22][6] ),
    .Y(_2949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5544_ (.A(net1323),
    .B(_2948_),
    .C(_2949_),
    .Y(_2950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5545_ (.Y(_2951_),
    .A(net1319),
    .B(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5546_ (.A0(\s0.data_out[23][6] ),
    .A1(\s0.data_out[22][6] ),
    .S(net1318),
    .X(_2952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5547_ (.A(net1311),
    .B_N(net1147),
    .Y(_2953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5548_ (.A2(_2952_),
    .A1(net1311),
    .B1(_2953_),
    .X(_2954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5549_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1323),
    .A2(_2954_),
    .Y(_2955_),
    .B1(_2950_));
 sg13g2_a22oi_1 _5550_ (.Y(_2956_),
    .B1(_2955_),
    .B2(net1407),
    .A2(_2947_),
    .A1(net1398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5551_ (.A(net1398),
    .B(_2947_),
    .Y(_2957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5552_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2958_),
    .B(_2955_),
    .A(net1407));
 sg13g2_nand3b_1 _5553_ (.B(_2958_),
    .C(_2956_),
    .Y(_2959_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2957_));
 sg13g2_nor2b_1 _5554_ (.A(net416),
    .B_N(net1327),
    .Y(_2960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5555_ (.A(net1327),
    .B(\s0.data_out[22][4] ),
    .Y(_2961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5556_ (.A(net1324),
    .B(_2960_),
    .C(_2961_),
    .Y(_2962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5557_ (.A0(\s0.data_out[23][4] ),
    .A1(\s0.data_out[22][4] ),
    .S(net1318),
    .X(_2963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5558_ (.A(net1312),
    .B_N(net1156),
    .Y(_2964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5559_ (.A2(_2963_),
    .A1(net1311),
    .B1(_2964_),
    .X(_2965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5560_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1324),
    .A2(_2965_),
    .Y(_2966_),
    .B1(_2962_));
 sg13g2_nor2b_1 _5561_ (.A(net459),
    .B_N(net1327),
    .Y(_2967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5562_ (.A(net1327),
    .B(\s0.data_out[22][5] ),
    .Y(_2968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5563_ (.A(net1323),
    .B(_2967_),
    .C(_2968_),
    .Y(_2969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5564_ (.A0(\s0.data_out[23][5] ),
    .A1(\s0.data_out[22][5] ),
    .S(net1318),
    .X(_2970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5565_ (.A(net1311),
    .B_N(net1151),
    .Y(_2971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5566_ (.A2(_2970_),
    .A1(net1311),
    .B1(_2971_),
    .X(_2972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5567_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1323),
    .A2(_2972_),
    .Y(_2973_),
    .B1(_2969_));
 sg13g2_a22oi_1 _5568_ (.Y(_2974_),
    .B1(_2973_),
    .B2(net1416),
    .A2(_2966_),
    .A1(net1426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5569_ (.A(net1435),
    .B(_2937_),
    .Y(_2975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5570_ (.A(net1416),
    .B(_2973_),
    .Y(_2976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5571_ (.B1(_2974_),
    .VDD(VPWR),
    .Y(_2977_),
    .VSS(VGND),
    .A1(net1426),
    .A2(_2966_));
 sg13g2_nor4_1 _5572_ (.A(_2959_),
    .B(_2975_),
    .C(_2976_),
    .D(_2977_),
    .Y(_2978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5573_ (.B1(_2978_),
    .VDD(VPWR),
    .Y(_2979_),
    .VSS(VGND),
    .A1(_2930_),
    .A2(_2939_));
 sg13g2_nor3_1 _5574_ (.A(_2959_),
    .B(_2974_),
    .C(_2976_),
    .Y(_2980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5575_ (.A(_2956_),
    .B(_2957_),
    .Y(_2981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5576_ (.A(_2898_),
    .B(_2980_),
    .C(_2981_),
    .Y(_2982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5577_ (.Y(_2983_),
    .A(net1390),
    .B(net1464),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5578_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2984_),
    .B(net1329),
    .A(net335));
 sg13g2_a21oi_1 _5579_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2979_),
    .A2(_2982_),
    .Y(_0004_),
    .B1(_2984_));
 sg13g2_nor2_1 _5580_ (.A(net1011),
    .B(_2777_),
    .Y(_2985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5581_ (.B1(net1326),
    .VDD(VPWR),
    .Y(_2986_),
    .VSS(VGND),
    .A1(_2925_),
    .A2(_2985_));
 sg13g2_nor2_1 _5582_ (.A(net1341),
    .B(_2922_),
    .Y(_2987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5583_ (.Y(_0005_),
    .B1(_2986_),
    .B2(_2987_),
    .A2(_2778_),
    .A1(net1341),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5584_ (.A(net1011),
    .B(_2775_),
    .Y(_2988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5585_ (.B1(net1325),
    .VDD(VPWR),
    .Y(_2989_),
    .VSS(VGND),
    .A1(_2917_),
    .A2(_2988_));
 sg13g2_nor2_1 _5586_ (.A(net1341),
    .B(_2914_),
    .Y(_2990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5587_ (.Y(_0006_),
    .B1(_2989_),
    .B2(_2990_),
    .A2(_2776_),
    .A1(net1341),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5588_ (.A(net1317),
    .B(\s0.data_out[22][2] ),
    .X(_2991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5589_ (.B1(net1325),
    .VDD(VPWR),
    .Y(_2992_),
    .VSS(VGND),
    .A1(_2909_),
    .A2(_2991_));
 sg13g2_nor2_1 _5590_ (.A(net1341),
    .B(_2907_),
    .Y(_2993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5591_ (.Y(_0007_),
    .B1(_2992_),
    .B2(_2993_),
    .A2(_2773_),
    .A1(net1341),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5592_ (.A(net1011),
    .B(_2770_),
    .Y(_2994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5593_ (.B1(net1326),
    .VDD(VPWR),
    .Y(_2995_),
    .VSS(VGND),
    .A1(_2935_),
    .A2(_2994_));
 sg13g2_nor2_1 _5594_ (.A(net1340),
    .B(net355),
    .Y(_2996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5595_ (.Y(_0008_),
    .B1(net399),
    .B2(_2996_),
    .A2(_2771_),
    .A1(net1340),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5596_ (.A(net1312),
    .B(\s0.data_out[22][4] ),
    .X(_2997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5597_ (.B1(net1324),
    .VDD(VPWR),
    .Y(_2998_),
    .VSS(VGND),
    .A1(_2964_),
    .A2(_2997_));
 sg13g2_nor2_1 _5598_ (.A(net1339),
    .B(_2962_),
    .Y(_2999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5599_ (.Y(_0009_),
    .B1(_2998_),
    .B2(_2999_),
    .A2(_2769_),
    .A1(net1339),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5600_ (.A(net1311),
    .B(\s0.data_out[22][5] ),
    .X(_3000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5601_ (.B1(net1323),
    .VDD(VPWR),
    .Y(_3001_),
    .VSS(VGND),
    .A1(_2971_),
    .A2(_3000_));
 sg13g2_nor2_1 _5602_ (.A(net1339),
    .B(_2969_),
    .Y(_3002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5603_ (.Y(_0010_),
    .B1(_3001_),
    .B2(_3002_),
    .A2(_2767_),
    .A1(net1339),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5604_ (.A(net1012),
    .B(_2765_),
    .Y(_3003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5605_ (.B1(net1324),
    .VDD(VPWR),
    .Y(_3004_),
    .VSS(VGND),
    .A1(_2953_),
    .A2(_3003_));
 sg13g2_nor2_1 _5606_ (.A(net1339),
    .B(_2950_),
    .Y(_3005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5607_ (.Y(_0011_),
    .B1(_3004_),
    .B2(_3005_),
    .A2(_2766_),
    .A1(net1339),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5608_ (.A(net1012),
    .B(_2763_),
    .Y(_3006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5609_ (.B1(net1323),
    .VDD(VPWR),
    .Y(_3007_),
    .VSS(VGND),
    .A1(_2945_),
    .A2(_3006_));
 sg13g2_nor2_1 _5610_ (.A(net1339),
    .B(_2942_),
    .Y(_3008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5611_ (.Y(_0012_),
    .B1(_3007_),
    .B2(_3008_),
    .A2(_2764_),
    .A1(net1339),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5612_ (.B1(net1313),
    .VDD(VPWR),
    .Y(_3009_),
    .VSS(VGND),
    .A1(net1392),
    .A2(net1300));
 sg13g2_a21oi_1 _5613_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1336),
    .A2(net1307),
    .Y(_3010_),
    .B1(_3009_));
 sg13g2_a21oi_1 _5614_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1012),
    .A2(_2895_),
    .Y(_3011_),
    .B1(_3010_));
 sg13g2_o21ai_1 _5615_ (.B1(_3010_),
    .VDD(VPWR),
    .Y(_3012_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[21] [0]),
    .A2(net1307));
 sg13g2_nor2_1 _5616_ (.A(net1302),
    .B(_3009_),
    .Y(_3013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5617_ (.B1(net1012),
    .VDD(VPWR),
    .Y(_3014_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[21] [0]),
    .A2(net1318));
 sg13g2_nand2_1 _5618_ (.Y(_3015_),
    .A(_3012_),
    .B(_3014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5619_ (.B1(net1463),
    .VDD(VPWR),
    .Y(_3016_),
    .VSS(VGND),
    .A1(_3013_),
    .A2(_3015_));
 sg13g2_a21oi_1 _5620_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2739_),
    .A2(_3011_),
    .Y(_0013_),
    .B1(_3016_));
 sg13g2_and2_1 _5621_ (.A(net1463),
    .B(_3011_),
    .X(_0014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5622_ (.A(net1462),
    .B(net332),
    .X(_0015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5623_ (.Y(_3017_),
    .A(net1309),
    .B(net557),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5624_ (.A0(\s0.data_out[22][1] ),
    .A1(\s0.data_out[21][1] ),
    .S(net1307),
    .X(_3018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5625_ (.A(net1303),
    .B_N(net1166),
    .Y(_3019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5626_ (.A2(_3018_),
    .A1(net1303),
    .B1(_3019_),
    .X(_3020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5627_ (.Y(_3021_),
    .B(net557),
    .A_N(net1320),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5628_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2915_),
    .A2(_3021_),
    .Y(_3022_),
    .B1(net1316));
 sg13g2_a21oi_1 _5629_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1317),
    .A2(_3020_),
    .Y(_3023_),
    .B1(_3022_));
 sg13g2_o21ai_1 _5630_ (.B1(_2923_),
    .VDD(VPWR),
    .Y(_3024_),
    .VSS(VGND),
    .A1(net1321),
    .A2(_2783_));
 sg13g2_nand2_1 _5631_ (.Y(_3025_),
    .A(net1011),
    .B(_3024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5632_ (.A(net1303),
    .B_N(net1170),
    .Y(_3026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5633_ (.A0(\s0.data_out[22][0] ),
    .A1(\s0.data_out[21][0] ),
    .S(net1310),
    .X(_3027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5634_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1303),
    .A2(_3027_),
    .Y(_3028_),
    .B1(_3026_));
 sg13g2_nand2b_1 _5635_ (.Y(_3029_),
    .B(net1316),
    .A_N(_3028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5636_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_3029_),
    .C1(net1458),
    .B1(_3025_),
    .A1(net1449),
    .Y(_3030_),
    .A2(_3023_));
 sg13g2_nor2_1 _5637_ (.A(net1449),
    .B(_3023_),
    .Y(_3031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5638_ (.Y(_3032_),
    .A(net1309),
    .B(net519),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5639_ (.A0(\s0.data_out[22][3] ),
    .A1(\s0.data_out[21][3] ),
    .S(net1307),
    .X(_3033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5640_ (.A(net1303),
    .B_N(net1161),
    .Y(_3034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5641_ (.A2(_3033_),
    .A1(net1303),
    .B1(_3034_),
    .X(_3035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5642_ (.Y(_3036_),
    .B(net519),
    .A_N(net1320),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5643_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2933_),
    .A2(_3036_),
    .Y(_3037_),
    .B1(net1316));
 sg13g2_a21oi_1 _5644_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1316),
    .A2(_3035_),
    .Y(_3038_),
    .B1(_3037_));
 sg13g2_nor2_1 _5645_ (.A(net1435),
    .B(_3038_),
    .Y(_3039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5646_ (.A0(\s0.data_out[22][2] ),
    .A1(\s0.data_out[21][2] ),
    .S(net1310),
    .X(_3040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5647_ (.A(net1303),
    .B_N(net1162),
    .Y(_3041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5648_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1304),
    .A2(_3040_),
    .Y(_3042_),
    .B1(_3041_));
 sg13g2_mux2_1 _5649_ (.A0(\s0.data_out[21][2] ),
    .A1(\s0.data_out[22][2] ),
    .S(net1320),
    .X(_3043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5650_ (.Y(_3044_),
    .A(_2749_),
    .B(_3043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5651_ (.B1(_3044_),
    .VDD(VPWR),
    .Y(_3045_),
    .VSS(VGND),
    .A1(net1011),
    .A2(_3042_));
 sg13g2_or2_1 _5652_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_3046_),
    .B(_3045_),
    .A(net1334));
 sg13g2_xnor2_1 _5653_ (.Y(_3047_),
    .A(net1334),
    .B(_3045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _5654_ (.A(_3030_),
    .B(_3031_),
    .C(_3039_),
    .D(_3047_),
    .Y(_3048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5655_ (.Y(_3049_),
    .A(net1435),
    .B(_3038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5656_ (.B1(_3049_),
    .VDD(VPWR),
    .Y(_3050_),
    .VSS(VGND),
    .A1(_3039_),
    .A2(_3046_));
 sg13g2_nor2_1 _5657_ (.A(_3048_),
    .B(_3050_),
    .Y(_3051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5658_ (.Y(_3052_),
    .A(net1308),
    .B(net527),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5659_ (.A0(\s0.data_out[22][7] ),
    .A1(\s0.data_out[21][7] ),
    .S(net1307),
    .X(_3053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5660_ (.A(net1300),
    .B_N(net1142),
    .Y(_3054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5661_ (.A2(_3053_),
    .A1(net1300),
    .B1(_3054_),
    .X(_3055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5662_ (.Y(_3056_),
    .B(\s0.data_out[21][7] ),
    .A_N(net1318),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5663_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2943_),
    .A2(_3056_),
    .Y(_3057_),
    .B1(net1313));
 sg13g2_a21oi_1 _5664_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1313),
    .A2(_3055_),
    .Y(_3058_),
    .B1(_3057_));
 sg13g2_nand2_1 _5665_ (.Y(_3059_),
    .A(net1308),
    .B(net650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5666_ (.A0(\s0.data_out[22][6] ),
    .A1(\s0.data_out[21][6] ),
    .S(net1307),
    .X(_3060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5667_ (.A(net1300),
    .B_N(net1147),
    .Y(_3061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5668_ (.A2(_3060_),
    .A1(net1300),
    .B1(_3061_),
    .X(_3062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5669_ (.Y(_3063_),
    .B(\s0.data_out[21][6] ),
    .A_N(net1319),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5670_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2951_),
    .A2(_3063_),
    .Y(_3064_),
    .B1(net1313));
 sg13g2_a21oi_1 _5671_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1313),
    .A2(_3062_),
    .Y(_3065_),
    .B1(_3064_));
 sg13g2_a22oi_1 _5672_ (.Y(_3066_),
    .B1(_3065_),
    .B2(net1407),
    .A2(_3058_),
    .A1(net1398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5673_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_3067_),
    .B(_3065_),
    .A(net1407));
 sg13g2_nor2_1 _5674_ (.A(net1398),
    .B(_3058_),
    .Y(_3068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _5675_ (.B(_3066_),
    .C(_3067_),
    .Y(_3069_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_3068_));
 sg13g2_nor2b_1 _5676_ (.A(net1304),
    .B_N(net1156),
    .Y(_3070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5677_ (.Y(_3071_),
    .A(net1309),
    .B(\s0.data_out[21][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5678_ (.A0(\s0.data_out[22][4] ),
    .A1(\s0.data_out[21][4] ),
    .S(net1307),
    .X(_3072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5679_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1304),
    .A2(_3072_),
    .Y(_3073_),
    .B1(_3070_));
 sg13g2_nand2b_1 _5680_ (.Y(_3074_),
    .B(net1314),
    .A_N(_3073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5681_ (.A0(\s0.data_out[21][4] ),
    .A1(\s0.data_out[22][4] ),
    .S(net1321),
    .X(_3075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5682_ (.Y(_3076_),
    .A(net1012),
    .B(_3075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5683_ (.B(_3074_),
    .C(_3076_),
    .A(net1426),
    .Y(_3077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5684_ (.Y(_3078_),
    .A(net1308),
    .B(\s0.data_out[21][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5685_ (.A0(\s0.data_out[22][5] ),
    .A1(\s0.data_out[21][5] ),
    .S(net1307),
    .X(_3079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5686_ (.A(net1300),
    .B_N(net1151),
    .Y(_3080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5687_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1300),
    .A2(_3079_),
    .Y(_3081_),
    .B1(_3080_));
 sg13g2_nand2b_1 _5688_ (.Y(_3082_),
    .B(net1313),
    .A_N(_3081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5689_ (.A0(\s0.data_out[21][5] ),
    .A1(\s0.data_out[22][5] ),
    .S(net1319),
    .X(_3083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5690_ (.Y(_3084_),
    .A(net1012),
    .B(_3083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5691_ (.B(_3082_),
    .C(_3084_),
    .A(net1416),
    .Y(_3085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5692_ (.Y(_3086_),
    .A(_3077_),
    .B(_3085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5693_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_3074_),
    .A2(_3076_),
    .Y(_3087_),
    .B1(net1426));
 sg13g2_a21oi_1 _5694_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_3082_),
    .A2(_3084_),
    .Y(_3088_),
    .B1(net1416));
 sg13g2_or2_1 _5695_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_3089_),
    .B(_3088_),
    .A(_3087_));
 sg13g2_or4_1 _5696_ (.A(_3051_),
    .B(_3069_),
    .C(_3086_),
    .D(_3089_),
    .X(_3090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5697_ (.B1(_3085_),
    .VDD(VPWR),
    .Y(_3091_),
    .VSS(VGND),
    .A1(_3077_),
    .A2(_3088_));
 sg13g2_nand2b_1 _5698_ (.Y(_3092_),
    .B(_3091_),
    .A_N(_3069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5699_ (.B1(_3011_),
    .VDD(VPWR),
    .Y(_0296_),
    .VSS(VGND),
    .A1(_3066_),
    .A2(_3068_));
 sg13g2_nor2b_1 _5700_ (.A(_0296_),
    .B_N(_3092_),
    .Y(_0297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5701_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0298_),
    .B(net1329),
    .A(net330));
 sg13g2_a21oi_1 _5702_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_3090_),
    .A2(_0297_),
    .Y(_0016_),
    .B1(_0298_));
 sg13g2_and2_1 _5703_ (.A(net1303),
    .B(\s0.data_out[21][0] ),
    .X(_0299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5704_ (.B1(net1317),
    .VDD(VPWR),
    .Y(_0300_),
    .VSS(VGND),
    .A1(_3026_),
    .A2(_0299_));
 sg13g2_a21oi_1 _5705_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1011),
    .A2(_3024_),
    .Y(_0301_),
    .B1(net1341));
 sg13g2_a22oi_1 _5706_ (.Y(_0017_),
    .B1(_0300_),
    .B2(_0301_),
    .A2(_2777_),
    .A1(net1342),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5707_ (.A(net1007),
    .B(_2782_),
    .Y(_0302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5708_ (.B1(net1316),
    .VDD(VPWR),
    .Y(_0303_),
    .VSS(VGND),
    .A1(_3019_),
    .A2(_0302_));
 sg13g2_nor2_1 _5709_ (.A(net1342),
    .B(_3022_),
    .Y(_0304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5710_ (.Y(_0018_),
    .B1(_0303_),
    .B2(_0304_),
    .A2(_2775_),
    .A1(net1342),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5711_ (.A(net1304),
    .B(\s0.data_out[21][2] ),
    .X(_0305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5712_ (.B1(net1316),
    .VDD(VPWR),
    .Y(_0306_),
    .VSS(VGND),
    .A1(_3041_),
    .A2(_0305_));
 sg13g2_nand3_1 _5713_ (.B(_3044_),
    .C(_0306_),
    .A(net1476),
    .Y(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5714_ (.B1(_0307_),
    .VDD(VPWR),
    .Y(_0308_),
    .VSS(VGND),
    .A1(net1463),
    .A2(net646));
 sg13g2_inv_1 _5715_ (.VDD(VPWR),
    .Y(_0019_),
    .A(_0308_),
    .VSS(VGND));
 sg13g2_nor2_1 _5716_ (.A(net1007),
    .B(_2781_),
    .Y(_0309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5717_ (.B1(net1316),
    .VDD(VPWR),
    .Y(_0310_),
    .VSS(VGND),
    .A1(_3034_),
    .A2(_0309_));
 sg13g2_nor2_1 _5718_ (.A(net1341),
    .B(_3037_),
    .Y(_0311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5719_ (.Y(_0020_),
    .B1(_0310_),
    .B2(_0311_),
    .A2(_2770_),
    .A1(net1342),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5720_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1304),
    .A2(net609),
    .Y(_0312_),
    .B1(_3070_));
 sg13g2_a21oi_1 _5721_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1011),
    .A2(_3075_),
    .Y(_0313_),
    .B1(net1344));
 sg13g2_o21ai_1 _5722_ (.B1(_0313_),
    .VDD(VPWR),
    .Y(_0314_),
    .VSS(VGND),
    .A1(net1011),
    .A2(_0312_));
 sg13g2_o21ai_1 _5723_ (.B1(_0314_),
    .VDD(VPWR),
    .Y(_0315_),
    .VSS(VGND),
    .A1(net1462),
    .A2(net635));
 sg13g2_inv_1 _5724_ (.VDD(VPWR),
    .Y(_0021_),
    .A(_0315_),
    .VSS(VGND));
 sg13g2_a21oi_1 _5725_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1300),
    .A2(\s0.data_out[21][5] ),
    .Y(_0316_),
    .B1(_3080_));
 sg13g2_a21oi_1 _5726_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1012),
    .A2(_3083_),
    .Y(_0317_),
    .B1(net1340));
 sg13g2_o21ai_1 _5727_ (.B1(_0317_),
    .VDD(VPWR),
    .Y(_0318_),
    .VSS(VGND),
    .A1(net1012),
    .A2(_0316_));
 sg13g2_o21ai_1 _5728_ (.B1(_0318_),
    .VDD(VPWR),
    .Y(_0319_),
    .VSS(VGND),
    .A1(net1463),
    .A2(net564));
 sg13g2_inv_1 _5729_ (.VDD(VPWR),
    .Y(_0022_),
    .A(net565),
    .VSS(VGND));
 sg13g2_nor2_1 _5730_ (.A(net1008),
    .B(_2780_),
    .Y(_0320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5731_ (.B1(net1313),
    .VDD(VPWR),
    .Y(_0321_),
    .VSS(VGND),
    .A1(_3061_),
    .A2(_0320_));
 sg13g2_nor2_1 _5732_ (.A(net1340),
    .B(_3064_),
    .Y(_0322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5733_ (.Y(_0023_),
    .B1(_0321_),
    .B2(_0322_),
    .A2(_2765_),
    .A1(net1340),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5734_ (.A(net1008),
    .B(_2779_),
    .Y(_0323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5735_ (.B1(net1313),
    .VDD(VPWR),
    .Y(_0324_),
    .VSS(VGND),
    .A1(_3054_),
    .A2(_0323_));
 sg13g2_nor2_1 _5736_ (.A(net1343),
    .B(net378),
    .Y(_0325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5737_ (.Y(_0024_),
    .B1(net528),
    .B2(_0325_),
    .A2(_2763_),
    .A1(net1340),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5738_ (.B1(net1301),
    .VDD(VPWR),
    .Y(_0326_),
    .VSS(VGND),
    .A1(net1393),
    .A2(net1286));
 sg13g2_nor2_1 _5739_ (.A(net1393),
    .B(_2753_),
    .Y(_0327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5740_ (.A(_0326_),
    .B(_0327_),
    .Y(_0328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5741_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1336),
    .A2(net1308),
    .Y(_0329_),
    .B1(net1301));
 sg13g2_nor2_1 _5742_ (.A(_0328_),
    .B(_0329_),
    .Y(_0330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5743_ (.Y(_0331_),
    .B(_0330_),
    .A_N(net698),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5744_ (.B1(_0328_),
    .VDD(VPWR),
    .Y(_0332_),
    .VSS(VGND),
    .A1(net649),
    .A2(net1296));
 sg13g2_or2_1 _5745_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0333_),
    .B(_0326_),
    .A(net1286));
 sg13g2_o21ai_1 _5746_ (.B1(net1008),
    .VDD(VPWR),
    .Y(_0334_),
    .VSS(VGND),
    .A1(net649),
    .A2(net1308));
 sg13g2_nand3_1 _5747_ (.B(_0333_),
    .C(_0334_),
    .A(_0332_),
    .Y(_0335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5748_ (.X(_0025_),
    .A(net1462),
    .B(_0331_),
    .C(_0335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5749_ (.A(net1344),
    .B(_0328_),
    .C(_0329_),
    .Y(_0026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5750_ (.A(net1472),
    .B(net338),
    .X(_0027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5751_ (.Y(_0336_),
    .A(net1297),
    .B(net633),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5752_ (.A0(\s0.data_out[21][1] ),
    .A1(\s0.data_out[20][1] ),
    .S(net1297),
    .X(_0337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5753_ (.A(net1290),
    .B_N(net1166),
    .Y(_0338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5754_ (.A2(_0337_),
    .A1(net1290),
    .B1(_0338_),
    .X(_0339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5755_ (.Y(_0340_),
    .B(\s0.data_out[20][1] ),
    .A_N(net1309),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5756_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_3017_),
    .A2(_0340_),
    .Y(_0341_),
    .B1(net1306));
 sg13g2_a21oi_1 _5757_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1305),
    .A2(_0339_),
    .Y(_0342_),
    .B1(_0341_));
 sg13g2_mux2_1 _5758_ (.A0(\s0.data_out[20][0] ),
    .A1(\s0.data_out[21][0] ),
    .S(net1309),
    .X(_0343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5759_ (.Y(_0344_),
    .A(net1007),
    .B(_0343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5760_ (.A(net1290),
    .B_N(net1170),
    .Y(_0345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5761_ (.A0(\s0.data_out[21][0] ),
    .A1(\s0.data_out[20][0] ),
    .S(net1297),
    .X(_0346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5762_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1290),
    .A2(_0346_),
    .Y(_0347_),
    .B1(_0345_));
 sg13g2_nand2b_1 _5763_ (.Y(_0348_),
    .B(net1305),
    .A_N(_0347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5764_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0348_),
    .C1(net1461),
    .B1(_0344_),
    .A1(net1451),
    .Y(_0349_),
    .A2(_0342_));
 sg13g2_nor2b_1 _5765_ (.A(net1291),
    .B_N(net1163),
    .Y(_0350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5766_ (.Y(_0351_),
    .A(net1298),
    .B(net424),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5767_ (.A0(\s0.data_out[21][2] ),
    .A1(\s0.data_out[20][2] ),
    .S(net1297),
    .X(_0352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5768_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1291),
    .A2(_0352_),
    .Y(_0353_),
    .B1(_0350_));
 sg13g2_mux2_1 _5769_ (.A0(\s0.data_out[20][2] ),
    .A1(\s0.data_out[21][2] ),
    .S(net1309),
    .X(_0354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5770_ (.Y(_0355_),
    .A(net1007),
    .B(_0354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5771_ (.B1(_0355_),
    .VDD(VPWR),
    .Y(_0356_),
    .VSS(VGND),
    .A1(net1007),
    .A2(_0353_));
 sg13g2_or2_1 _5772_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0357_),
    .B(_0356_),
    .A(net1334));
 sg13g2_xnor2_1 _5773_ (.Y(_0358_),
    .A(net1334),
    .B(_0356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5774_ (.Y(_0359_),
    .A(net1297),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5775_ (.A0(\s0.data_out[21][3] ),
    .A1(\s0.data_out[20][3] ),
    .S(net1297),
    .X(_0360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5776_ (.A(net1290),
    .B_N(net1161),
    .Y(_0361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5777_ (.A2(_0360_),
    .A1(net1290),
    .B1(_0361_),
    .X(_0362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5778_ (.Y(_0363_),
    .B(\s0.data_out[20][3] ),
    .A_N(net1309),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5779_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_3032_),
    .A2(_0363_),
    .Y(_0364_),
    .B1(net1305));
 sg13g2_a21oi_1 _5780_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1305),
    .A2(_0362_),
    .Y(_0365_),
    .B1(_0364_));
 sg13g2_nor2_1 _5781_ (.A(net1437),
    .B(_0365_),
    .Y(_0366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5782_ (.A(net1451),
    .B(_0342_),
    .Y(_0367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _5783_ (.A(_0349_),
    .B(_0358_),
    .C(_0366_),
    .D(_0367_),
    .Y(_0368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5784_ (.Y(_0369_),
    .A(net1437),
    .B(_0365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5785_ (.B1(_0369_),
    .VDD(VPWR),
    .Y(_0370_),
    .VSS(VGND),
    .A1(_0357_),
    .A2(_0366_));
 sg13g2_nor2_1 _5786_ (.A(_0368_),
    .B(_0370_),
    .Y(_0371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5787_ (.Y(_0372_),
    .A(net1296),
    .B(net473),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5788_ (.A0(\s0.data_out[21][7] ),
    .A1(\s0.data_out[20][7] ),
    .S(net1296),
    .X(_0373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5789_ (.A(net1286),
    .B_N(net1142),
    .Y(_0374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5790_ (.A2(_0373_),
    .A1(net1286),
    .B1(_0374_),
    .X(_0375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5791_ (.Y(_0376_),
    .B(net473),
    .A_N(net1308),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5792_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_3052_),
    .A2(_0376_),
    .Y(_0377_),
    .B1(net1301));
 sg13g2_a21oi_1 _5793_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1301),
    .A2(_0375_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_nand2_1 _5794_ (.Y(_0379_),
    .A(net1296),
    .B(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5795_ (.A0(\s0.data_out[21][6] ),
    .A1(\s0.data_out[20][6] ),
    .S(net1296),
    .X(_0380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5796_ (.A(net1286),
    .B_N(net1147),
    .Y(_0381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5797_ (.A2(_0380_),
    .A1(net1286),
    .B1(_0381_),
    .X(_0382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5798_ (.Y(_0383_),
    .B(net432),
    .A_N(net1308),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5799_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_3059_),
    .A2(_0383_),
    .Y(_0384_),
    .B1(net1301));
 sg13g2_a21oi_1 _5800_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1301),
    .A2(_0382_),
    .Y(_0385_),
    .B1(_0384_));
 sg13g2_a22oi_1 _5801_ (.Y(_0386_),
    .B1(_0385_),
    .B2(net1407),
    .A2(_0378_),
    .A1(net1398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5802_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0387_),
    .B(_0385_),
    .A(net1407));
 sg13g2_nor2_1 _5803_ (.A(net1398),
    .B(_0378_),
    .Y(_0388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _5804_ (.B(_0386_),
    .C(_0387_),
    .Y(_0389_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0388_));
 sg13g2_nor2b_1 _5805_ (.A(net1292),
    .B_N(net1157),
    .Y(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5806_ (.Y(_0391_),
    .A(net1298),
    .B(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5807_ (.A0(\s0.data_out[21][4] ),
    .A1(\s0.data_out[20][4] ),
    .S(net1297),
    .X(_0392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5808_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1292),
    .A2(_0392_),
    .Y(_0393_),
    .B1(_0390_));
 sg13g2_nand2b_1 _5809_ (.Y(_0394_),
    .B(net1305),
    .A_N(_0393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5810_ (.B1(_3071_),
    .VDD(VPWR),
    .Y(_0395_),
    .VSS(VGND),
    .A1(net1309),
    .A2(_2787_));
 sg13g2_nand2_1 _5811_ (.Y(_0396_),
    .A(net1007),
    .B(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5812_ (.B(_0394_),
    .C(_0396_),
    .A(net1427),
    .Y(_0397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5813_ (.Y(_0398_),
    .A(net1299),
    .B(\s0.data_out[20][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5814_ (.A0(\s0.data_out[21][5] ),
    .A1(\s0.data_out[20][5] ),
    .S(net1296),
    .X(_0399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5815_ (.A(net1289),
    .B_N(net1151),
    .Y(_0400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5816_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1289),
    .A2(_0399_),
    .Y(_0401_),
    .B1(_0400_));
 sg13g2_nand2b_1 _5817_ (.Y(_0402_),
    .B(net1302),
    .A_N(_0401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5818_ (.B1(_3078_),
    .VDD(VPWR),
    .Y(_0403_),
    .VSS(VGND),
    .A1(net1308),
    .A2(_2786_));
 sg13g2_nand2_1 _5819_ (.Y(_0404_),
    .A(net1008),
    .B(_0403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5820_ (.B(_0402_),
    .C(_0404_),
    .A(net1418),
    .Y(_0405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5821_ (.Y(_0406_),
    .A(_0397_),
    .B(_0405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5822_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0394_),
    .A2(_0396_),
    .Y(_0407_),
    .B1(net1427));
 sg13g2_a21oi_1 _5823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0402_),
    .A2(_0404_),
    .Y(_0408_),
    .B1(net1418));
 sg13g2_or2_1 _5824_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0409_),
    .B(_0408_),
    .A(_0407_));
 sg13g2_or4_1 _5825_ (.A(_0371_),
    .B(_0389_),
    .C(_0406_),
    .D(_0409_),
    .X(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5826_ (.B1(_0405_),
    .VDD(VPWR),
    .Y(_0411_),
    .VSS(VGND),
    .A1(_0397_),
    .A2(_0408_));
 sg13g2_nor2b_1 _5827_ (.A(_0389_),
    .B_N(_0411_),
    .Y(_0412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5828_ (.B1(_0330_),
    .VDD(VPWR),
    .Y(_0413_),
    .VSS(VGND),
    .A1(_0386_),
    .A2(_0388_));
 sg13g2_nor2_1 _5829_ (.A(_0412_),
    .B(_0413_),
    .Y(_0414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5830_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0415_),
    .B(net1329),
    .A(net332));
 sg13g2_a21oi_1 _5831_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0410_),
    .A2(_0414_),
    .Y(_0028_),
    .B1(_0415_));
 sg13g2_and2_1 _5832_ (.A(net1291),
    .B(\s0.data_out[20][0] ),
    .X(_0416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5833_ (.B1(net1305),
    .VDD(VPWR),
    .Y(_0417_),
    .VSS(VGND),
    .A1(_0345_),
    .A2(_0416_));
 sg13g2_nand3_1 _5834_ (.B(_0344_),
    .C(_0417_),
    .A(net1462),
    .Y(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5835_ (.B1(_0418_),
    .VDD(VPWR),
    .Y(_0419_),
    .VSS(VGND),
    .A1(net1463),
    .A2(net648));
 sg13g2_inv_1 _5836_ (.VDD(VPWR),
    .Y(_0029_),
    .A(_0419_),
    .VSS(VGND));
 sg13g2_and2_1 _5837_ (.A(net1290),
    .B(\s0.data_out[20][1] ),
    .X(_0420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5838_ (.B1(net1306),
    .VDD(VPWR),
    .Y(_0421_),
    .VSS(VGND),
    .A1(_0338_),
    .A2(_0420_));
 sg13g2_nor2_1 _5839_ (.A(net1345),
    .B(_0341_),
    .Y(_0422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5840_ (.Y(_0030_),
    .B1(_0421_),
    .B2(_0422_),
    .A2(_2782_),
    .A1(net1345),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5841_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1291),
    .A2(net424),
    .Y(_0423_),
    .B1(_0350_));
 sg13g2_a21oi_1 _5842_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1007),
    .A2(_0354_),
    .Y(_0424_),
    .B1(net1345));
 sg13g2_o21ai_1 _5843_ (.B1(_0424_),
    .VDD(VPWR),
    .Y(_0425_),
    .VSS(VGND),
    .A1(net1007),
    .A2(_0423_));
 sg13g2_o21ai_1 _5844_ (.B1(_0425_),
    .VDD(VPWR),
    .Y(_0426_),
    .VSS(VGND),
    .A1(net1462),
    .A2(net624));
 sg13g2_inv_1 _5845_ (.VDD(VPWR),
    .Y(_0031_),
    .A(_0426_),
    .VSS(VGND));
 sg13g2_and2_1 _5846_ (.A(net1290),
    .B(\s0.data_out[20][3] ),
    .X(_0427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5847_ (.B1(net1305),
    .VDD(VPWR),
    .Y(_0428_),
    .VSS(VGND),
    .A1(_0361_),
    .A2(_0427_));
 sg13g2_nor2_1 _5848_ (.A(net1345),
    .B(_0364_),
    .Y(_0429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5849_ (.Y(_0032_),
    .B1(_0428_),
    .B2(_0429_),
    .A2(_2781_),
    .A1(net1345),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1292),
    .A2(net496),
    .Y(_0430_),
    .B1(_0390_));
 sg13g2_a21oi_1 _5851_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1008),
    .A2(_0395_),
    .Y(_0431_),
    .B1(net1344));
 sg13g2_o21ai_1 _5852_ (.B1(_0431_),
    .VDD(VPWR),
    .Y(_0432_),
    .VSS(VGND),
    .A1(_2752_),
    .A2(_0430_));
 sg13g2_o21ai_1 _5853_ (.B1(_0432_),
    .VDD(VPWR),
    .Y(_0433_),
    .VSS(VGND),
    .A1(net1462),
    .A2(net609));
 sg13g2_inv_1 _5854_ (.VDD(VPWR),
    .Y(_0033_),
    .A(_0433_),
    .VSS(VGND));
 sg13g2_a21oi_1 _5855_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1289),
    .A2(net468),
    .Y(_0434_),
    .B1(_0400_));
 sg13g2_a21oi_1 _5856_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1008),
    .A2(_0403_),
    .Y(_0435_),
    .B1(net1344));
 sg13g2_o21ai_1 _5857_ (.B1(_0435_),
    .VDD(VPWR),
    .Y(_0436_),
    .VSS(VGND),
    .A1(net1008),
    .A2(_0434_));
 sg13g2_o21ai_1 _5858_ (.B1(_0436_),
    .VDD(VPWR),
    .Y(_0437_),
    .VSS(VGND),
    .A1(net1462),
    .A2(net659));
 sg13g2_inv_1 _5859_ (.VDD(VPWR),
    .Y(_0034_),
    .A(_0437_),
    .VSS(VGND));
 sg13g2_and2_1 _5860_ (.A(net1286),
    .B(net432),
    .X(_0438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5861_ (.B1(net1301),
    .VDD(VPWR),
    .Y(_0439_),
    .VSS(VGND),
    .A1(_0381_),
    .A2(_0438_));
 sg13g2_nor2_1 _5862_ (.A(net1344),
    .B(_0384_),
    .Y(_0440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5863_ (.Y(_0035_),
    .B1(_0439_),
    .B2(_0440_),
    .A2(_2780_),
    .A1(net1344),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5864_ (.A(net1286),
    .B(net473),
    .X(_0441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5865_ (.B1(net1301),
    .VDD(VPWR),
    .Y(_0442_),
    .VSS(VGND),
    .A1(_0374_),
    .A2(_0441_));
 sg13g2_nor2_1 _5866_ (.A(net1344),
    .B(_0377_),
    .Y(_0443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5867_ (.Y(_0036_),
    .B1(_0442_),
    .B2(_0443_),
    .A2(_2779_),
    .A1(net1344),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5868_ (.B1(net1287),
    .VDD(VPWR),
    .Y(_0444_),
    .VSS(VGND),
    .A1(net1393),
    .A2(net1273));
 sg13g2_nand2_1 _5869_ (.Y(_0445_),
    .A(net1336),
    .B(net1282),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5870_ (.Y(_0446_),
    .B(_0445_),
    .A_N(_0444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5871_ (.B1(_0446_),
    .VDD(VPWR),
    .Y(_0447_),
    .VSS(VGND),
    .A1(net1287),
    .A2(_0327_));
 sg13g2_nor2_1 _5872_ (.A(net366),
    .B(net1281),
    .Y(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5873_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0449_),
    .B(_0448_),
    .A(_0446_));
 sg13g2_nor2_1 _5874_ (.A(net1273),
    .B(_0444_),
    .Y(_0450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5875_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2738_),
    .A2(_2753_),
    .Y(_0451_),
    .B1(net1288));
 sg13g2_nor2_1 _5876_ (.A(_0450_),
    .B(_0451_),
    .Y(_0452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5877_ (.B1(net1472),
    .VDD(VPWR),
    .Y(_0453_),
    .VSS(VGND),
    .A1(net649),
    .A2(_0447_));
 sg13g2_a21oi_1 _5878_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0449_),
    .A2(_0452_),
    .Y(_0037_),
    .B1(_0453_));
 sg13g2_nor2_1 _5879_ (.A(net1352),
    .B(_0447_),
    .Y(_0038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5880_ (.A(net1466),
    .B(net325),
    .X(_0039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5881_ (.Y(_0454_),
    .A(net1284),
    .B(net657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5882_ (.A0(\s0.data_out[20][2] ),
    .A1(\s0.data_out[19][2] ),
    .S(net1283),
    .X(_0455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5883_ (.A(net1276),
    .B_N(net1162),
    .Y(_0456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5884_ (.A2(_0455_),
    .A1(net1276),
    .B1(_0456_),
    .X(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5885_ (.Y(_0458_),
    .B(\s0.data_out[19][2] ),
    .A_N(net1298),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5886_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0351_),
    .A2(_0458_),
    .Y(_0459_),
    .B1(net1293));
 sg13g2_a21oi_1 _5887_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1293),
    .A2(_0457_),
    .Y(_0460_),
    .B1(_0459_));
 sg13g2_or2_1 _5888_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0461_),
    .B(_0460_),
    .A(net1444));
 sg13g2_nand2_1 _5889_ (.Y(_0462_),
    .A(net1284),
    .B(net695),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5890_ (.B1(_0462_),
    .VDD(VPWR),
    .Y(_0463_),
    .VSS(VGND),
    .A1(net1283),
    .A2(_2790_));
 sg13g2_nor2b_1 _5891_ (.A(net1277),
    .B_N(net1166),
    .Y(_0464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5892_ (.A2(_0463_),
    .A1(net1276),
    .B1(_0464_),
    .X(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5893_ (.Y(_0466_),
    .A(_2753_),
    .B(\s0.data_out[19][1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5894_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0336_),
    .A2(_0466_),
    .Y(_0467_),
    .B1(net1294));
 sg13g2_a21oi_1 _5895_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1294),
    .A2(_0465_),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_mux2_1 _5896_ (.A0(\s0.data_out[20][0] ),
    .A1(\s0.data_out[19][0] ),
    .S(net1283),
    .X(_0469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5897_ (.A(net1276),
    .B_N(net1173),
    .Y(_0470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5898_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1276),
    .A2(_0469_),
    .Y(_0471_),
    .B1(_0470_));
 sg13g2_nand2b_1 _5899_ (.Y(_0472_),
    .B(net1293),
    .A_N(_0471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5900_ (.A0(\s0.data_out[19][0] ),
    .A1(\s0.data_out[20][0] ),
    .S(net1298),
    .X(_0473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5901_ (.Y(_0474_),
    .B(_0473_),
    .A_N(net1293),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5902_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0474_),
    .C1(net1461),
    .B1(_0472_),
    .A1(net1451),
    .Y(_0475_),
    .A2(_0468_));
 sg13g2_o21ai_1 _5903_ (.B1(_0461_),
    .VDD(VPWR),
    .Y(_0476_),
    .VSS(VGND),
    .A1(net1451),
    .A2(_0468_));
 sg13g2_nand2_1 _5904_ (.Y(_0477_),
    .A(net1284),
    .B(net690),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5905_ (.B1(_0477_),
    .VDD(VPWR),
    .Y(_0478_),
    .VSS(VGND),
    .A1(net1283),
    .A2(_2788_));
 sg13g2_nor2_1 _5906_ (.A(net1276),
    .B(net993),
    .Y(_0479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5907_ (.A2(_0478_),
    .A1(net1276),
    .B1(_0479_),
    .X(_0480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5908_ (.Y(_0481_),
    .A(_2753_),
    .B(\s0.data_out[19][3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5909_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0359_),
    .A2(_0481_),
    .Y(_0482_),
    .B1(net1293));
 sg13g2_a21oi_1 _5910_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1294),
    .A2(_0480_),
    .Y(_0483_),
    .B1(_0482_));
 sg13g2_a22oi_1 _5911_ (.Y(_0484_),
    .B1(_0483_),
    .B2(net1437),
    .A2(_0460_),
    .A1(net1444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5912_ (.B1(_0484_),
    .VDD(VPWR),
    .Y(_0485_),
    .VSS(VGND),
    .A1(_0475_),
    .A2(_0476_));
 sg13g2_nand2_1 _5913_ (.Y(_0486_),
    .A(net1282),
    .B(net506),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5914_ (.A0(\s0.data_out[20][7] ),
    .A1(\s0.data_out[19][7] ),
    .S(net1281),
    .X(_0487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5915_ (.A(net1273),
    .B_N(net1143),
    .Y(_0488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5916_ (.A2(_0487_),
    .A1(net1273),
    .B1(_0488_),
    .X(_0489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5917_ (.Y(_0490_),
    .B(\s0.data_out[19][7] ),
    .A_N(net1296),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5918_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0372_),
    .A2(_0490_),
    .Y(_0491_),
    .B1(net1287));
 sg13g2_a21oi_1 _5919_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1287),
    .A2(_0489_),
    .Y(_0492_),
    .B1(_0491_));
 sg13g2_nand2_1 _5920_ (.Y(_0493_),
    .A(net1282),
    .B(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5921_ (.A0(\s0.data_out[20][6] ),
    .A1(\s0.data_out[19][6] ),
    .S(net1281),
    .X(_0494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5922_ (.A(net1273),
    .B_N(net1148),
    .Y(_0495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5923_ (.A2(_0494_),
    .A1(net1273),
    .B1(_0495_),
    .X(_0496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5924_ (.Y(_0497_),
    .B(\s0.data_out[19][6] ),
    .A_N(net1296),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5925_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0379_),
    .A2(_0497_),
    .Y(_0498_),
    .B1(net1287));
 sg13g2_a21oi_1 _5926_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1287),
    .A2(_0496_),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_a22oi_1 _5927_ (.Y(_0500_),
    .B1(_0499_),
    .B2(net1409),
    .A2(_0492_),
    .A1(net1400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5928_ (.VDD(VPWR),
    .Y(_0501_),
    .A(_0500_),
    .VSS(VGND));
 sg13g2_or2_1 _5929_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0502_),
    .B(_0492_),
    .A(net1400));
 sg13g2_o21ai_1 _5930_ (.B1(_0502_),
    .VDD(VPWR),
    .Y(_0503_),
    .VSS(VGND),
    .A1(net1409),
    .A2(_0499_));
 sg13g2_nor2_1 _5931_ (.A(_0501_),
    .B(_0503_),
    .Y(_0504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5932_ (.Y(_0505_),
    .A(net1283),
    .B(net486),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5933_ (.B1(_0505_),
    .VDD(VPWR),
    .Y(_0506_),
    .VSS(VGND),
    .A1(net1283),
    .A2(_2787_));
 sg13g2_nor2b_1 _5934_ (.A(net1277),
    .B_N(net1156),
    .Y(_0507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5935_ (.A2(_0506_),
    .A1(net1277),
    .B1(_0507_),
    .X(_0508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5936_ (.Y(_0509_),
    .A(_2753_),
    .B(net486),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5937_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0391_),
    .A2(_0509_),
    .Y(_0510_),
    .B1(net1295));
 sg13g2_a21oi_1 _5938_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1295),
    .A2(_0508_),
    .Y(_0511_),
    .B1(_0510_));
 sg13g2_nand2_1 _5939_ (.Y(_0512_),
    .A(net1281),
    .B(net352),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5940_ (.B1(_0512_),
    .VDD(VPWR),
    .Y(_0513_),
    .VSS(VGND),
    .A1(net1281),
    .A2(_2786_));
 sg13g2_nor2b_1 _5941_ (.A(net1275),
    .B_N(net1152),
    .Y(_0514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5942_ (.A2(_0513_),
    .A1(net1273),
    .B1(_0514_),
    .X(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5943_ (.Y(_0516_),
    .A(_2753_),
    .B(net352),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5944_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0398_),
    .A2(_0516_),
    .Y(_0517_),
    .B1(net1288));
 sg13g2_a21oi_1 _5945_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1288),
    .A2(_0515_),
    .Y(_0518_),
    .B1(_0517_));
 sg13g2_a22oi_1 _5946_ (.Y(_0519_),
    .B1(_0518_),
    .B2(net1418),
    .A2(_0511_),
    .A1(net1427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5947_ (.A(net1437),
    .B(_0483_),
    .Y(_0520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5948_ (.A(net1418),
    .B(_0518_),
    .Y(_0521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5949_ (.A(net1427),
    .B(_0511_),
    .Y(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5950_ (.A(_0520_),
    .B(_0521_),
    .C(_0522_),
    .Y(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5951_ (.B(_0504_),
    .C(_0519_),
    .A(_0485_),
    .Y(_0524_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0523_));
 sg13g2_nor2_1 _5952_ (.A(_0519_),
    .B(_0521_),
    .Y(_0525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5953_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0525_),
    .C1(_0447_),
    .B1(_0504_),
    .A1(_0501_),
    .Y(_0526_),
    .A2(_0502_));
 sg13g2_or2_1 _5954_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0527_),
    .B(net1329),
    .A(net338));
 sg13g2_a21oi_1 _5955_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0524_),
    .A2(_0526_),
    .Y(_0040_),
    .B1(_0527_));
 sg13g2_and2_1 _5956_ (.A(net1276),
    .B(\s0.data_out[19][0] ),
    .X(_0528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5957_ (.B1(net1293),
    .VDD(VPWR),
    .Y(_0529_),
    .VSS(VGND),
    .A1(_0470_),
    .A2(_0528_));
 sg13g2_nand3_1 _5958_ (.B(_0474_),
    .C(_0529_),
    .A(net1472),
    .Y(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5959_ (.B1(_0530_),
    .VDD(VPWR),
    .Y(_0531_),
    .VSS(VGND),
    .A1(net1472),
    .A2(net672));
 sg13g2_inv_1 _5960_ (.VDD(VPWR),
    .Y(_0041_),
    .A(_0531_),
    .VSS(VGND));
 sg13g2_nor2_1 _5961_ (.A(net1003),
    .B(_2796_),
    .Y(_0532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5962_ (.B1(net1294),
    .VDD(VPWR),
    .Y(_0533_),
    .VSS(VGND),
    .A1(_0464_),
    .A2(_0532_));
 sg13g2_nor2_1 _5963_ (.A(net1354),
    .B(_0467_),
    .Y(_0534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5964_ (.Y(_0042_),
    .B1(_0533_),
    .B2(_0534_),
    .A2(_2790_),
    .A1(net1354),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5965_ (.A(net1003),
    .B(_2795_),
    .Y(_0535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5966_ (.B1(net1293),
    .VDD(VPWR),
    .Y(_0536_),
    .VSS(VGND),
    .A1(_0456_),
    .A2(_0535_));
 sg13g2_nor2_1 _5967_ (.A(net1354),
    .B(_0459_),
    .Y(_0537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5968_ (.Y(_0043_),
    .B1(_0536_),
    .B2(_0537_),
    .A2(_2789_),
    .A1(net1354),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5969_ (.A(_2755_),
    .B(_2794_),
    .Y(_0538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5970_ (.B1(net1293),
    .VDD(VPWR),
    .Y(_0539_),
    .VSS(VGND),
    .A1(_0479_),
    .A2(_0538_));
 sg13g2_nor2_1 _5971_ (.A(net1354),
    .B(_0482_),
    .Y(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5972_ (.Y(_0044_),
    .B1(_0539_),
    .B2(_0540_),
    .A2(_2788_),
    .A1(net1354),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5973_ (.A(_2755_),
    .B(_2793_),
    .Y(_0541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5974_ (.B1(net1295),
    .VDD(VPWR),
    .Y(_0542_),
    .VSS(VGND),
    .A1(_0507_),
    .A2(_0541_));
 sg13g2_nor2_1 _5975_ (.A(net1352),
    .B(_0510_),
    .Y(_0543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5976_ (.Y(_0045_),
    .B1(_0542_),
    .B2(_0543_),
    .A2(_2787_),
    .A1(net1352),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5977_ (.A(net1003),
    .B(_2792_),
    .Y(_0544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5978_ (.B1(net1288),
    .VDD(VPWR),
    .Y(_0545_),
    .VSS(VGND),
    .A1(_0514_),
    .A2(_0544_));
 sg13g2_nor2_1 _5979_ (.A(net1352),
    .B(net353),
    .Y(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5980_ (.Y(_0046_),
    .B1(_0545_),
    .B2(_0546_),
    .A2(_2786_),
    .A1(net1352),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5981_ (.A(net1273),
    .B(\s0.data_out[19][6] ),
    .X(_0547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5982_ (.B1(net1287),
    .VDD(VPWR),
    .Y(_0548_),
    .VSS(VGND),
    .A1(_0495_),
    .A2(_0547_));
 sg13g2_nor2_1 _5983_ (.A(net1352),
    .B(_0498_),
    .Y(_0549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5984_ (.Y(_0047_),
    .B1(_0548_),
    .B2(_0549_),
    .A2(_2785_),
    .A1(net1352),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5985_ (.A(net1003),
    .B(_2791_),
    .Y(_0550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5986_ (.B1(net1287),
    .VDD(VPWR),
    .Y(_0551_),
    .VSS(VGND),
    .A1(_0488_),
    .A2(_0550_));
 sg13g2_nor2_1 _5987_ (.A(net1353),
    .B(_0491_),
    .Y(_0552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5988_ (.Y(_0048_),
    .B1(_0551_),
    .B2(_0552_),
    .A2(_2784_),
    .A1(net1353),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5989_ (.B1(net1274),
    .VDD(VPWR),
    .Y(_0553_),
    .VSS(VGND),
    .A1(net1393),
    .A2(net1261));
 sg13g2_nor2_1 _5990_ (.A(net1394),
    .B(_2756_),
    .Y(_0554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5991_ (.A(_0553_),
    .B(_0554_),
    .Y(_0555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5992_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1003),
    .A2(_0445_),
    .Y(_0556_),
    .B1(_0555_));
 sg13g2_o21ai_1 _5993_ (.B1(_0555_),
    .VDD(VPWR),
    .Y(_0557_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[18] [0]),
    .A2(net1269));
 sg13g2_nor2_1 _5994_ (.A(net1261),
    .B(_0553_),
    .Y(_0558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5995_ (.B1(net1003),
    .VDD(VPWR),
    .Y(_0559_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[18] [0]),
    .A2(net1281));
 sg13g2_nand2_1 _5996_ (.Y(_0560_),
    .A(_0557_),
    .B(_0559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5997_ (.B1(net1470),
    .VDD(VPWR),
    .Y(_0561_),
    .VSS(VGND),
    .A1(_0558_),
    .A2(_0560_));
 sg13g2_a21oi_1 _5998_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2738_),
    .A2(_0556_),
    .Y(_0049_),
    .B1(_0561_));
 sg13g2_and2_1 _5999_ (.A(net1470),
    .B(_0556_),
    .X(_0050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6000_ (.A(net1470),
    .B(net337),
    .X(_0051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6001_ (.Y(_0562_),
    .A(net1271),
    .B(net428),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6002_ (.A0(\s0.data_out[19][2] ),
    .A1(\s0.data_out[18][2] ),
    .S(net1270),
    .X(_0563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6003_ (.A(net1266),
    .B_N(net1162),
    .Y(_0564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6004_ (.A2(_0563_),
    .A1(net1265),
    .B1(_0564_),
    .X(_0565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6005_ (.Y(_0566_),
    .B(net428),
    .A_N(net1283),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6006_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0454_),
    .A2(_0566_),
    .Y(_0567_),
    .B1(net1278));
 sg13g2_a21oi_1 _6007_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1278),
    .A2(_0565_),
    .Y(_0568_),
    .B1(_0567_));
 sg13g2_or2_1 _6008_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0569_),
    .B(_0568_),
    .A(net1443));
 sg13g2_nand2_1 _6009_ (.Y(_0570_),
    .A(net1271),
    .B(net418),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6010_ (.B1(_0570_),
    .VDD(VPWR),
    .Y(_0571_),
    .VSS(VGND),
    .A1(net1270),
    .A2(_2796_));
 sg13g2_nor2b_1 _6011_ (.A(net1265),
    .B_N(net1167),
    .Y(_0572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6012_ (.A2(_0571_),
    .A1(net1266),
    .B1(_0572_),
    .X(_0573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6013_ (.Y(_0574_),
    .B(net418),
    .A_N(net1283),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6014_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0462_),
    .A2(_0574_),
    .Y(_0575_),
    .B1(net1279));
 sg13g2_a21oi_1 _6015_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1278),
    .A2(_0573_),
    .Y(_0576_),
    .B1(_0575_));
 sg13g2_mux2_1 _6016_ (.A0(\s0.data_out[19][0] ),
    .A1(\s0.data_out[18][0] ),
    .S(net1270),
    .X(_0577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6017_ (.A(net1265),
    .B_N(net1173),
    .Y(_0578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6018_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1265),
    .A2(_0577_),
    .Y(_0579_),
    .B1(_0578_));
 sg13g2_nand2b_1 _6019_ (.Y(_0580_),
    .B(net1278),
    .A_N(_0579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6020_ (.A0(\s0.data_out[18][0] ),
    .A1(\s0.data_out[19][0] ),
    .S(net1284),
    .X(_0581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6021_ (.Y(_0582_),
    .A(net1003),
    .B(_0581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _6022_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0582_),
    .C1(net1460),
    .B1(_0580_),
    .A1(net1452),
    .Y(_0583_),
    .A2(_0576_));
 sg13g2_o21ai_1 _6023_ (.B1(_0569_),
    .VDD(VPWR),
    .Y(_0584_),
    .VSS(VGND),
    .A1(net1452),
    .A2(_0576_));
 sg13g2_nand2_1 _6024_ (.Y(_0585_),
    .A(net1270),
    .B(net410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6025_ (.B1(_0585_),
    .VDD(VPWR),
    .Y(_0586_),
    .VSS(VGND),
    .A1(net1270),
    .A2(_2794_));
 sg13g2_nor2_1 _6026_ (.A(net1265),
    .B(net993),
    .Y(_0587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6027_ (.A2(_0586_),
    .A1(net1265),
    .B1(_0587_),
    .X(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6028_ (.Y(_0589_),
    .B(net410),
    .A_N(net1284),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6029_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0477_),
    .A2(_0589_),
    .Y(_0590_),
    .B1(net1278));
 sg13g2_a21oi_1 _6030_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1279),
    .A2(_0588_),
    .Y(_0591_),
    .B1(_0590_));
 sg13g2_a22oi_1 _6031_ (.Y(_0592_),
    .B1(_0591_),
    .B2(net1437),
    .A2(_0568_),
    .A1(net1444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6032_ (.B1(_0592_),
    .VDD(VPWR),
    .Y(_0593_),
    .VSS(VGND),
    .A1(_0583_),
    .A2(_0584_));
 sg13g2_nand2_1 _6033_ (.Y(_0594_),
    .A(net1269),
    .B(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6034_ (.A0(\s0.data_out[19][7] ),
    .A1(\s0.data_out[18][7] ),
    .S(net1269),
    .X(_0595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6035_ (.A(net1261),
    .B_N(net1143),
    .Y(_0596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6036_ (.A2(_0595_),
    .A1(net1261),
    .B1(_0596_),
    .X(_0597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6037_ (.Y(_0598_),
    .B(net499),
    .A_N(net1281),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6038_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0486_),
    .A2(_0598_),
    .Y(_0599_),
    .B1(net1274));
 sg13g2_a21oi_1 _6039_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1274),
    .A2(_0597_),
    .Y(_0600_),
    .B1(_0599_));
 sg13g2_nand2_1 _6040_ (.Y(_0601_),
    .A(net1272),
    .B(net534),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6041_ (.A0(\s0.data_out[19][6] ),
    .A1(\s0.data_out[18][6] ),
    .S(net1269),
    .X(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6042_ (.A(net1261),
    .B_N(net1148),
    .Y(_0603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6043_ (.A2(_0602_),
    .A1(net1261),
    .B1(_0603_),
    .X(_0604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6044_ (.Y(_0605_),
    .B(net534),
    .A_N(net1281),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6045_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0493_),
    .A2(_0605_),
    .Y(_0606_),
    .B1(net1274));
 sg13g2_a21oi_1 _6046_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1274),
    .A2(_0604_),
    .Y(_0607_),
    .B1(_0606_));
 sg13g2_a22oi_1 _6047_ (.Y(_0608_),
    .B1(_0607_),
    .B2(net1409),
    .A2(_0600_),
    .A1(net1400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _6048_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0609_),
    .B(_0607_),
    .A(net1409));
 sg13g2_or2_1 _6049_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0610_),
    .B(_0600_),
    .A(net1400));
 sg13g2_inv_1 _6050_ (.VDD(VPWR),
    .Y(_0611_),
    .A(_0610_),
    .VSS(VGND));
 sg13g2_and3_1 _6051_ (.X(_0612_),
    .A(_0608_),
    .B(_0609_),
    .C(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6052_ (.Y(_0613_),
    .A(net1271),
    .B(net440),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6053_ (.A0(\s0.data_out[19][4] ),
    .A1(\s0.data_out[18][4] ),
    .S(net1270),
    .X(_0614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6054_ (.A(net1266),
    .B_N(net1156),
    .Y(_0615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6055_ (.A2(_0614_),
    .A1(net1266),
    .B1(_0615_),
    .X(_0616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6056_ (.Y(_0617_),
    .B(net440),
    .A_N(net1284),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6057_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0505_),
    .A2(_0617_),
    .Y(_0618_),
    .B1(net1277));
 sg13g2_a21oi_1 _6058_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1278),
    .A2(_0616_),
    .Y(_0619_),
    .B1(_0618_));
 sg13g2_nand2_1 _6059_ (.Y(_0620_),
    .A(net1272),
    .B(\s0.data_out[18][5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6060_ (.A0(\s0.data_out[19][5] ),
    .A1(\s0.data_out[18][5] ),
    .S(net1269),
    .X(_0621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6061_ (.A(net1264),
    .B_N(net1152),
    .Y(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6062_ (.A2(_0621_),
    .A1(net1264),
    .B1(_0622_),
    .X(_0623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6063_ (.Y(_0624_),
    .B(net436),
    .A_N(net1282),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6064_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0512_),
    .A2(_0624_),
    .Y(_0625_),
    .B1(net1275));
 sg13g2_a21oi_1 _6065_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1274),
    .A2(_0623_),
    .Y(_0626_),
    .B1(_0625_));
 sg13g2_a22oi_1 _6066_ (.Y(_0627_),
    .B1(_0626_),
    .B2(net1418),
    .A2(_0619_),
    .A1(net1427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6067_ (.A(net1427),
    .B(_0619_),
    .Y(_0628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _6068_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0629_),
    .B(_0591_),
    .A(net1437));
 sg13g2_nor2_1 _6069_ (.A(net1418),
    .B(_0626_),
    .Y(_0630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6070_ (.A(_0628_),
    .B(_0630_),
    .Y(_0631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _6071_ (.A(_0612_),
    .B(_0627_),
    .C(_0629_),
    .D(_0631_),
    .X(_0632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6072_ (.A(_0627_),
    .B(_0630_),
    .Y(_0633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6073_ (.B1(_0556_),
    .VDD(VPWR),
    .Y(_0634_),
    .VSS(VGND),
    .A1(_0608_),
    .A2(_0611_));
 sg13g2_a221oi_1 _6074_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0612_),
    .C1(_0634_),
    .B1(_0633_),
    .A1(_0593_),
    .Y(_0635_),
    .A2(_0632_));
 sg13g2_nor3_1 _6075_ (.A(net327),
    .B(net1330),
    .C(_0635_),
    .Y(_0052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6076_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1265),
    .A2(\s0.data_out[18][0] ),
    .Y(_0636_),
    .B1(_0578_));
 sg13g2_a21oi_1 _6077_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1003),
    .A2(_0581_),
    .Y(_0637_),
    .B1(net1355));
 sg13g2_o21ai_1 _6078_ (.B1(_0637_),
    .VDD(VPWR),
    .Y(_0638_),
    .VSS(VGND),
    .A1(_2755_),
    .A2(_0636_));
 sg13g2_o21ai_1 _6079_ (.B1(_0638_),
    .VDD(VPWR),
    .Y(_0639_),
    .VSS(VGND),
    .A1(net1471),
    .A2(net597));
 sg13g2_inv_1 _6080_ (.VDD(VPWR),
    .Y(_0053_),
    .A(net598),
    .VSS(VGND));
 sg13g2_and2_1 _6081_ (.A(net1266),
    .B(net418),
    .X(_0640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6082_ (.B1(net1279),
    .VDD(VPWR),
    .Y(_0641_),
    .VSS(VGND),
    .A1(_0572_),
    .A2(_0640_));
 sg13g2_nor2_1 _6083_ (.A(net1355),
    .B(_0575_),
    .Y(_0642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6084_ (.Y(_0054_),
    .B1(_0641_),
    .B2(_0642_),
    .A2(_2796_),
    .A1(net1355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6085_ (.A(net1266),
    .B(net428),
    .X(_0643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6086_ (.B1(net1278),
    .VDD(VPWR),
    .Y(_0644_),
    .VSS(VGND),
    .A1(_0564_),
    .A2(_0643_));
 sg13g2_nor2_1 _6087_ (.A(net1355),
    .B(_0567_),
    .Y(_0645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6088_ (.Y(_0055_),
    .B1(_0644_),
    .B2(_0645_),
    .A2(_2795_),
    .A1(net1355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6089_ (.A(net1265),
    .B(net410),
    .X(_0646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6090_ (.B1(net1279),
    .VDD(VPWR),
    .Y(_0647_),
    .VSS(VGND),
    .A1(_0587_),
    .A2(_0646_));
 sg13g2_nor2_1 _6091_ (.A(net1355),
    .B(_0590_),
    .Y(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6092_ (.Y(_0056_),
    .B1(_0647_),
    .B2(_0648_),
    .A2(_2794_),
    .A1(net1355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6093_ (.A(net1266),
    .B(net440),
    .X(_0649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6094_ (.B1(net1278),
    .VDD(VPWR),
    .Y(_0650_),
    .VSS(VGND),
    .A1(_0615_),
    .A2(_0649_));
 sg13g2_nor2_1 _6095_ (.A(net1352),
    .B(_0618_),
    .Y(_0651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6096_ (.Y(_0057_),
    .B1(_0650_),
    .B2(_0651_),
    .A2(_2793_),
    .A1(net1353),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6097_ (.A(net1264),
    .B(net436),
    .X(_0652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6098_ (.B1(net1275),
    .VDD(VPWR),
    .Y(_0653_),
    .VSS(VGND),
    .A1(_0622_),
    .A2(_0652_));
 sg13g2_nor2_1 _6099_ (.A(net1353),
    .B(_0625_),
    .Y(_0654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6100_ (.Y(_0058_),
    .B1(net437),
    .B2(_0654_),
    .A2(_2792_),
    .A1(net1353),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6101_ (.A(net1261),
    .B(\s0.data_out[18][6] ),
    .X(_0655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6102_ (.B1(net1274),
    .VDD(VPWR),
    .Y(_0656_),
    .VSS(VGND),
    .A1(_0603_),
    .A2(_0655_));
 sg13g2_nand3b_1 _6103_ (.B(_0656_),
    .C(net1470),
    .Y(_0657_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0606_));
 sg13g2_o21ai_1 _6104_ (.B1(_0657_),
    .VDD(VPWR),
    .Y(_0658_),
    .VSS(VGND),
    .A1(net1470),
    .A2(net622));
 sg13g2_inv_1 _6105_ (.VDD(VPWR),
    .Y(_0059_),
    .A(net623),
    .VSS(VGND));
 sg13g2_and2_1 _6106_ (.A(net1261),
    .B(net499),
    .X(_0659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6107_ (.B1(net1274),
    .VDD(VPWR),
    .Y(_0660_),
    .VSS(VGND),
    .A1(_0596_),
    .A2(_0659_));
 sg13g2_nor2_1 _6108_ (.A(net1356),
    .B(_0599_),
    .Y(_0661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6109_ (.Y(_0060_),
    .B1(_0660_),
    .B2(_0661_),
    .A2(_2791_),
    .A1(net1356),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6110_ (.B1(net1262),
    .VDD(VPWR),
    .Y(_0662_),
    .VSS(VGND),
    .A1(net1394),
    .A2(net1249));
 sg13g2_nand2_1 _6111_ (.Y(_0663_),
    .A(net1337),
    .B(net1258),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6112_ (.Y(_0664_),
    .B(_0663_),
    .A_N(_0662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6113_ (.B1(_0664_),
    .VDD(VPWR),
    .Y(_0665_),
    .VSS(VGND),
    .A1(net1262),
    .A2(_0554_));
 sg13g2_nor2_1 _6114_ (.A(net383),
    .B(net1258),
    .Y(_0666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _6115_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0667_),
    .B(_0666_),
    .A(_0664_));
 sg13g2_nor2_1 _6116_ (.A(net1249),
    .B(_0662_),
    .Y(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6117_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2737_),
    .A2(_2756_),
    .Y(_0669_),
    .B1(net1262));
 sg13g2_nor2_1 _6118_ (.A(_0668_),
    .B(_0669_),
    .Y(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6119_ (.B1(net1470),
    .VDD(VPWR),
    .Y(_0671_),
    .VSS(VGND),
    .A1(net543),
    .A2(_0665_));
 sg13g2_a21oi_1 _6120_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0667_),
    .A2(_0670_),
    .Y(_0061_),
    .B1(_0671_));
 sg13g2_nor2_1 _6121_ (.A(net1356),
    .B(_0665_),
    .Y(_0062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6122_ (.A(net1478),
    .B(net322),
    .X(_0063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6123_ (.Y(_0672_),
    .A(net1260),
    .B(net511),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6124_ (.A0(\s0.data_out[18][2] ),
    .A1(\s0.data_out[17][2] ),
    .S(net1259),
    .X(_0673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6125_ (.A(net1252),
    .B_N(net1165),
    .Y(_0674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6126_ (.A2(_0673_),
    .A1(net1252),
    .B1(_0674_),
    .X(_0675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6127_ (.Y(_0676_),
    .B(\s0.data_out[17][2] ),
    .A_N(net1271),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6128_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0562_),
    .A2(_0676_),
    .Y(_0677_),
    .B1(net1268));
 sg13g2_a21oi_1 _6129_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1268),
    .A2(_0675_),
    .Y(_0678_),
    .B1(_0677_));
 sg13g2_nor2_1 _6130_ (.A(net1447),
    .B(_0678_),
    .Y(_0679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6131_ (.Y(_0680_),
    .A(net1260),
    .B(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6132_ (.A0(\s0.data_out[18][1] ),
    .A1(\s0.data_out[17][1] ),
    .S(net1259),
    .X(_0681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6133_ (.A(net1253),
    .B_N(net1169),
    .Y(_0682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6134_ (.A2(_0681_),
    .A1(net1253),
    .B1(_0682_),
    .X(_0683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6135_ (.Y(_0684_),
    .B(\s0.data_out[17][1] ),
    .A_N(net1271),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6136_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0570_),
    .A2(_0684_),
    .Y(_0685_),
    .B1(net1267));
 sg13g2_a21oi_1 _6137_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1267),
    .A2(_0683_),
    .Y(_0686_),
    .B1(_0685_));
 sg13g2_mux2_1 _6138_ (.A0(\s0.data_out[18][0] ),
    .A1(\s0.data_out[17][0] ),
    .S(net1259),
    .X(_0687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6139_ (.A(net1252),
    .B_N(net1172),
    .Y(_0688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6140_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1252),
    .A2(_0687_),
    .Y(_0689_),
    .B1(_0688_));
 sg13g2_nand2b_1 _6141_ (.Y(_0690_),
    .B(net1267),
    .A_N(_0689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6142_ (.A0(\s0.data_out[17][0] ),
    .A1(\s0.data_out[18][0] ),
    .S(net1270),
    .X(_0691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6143_ (.Y(_0692_),
    .B(_0691_),
    .A_N(net1267),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6144_ (.A(net1452),
    .B(_0686_),
    .Y(_0693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _6145_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0692_),
    .C1(net1460),
    .B1(_0690_),
    .A1(net1452),
    .Y(_0694_),
    .A2(_0686_));
 sg13g2_nor3_1 _6146_ (.A(_0679_),
    .B(_0693_),
    .C(_0694_),
    .Y(_0695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6147_ (.Y(_0696_),
    .A(net1259),
    .B(net689),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6148_ (.A0(\s0.data_out[18][3] ),
    .A1(\s0.data_out[17][3] ),
    .S(net1259),
    .X(_0697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6149_ (.A(net1253),
    .B_N(\s0.data_new_delayed[3] ),
    .Y(_0698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6150_ (.A2(_0697_),
    .A1(net1253),
    .B1(_0698_),
    .X(_0699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6151_ (.Y(_0700_),
    .B(\s0.data_out[17][3] ),
    .A_N(net1270),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6152_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0585_),
    .A2(_0700_),
    .Y(_0701_),
    .B1(net1267));
 sg13g2_a21oi_1 _6153_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1267),
    .A2(_0699_),
    .Y(_0702_),
    .B1(_0701_));
 sg13g2_a221oi_1 _6154_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net1439),
    .C1(_0695_),
    .B1(_0702_),
    .A1(net1447),
    .Y(_0703_),
    .A2(_0678_));
 sg13g2_nand2_1 _6155_ (.Y(_0704_),
    .A(net1257),
    .B(net560),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6156_ (.A0(\s0.data_out[18][7] ),
    .A1(\s0.data_out[17][7] ),
    .S(net1258),
    .X(_0705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6157_ (.A(net1249),
    .B_N(net1143),
    .Y(_0706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6158_ (.A2(_0705_),
    .A1(net1249),
    .B1(_0706_),
    .X(_0707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6159_ (.Y(_0708_),
    .B(\s0.data_out[17][7] ),
    .A_N(net1269),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6160_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0594_),
    .A2(_0708_),
    .Y(_0709_),
    .B1(net1262));
 sg13g2_a21oi_1 _6161_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1262),
    .A2(_0707_),
    .Y(_0710_),
    .B1(_0709_));
 sg13g2_nand2_1 _6162_ (.Y(_0711_),
    .A(net1257),
    .B(net664),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6163_ (.A0(\s0.data_out[18][6] ),
    .A1(\s0.data_out[17][6] ),
    .S(net1258),
    .X(_0712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6164_ (.A(net1249),
    .B_N(net1148),
    .Y(_0713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6165_ (.A2(_0712_),
    .A1(net1249),
    .B1(_0713_),
    .X(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6166_ (.Y(_0715_),
    .B(\s0.data_out[17][6] ),
    .A_N(net1269),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6167_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0601_),
    .A2(_0715_),
    .Y(_0716_),
    .B1(net1262));
 sg13g2_a21oi_1 _6168_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1262),
    .A2(_0714_),
    .Y(_0717_),
    .B1(_0716_));
 sg13g2_a22oi_1 _6169_ (.Y(_0718_),
    .B1(_0717_),
    .B2(net1411),
    .A2(_0710_),
    .A1(net1402),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6170_ (.A(net1411),
    .B(_0717_),
    .Y(_0719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _6171_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0720_),
    .B(_0710_),
    .A(net1402));
 sg13g2_nand3b_1 _6172_ (.B(_0720_),
    .C(_0718_),
    .Y(_0721_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0719_));
 sg13g2_nand2_1 _6173_ (.Y(_0722_),
    .A(net1257),
    .B(\s0.data_out[17][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6174_ (.A0(\s0.data_out[18][4] ),
    .A1(\s0.data_out[17][4] ),
    .S(net1259),
    .X(_0723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6175_ (.A(net1252),
    .B_N(net1158),
    .Y(_0724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6176_ (.A2(_0723_),
    .A1(net1252),
    .B1(_0724_),
    .X(_0725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6177_ (.Y(_0726_),
    .B(\s0.data_out[17][4] ),
    .A_N(net1271),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6178_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0613_),
    .A2(_0726_),
    .Y(_0727_),
    .B1(net1268));
 sg13g2_a21oi_1 _6179_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1268),
    .A2(_0725_),
    .Y(_0728_),
    .B1(_0727_));
 sg13g2_nand2_1 _6180_ (.Y(_0729_),
    .A(net1257),
    .B(net368),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6181_ (.A0(\s0.data_out[18][5] ),
    .A1(\s0.data_out[17][5] ),
    .S(net1258),
    .X(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6182_ (.A(net1249),
    .B_N(net1153),
    .Y(_0731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6183_ (.A2(_0730_),
    .A1(net1251),
    .B1(_0731_),
    .X(_0732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6184_ (.Y(_0733_),
    .B(net368),
    .A_N(net1269),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6185_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0620_),
    .A2(_0733_),
    .Y(_0734_),
    .B1(net1263));
 sg13g2_a21oi_1 _6186_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1263),
    .A2(_0732_),
    .Y(_0735_),
    .B1(_0734_));
 sg13g2_a22oi_1 _6187_ (.Y(_0736_),
    .B1(_0735_),
    .B2(net1421),
    .A2(_0728_),
    .A1(net1430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6188_ (.A(net1430),
    .B(_0728_),
    .Y(_0737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6189_ (.A(net1421),
    .B(_0735_),
    .Y(_0738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6190_ (.A(net1439),
    .B(_0702_),
    .Y(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _6191_ (.A(_0737_),
    .B(_0738_),
    .C(_0739_),
    .Y(_0740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6192_ (.Y(_0741_),
    .A(_0736_),
    .B(_0740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _6193_ (.A(_0703_),
    .B(_0721_),
    .C(_0741_),
    .X(_0742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _6194_ (.A(_0721_),
    .B(_0736_),
    .C(_0738_),
    .Y(_0743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6195_ (.A(_0718_),
    .B_N(_0720_),
    .Y(_0744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _6196_ (.A(_0665_),
    .B(_0743_),
    .C(_0744_),
    .Y(_0745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _6197_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0746_),
    .B(net1330),
    .A(net337));
 sg13g2_a21oi_1 _6198_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0742_),
    .A2(_0745_),
    .Y(_0064_),
    .B1(_0746_));
 sg13g2_and2_1 _6199_ (.A(net1252),
    .B(\s0.data_out[17][0] ),
    .X(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6200_ (.B1(net1267),
    .VDD(VPWR),
    .Y(_0748_),
    .VSS(VGND),
    .A1(_0688_),
    .A2(_0747_));
 sg13g2_nand3_1 _6201_ (.B(_0692_),
    .C(_0748_),
    .A(net1471),
    .Y(_0749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6202_ (.B1(_0749_),
    .VDD(VPWR),
    .Y(_0750_),
    .VSS(VGND),
    .A1(net1471),
    .A2(net660));
 sg13g2_inv_1 _6203_ (.VDD(VPWR),
    .Y(_0065_),
    .A(_0750_),
    .VSS(VGND));
 sg13g2_nor2_1 _6204_ (.A(net1002),
    .B(_2807_),
    .Y(_0751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6205_ (.B1(net1268),
    .VDD(VPWR),
    .Y(_0752_),
    .VSS(VGND),
    .A1(_0682_),
    .A2(_0751_));
 sg13g2_nor2_1 _6206_ (.A(net1366),
    .B(_0685_),
    .Y(_0753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6207_ (.Y(_0066_),
    .B1(_0752_),
    .B2(_0753_),
    .A2(_2802_),
    .A1(net1366),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6208_ (.A(_2757_),
    .B(_2806_),
    .Y(_0754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6209_ (.B1(net1268),
    .VDD(VPWR),
    .Y(_0755_),
    .VSS(VGND),
    .A1(_0674_),
    .A2(_0754_));
 sg13g2_nor2_1 _6210_ (.A(net1357),
    .B(_0677_),
    .Y(_0756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6211_ (.Y(_0067_),
    .B1(_0755_),
    .B2(_0756_),
    .A2(_2801_),
    .A1(net1355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6212_ (.A(_2757_),
    .B(_2805_),
    .Y(_0757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6213_ (.B1(net1267),
    .VDD(VPWR),
    .Y(_0758_),
    .VSS(VGND),
    .A1(_0698_),
    .A2(_0757_));
 sg13g2_nor2_1 _6214_ (.A(net1357),
    .B(_0701_),
    .Y(_0759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6215_ (.Y(_0068_),
    .B1(_0758_),
    .B2(_0759_),
    .A2(_2800_),
    .A1(net1357),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6216_ (.A(net1252),
    .B(\s0.data_out[17][4] ),
    .X(_0760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6217_ (.B1(net1268),
    .VDD(VPWR),
    .Y(_0761_),
    .VSS(VGND),
    .A1(_0724_),
    .A2(_0760_));
 sg13g2_nor2_1 _6218_ (.A(net1356),
    .B(_0727_),
    .Y(_0762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6219_ (.Y(_0069_),
    .B1(_0761_),
    .B2(_0762_),
    .A2(_2799_),
    .A1(net1356),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6220_ (.A(net1002),
    .B(_2804_),
    .Y(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6221_ (.B1(net1263),
    .VDD(VPWR),
    .Y(_0764_),
    .VSS(VGND),
    .A1(_0731_),
    .A2(_0763_));
 sg13g2_nor2_1 _6222_ (.A(net1356),
    .B(net369),
    .Y(_0765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6223_ (.Y(_0070_),
    .B1(_0764_),
    .B2(_0765_),
    .A2(_2798_),
    .A1(net1356),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6224_ (.A(net1249),
    .B(\s0.data_out[17][6] ),
    .X(_0766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6225_ (.B1(net1262),
    .VDD(VPWR),
    .Y(_0767_),
    .VSS(VGND),
    .A1(_0713_),
    .A2(_0766_));
 sg13g2_nand3b_1 _6226_ (.B(_0767_),
    .C(net1470),
    .Y(_0768_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0716_));
 sg13g2_o21ai_1 _6227_ (.B1(_0768_),
    .VDD(VPWR),
    .Y(_0769_),
    .VSS(VGND),
    .A1(net1470),
    .A2(net534));
 sg13g2_inv_1 _6228_ (.VDD(VPWR),
    .Y(_0071_),
    .A(net535),
    .VSS(VGND));
 sg13g2_nor2_1 _6229_ (.A(net1002),
    .B(_2803_),
    .Y(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6230_ (.B1(net1263),
    .VDD(VPWR),
    .Y(_0771_),
    .VSS(VGND),
    .A1(_0706_),
    .A2(_0770_));
 sg13g2_nor2_1 _6231_ (.A(net1365),
    .B(_0709_),
    .Y(_0772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6232_ (.Y(_0072_),
    .B1(_0771_),
    .B2(_0772_),
    .A2(_2797_),
    .A1(net1365),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6233_ (.B1(net1250),
    .VDD(VPWR),
    .Y(_0773_),
    .VSS(VGND),
    .A1(net1394),
    .A2(net1236));
 sg13g2_a21oi_1 _6234_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1337),
    .A2(net1245),
    .Y(_0774_),
    .B1(_0773_));
 sg13g2_a21oi_1 _6235_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1002),
    .A2(_0663_),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_o21ai_1 _6236_ (.B1(_0774_),
    .VDD(VPWR),
    .Y(_0776_),
    .VSS(VGND),
    .A1(net370),
    .A2(net1245));
 sg13g2_nor2_1 _6237_ (.A(net1236),
    .B(_0773_),
    .Y(_0777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6238_ (.B1(net1002),
    .VDD(VPWR),
    .Y(_0778_),
    .VSS(VGND),
    .A1(net370),
    .A2(net1257));
 sg13g2_nand2_1 _6239_ (.Y(_0779_),
    .A(_0776_),
    .B(_0778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6240_ (.B1(net1478),
    .VDD(VPWR),
    .Y(_0780_),
    .VSS(VGND),
    .A1(_0777_),
    .A2(_0779_));
 sg13g2_a21oi_1 _6241_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2737_),
    .A2(_0775_),
    .Y(_0073_),
    .B1(_0780_));
 sg13g2_and2_1 _6242_ (.A(net1478),
    .B(_0775_),
    .X(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6243_ (.A(net1477),
    .B(net326),
    .X(_0075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6244_ (.Y(_0781_),
    .A(net1248),
    .B(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6245_ (.A0(\s0.data_out[17][2] ),
    .A1(\s0.data_out[16][2] ),
    .S(net1246),
    .X(_0782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6246_ (.A(net1238),
    .B_N(net1165),
    .Y(_0783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6247_ (.A2(_0782_),
    .A1(net1238),
    .B1(_0783_),
    .X(_0784_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6248_ (.Y(_0785_),
    .B(net426),
    .A_N(net1259),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6249_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0672_),
    .A2(_0785_),
    .Y(_0786_),
    .B1(net1254));
 sg13g2_a21oi_1 _6250_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1254),
    .A2(_0784_),
    .Y(_0787_),
    .B1(_0786_));
 sg13g2_or2_1 _6251_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0788_),
    .B(_0787_),
    .A(net1447));
 sg13g2_nor2b_1 _6252_ (.A(net1239),
    .B_N(net1169),
    .Y(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6253_ (.Y(_0790_),
    .A(net1245),
    .B(net479),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6254_ (.B1(_0790_),
    .VDD(VPWR),
    .Y(_0791_),
    .VSS(VGND),
    .A1(net1246),
    .A2(_2807_));
 sg13g2_a21o_1 _6255_ (.A2(_0791_),
    .A1(net1239),
    .B1(_0789_),
    .X(_0792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6256_ (.Y(_0793_),
    .B(net479),
    .A_N(net1260),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6257_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0680_),
    .A2(_0793_),
    .Y(_0794_),
    .B1(net1255));
 sg13g2_a21oi_1 _6258_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1254),
    .A2(_0792_),
    .Y(_0795_),
    .B1(_0794_));
 sg13g2_mux2_1 _6259_ (.A0(\s0.data_out[17][0] ),
    .A1(\s0.data_out[16][0] ),
    .S(net1245),
    .X(_0796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6260_ (.A(net1238),
    .B_N(net1172),
    .Y(_0797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6261_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1238),
    .A2(_0796_),
    .Y(_0798_),
    .B1(_0797_));
 sg13g2_nand2b_1 _6262_ (.Y(_0799_),
    .B(net1255),
    .A_N(_0798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6263_ (.A0(\s0.data_out[16][0] ),
    .A1(\s0.data_out[17][0] ),
    .S(net1260),
    .X(_0800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6264_ (.Y(_0801_),
    .A(_2757_),
    .B(_0800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6265_ (.B1(_0788_),
    .VDD(VPWR),
    .Y(_0802_),
    .VSS(VGND),
    .A1(net1453),
    .A2(_0795_));
 sg13g2_a221oi_1 _6266_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0801_),
    .C1(net1460),
    .B1(_0799_),
    .A1(net1453),
    .Y(_0803_),
    .A2(_0795_));
 sg13g2_nand2_1 _6267_ (.Y(_0804_),
    .A(net1246),
    .B(net482),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6268_ (.B1(_0804_),
    .VDD(VPWR),
    .Y(_0805_),
    .VSS(VGND),
    .A1(net1246),
    .A2(_2805_));
 sg13g2_nor2_1 _6269_ (.A(net1238),
    .B(net994),
    .Y(_0806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6270_ (.A2(_0805_),
    .A1(net1239),
    .B1(_0806_),
    .X(_0807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6271_ (.Y(_0808_),
    .B(net482),
    .A_N(net1259),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6272_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0696_),
    .A2(_0808_),
    .Y(_0809_),
    .B1(net1254));
 sg13g2_a21oi_1 _6273_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1254),
    .A2(_0807_),
    .Y(_0810_),
    .B1(_0809_));
 sg13g2_a22oi_1 _6274_ (.Y(_0811_),
    .B1(_0810_),
    .B2(net1439),
    .A2(_0787_),
    .A1(net1447),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6275_ (.B1(_0811_),
    .VDD(VPWR),
    .Y(_0812_),
    .VSS(VGND),
    .A1(_0802_),
    .A2(_0803_));
 sg13g2_nand2_1 _6276_ (.Y(_0813_),
    .A(net1247),
    .B(net503),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6277_ (.A0(\s0.data_out[17][7] ),
    .A1(\s0.data_out[16][7] ),
    .S(net1245),
    .X(_0814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6278_ (.A(net1236),
    .B_N(net1144),
    .Y(_0815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6279_ (.A2(_0814_),
    .A1(net1236),
    .B1(_0815_),
    .X(_0816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6280_ (.Y(_0817_),
    .B(net503),
    .A_N(net1257),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6281_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0704_),
    .A2(_0817_),
    .Y(_0818_),
    .B1(net1250));
 sg13g2_a21oi_1 _6282_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1250),
    .A2(_0816_),
    .Y(_0819_),
    .B1(_0818_));
 sg13g2_nand2_1 _6283_ (.Y(_0820_),
    .A(net1247),
    .B(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6284_ (.A0(\s0.data_out[17][6] ),
    .A1(\s0.data_out[16][6] ),
    .S(net1245),
    .X(_0821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6285_ (.A(net1237),
    .B_N(net1149),
    .Y(_0822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6286_ (.A2(_0821_),
    .A1(net1237),
    .B1(_0822_),
    .X(_0823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6287_ (.Y(_0824_),
    .B(net599),
    .A_N(net1257),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6288_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0711_),
    .A2(_0824_),
    .Y(_0825_),
    .B1(net1250));
 sg13g2_a21oi_1 _6289_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1250),
    .A2(_0823_),
    .Y(_0826_),
    .B1(_0825_));
 sg13g2_a22oi_1 _6290_ (.Y(_0827_),
    .B1(_0826_),
    .B2(net1411),
    .A2(_0819_),
    .A1(net1402),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _6291_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0828_),
    .B(_0826_),
    .A(net1411));
 sg13g2_or2_1 _6292_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0829_),
    .B(_0819_),
    .A(net1402));
 sg13g2_inv_1 _6293_ (.VDD(VPWR),
    .Y(_0830_),
    .A(_0829_),
    .VSS(VGND));
 sg13g2_and3_1 _6294_ (.X(_0831_),
    .A(_0827_),
    .B(_0828_),
    .C(_0829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _6295_ (.B(_0828_),
    .C(_0829_),
    .A(_0827_),
    .Y(_0832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6296_ (.Y(_0833_),
    .A(net1248),
    .B(net475),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6297_ (.A0(\s0.data_out[17][5] ),
    .A1(\s0.data_out[16][5] ),
    .S(net1245),
    .X(_0834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6298_ (.A(net1236),
    .B_N(net1153),
    .Y(_0835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6299_ (.A2(_0834_),
    .A1(net1236),
    .B1(_0835_),
    .X(_0836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6300_ (.Y(_0837_),
    .B(net475),
    .A_N(net1258),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6301_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0729_),
    .A2(_0837_),
    .Y(_0838_),
    .B1(net1251));
 sg13g2_a21oi_1 _6302_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1251),
    .A2(_0836_),
    .Y(_0839_),
    .B1(_0838_));
 sg13g2_nand2_1 _6303_ (.Y(_0840_),
    .A(net1421),
    .B(_0839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6304_ (.A(net1237),
    .B_N(net1158),
    .Y(_0841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6305_ (.Y(_0842_),
    .A(net1247),
    .B(net525),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6306_ (.A0(\s0.data_out[17][4] ),
    .A1(\s0.data_out[16][4] ),
    .S(net1245),
    .X(_0843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6307_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1237),
    .A2(_0843_),
    .Y(_0844_),
    .B1(_0841_));
 sg13g2_nand2b_1 _6308_ (.Y(_0845_),
    .B(net1250),
    .A_N(_0844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6309_ (.B1(_0722_),
    .VDD(VPWR),
    .Y(_0846_),
    .VSS(VGND),
    .A1(net1257),
    .A2(_2810_));
 sg13g2_nand2_1 _6310_ (.Y(_0847_),
    .A(net1002),
    .B(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _6311_ (.B(_0845_),
    .C(_0847_),
    .A(net1430),
    .Y(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6312_ (.A2(_0847_),
    .A1(_0845_),
    .B1(net1430),
    .X(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6313_ (.A(net1421),
    .B(_0839_),
    .Y(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6314_ (.Y(_0851_),
    .A(_0848_),
    .B(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6315_ (.B1(_0840_),
    .VDD(VPWR),
    .Y(_0852_),
    .VSS(VGND),
    .A1(net1439),
    .A2(_0810_));
 sg13g2_nor4_1 _6316_ (.A(_0832_),
    .B(_0850_),
    .C(_0851_),
    .D(_0852_),
    .Y(_0853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6317_ (.B1(_0840_),
    .VDD(VPWR),
    .Y(_0854_),
    .VSS(VGND),
    .A1(_0848_),
    .A2(_0850_));
 sg13g2_o21ai_1 _6318_ (.B1(_0775_),
    .VDD(VPWR),
    .Y(_0855_),
    .VSS(VGND),
    .A1(_0827_),
    .A2(_0830_));
 sg13g2_a221oi_1 _6319_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0831_),
    .C1(_0855_),
    .B1(_0854_),
    .A1(_0812_),
    .Y(_0856_),
    .A2(_0853_));
 sg13g2_nor3_1 _6320_ (.A(net322),
    .B(net1331),
    .C(_0856_),
    .Y(_0076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6321_ (.A(net1238),
    .B(\s0.data_out[16][0] ),
    .X(_0857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6322_ (.B1(net1255),
    .VDD(VPWR),
    .Y(_0858_),
    .VSS(VGND),
    .A1(_0797_),
    .A2(_0857_));
 sg13g2_nand3_1 _6323_ (.B(_0801_),
    .C(_0858_),
    .A(net1478),
    .Y(_0859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6324_ (.B1(_0859_),
    .VDD(VPWR),
    .Y(_0860_),
    .VSS(VGND),
    .A1(net1478),
    .A2(net653));
 sg13g2_inv_1 _6325_ (.VDD(VPWR),
    .Y(_0077_),
    .A(_0860_),
    .VSS(VGND));
 sg13g2_and2_1 _6326_ (.A(net1238),
    .B(net479),
    .X(_0861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6327_ (.B1(net1255),
    .VDD(VPWR),
    .Y(_0862_),
    .VSS(VGND),
    .A1(_0789_),
    .A2(_0861_));
 sg13g2_nor2_1 _6328_ (.A(net1366),
    .B(_0794_),
    .Y(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6329_ (.Y(_0078_),
    .B1(_0862_),
    .B2(_0863_),
    .A2(_2807_),
    .A1(net1366),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6330_ (.A(net1238),
    .B(net426),
    .X(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6331_ (.B1(net1254),
    .VDD(VPWR),
    .Y(_0865_),
    .VSS(VGND),
    .A1(_0783_),
    .A2(_0864_));
 sg13g2_nor2_1 _6332_ (.A(net1366),
    .B(_0786_),
    .Y(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6333_ (.Y(_0079_),
    .B1(_0865_),
    .B2(_0866_),
    .A2(_2806_),
    .A1(net1366),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6334_ (.A(net1239),
    .B(net482),
    .X(_0867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6335_ (.B1(net1254),
    .VDD(VPWR),
    .Y(_0868_),
    .VSS(VGND),
    .A1(_0806_),
    .A2(_0867_));
 sg13g2_nor2_1 _6336_ (.A(net1365),
    .B(_0809_),
    .Y(_0869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6337_ (.Y(_0080_),
    .B1(_0868_),
    .B2(_0869_),
    .A2(_2805_),
    .A1(net1366),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6338_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1237),
    .A2(net525),
    .Y(_0870_),
    .B1(_0841_));
 sg13g2_a21oi_1 _6339_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1002),
    .A2(_0846_),
    .Y(_0871_),
    .B1(net1365));
 sg13g2_o21ai_1 _6340_ (.B1(_0871_),
    .VDD(VPWR),
    .Y(_0872_),
    .VSS(VGND),
    .A1(net1002),
    .A2(_0870_));
 sg13g2_o21ai_1 _6341_ (.B1(_0872_),
    .VDD(VPWR),
    .Y(_0873_),
    .VSS(VGND),
    .A1(net1478),
    .A2(net668));
 sg13g2_inv_1 _6342_ (.VDD(VPWR),
    .Y(_0081_),
    .A(_0873_),
    .VSS(VGND));
 sg13g2_and2_1 _6343_ (.A(net1236),
    .B(net475),
    .X(_0874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6344_ (.B1(net1251),
    .VDD(VPWR),
    .Y(_0875_),
    .VSS(VGND),
    .A1(_0835_),
    .A2(_0874_));
 sg13g2_nor2_1 _6345_ (.A(net1365),
    .B(_0838_),
    .Y(_0876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6346_ (.Y(_0082_),
    .B1(_0875_),
    .B2(_0876_),
    .A2(_2804_),
    .A1(net1365),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6347_ (.A(net1237),
    .B(\s0.data_out[16][6] ),
    .X(_0877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6348_ (.B1(net1250),
    .VDD(VPWR),
    .Y(_0878_),
    .VSS(VGND),
    .A1(_0822_),
    .A2(_0877_));
 sg13g2_nand3b_1 _6349_ (.B(_0878_),
    .C(net1478),
    .Y(_0879_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0825_));
 sg13g2_o21ai_1 _6350_ (.B1(_0879_),
    .VDD(VPWR),
    .Y(_0880_),
    .VSS(VGND),
    .A1(net1478),
    .A2(net664));
 sg13g2_inv_1 _6351_ (.VDD(VPWR),
    .Y(_0083_),
    .A(net665),
    .VSS(VGND));
 sg13g2_and2_1 _6352_ (.A(net1236),
    .B(net503),
    .X(_0881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6353_ (.B1(net1250),
    .VDD(VPWR),
    .Y(_0882_),
    .VSS(VGND),
    .A1(_0815_),
    .A2(_0881_));
 sg13g2_nor2_1 _6354_ (.A(net1365),
    .B(_0818_),
    .Y(_0883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6355_ (.Y(_0084_),
    .B1(_0882_),
    .B2(_0883_),
    .A2(_2803_),
    .A1(net1365),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6356_ (.B1(net1240),
    .VDD(VPWR),
    .Y(_0884_),
    .VSS(VGND),
    .A1(net1394),
    .A2(net1223));
 sg13g2_a21oi_1 _6357_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1337),
    .A2(net1233),
    .Y(_0885_),
    .B1(_0884_));
 sg13g2_a21oi_1 _6358_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1337),
    .A2(net1247),
    .Y(_0886_),
    .B1(net1240));
 sg13g2_nor2_1 _6359_ (.A(_0885_),
    .B(_0886_),
    .Y(_0887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6360_ (.B1(_0885_),
    .VDD(VPWR),
    .Y(_0888_),
    .VSS(VGND),
    .A1(net362),
    .A2(net1233));
 sg13g2_nor2_1 _6361_ (.A(net1223),
    .B(_0884_),
    .Y(_0889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6362_ (.A(net362),
    .B(net1247),
    .Y(_0890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6363_ (.B1(_0888_),
    .VDD(VPWR),
    .Y(_0891_),
    .VSS(VGND),
    .A1(net1241),
    .A2(_0890_));
 sg13g2_o21ai_1 _6364_ (.B1(net1477),
    .VDD(VPWR),
    .Y(_0892_),
    .VSS(VGND),
    .A1(_0889_),
    .A2(_0891_));
 sg13g2_a21oi_1 _6365_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2736_),
    .A2(_0887_),
    .Y(_0085_),
    .B1(_0892_));
 sg13g2_nor3_1 _6366_ (.A(net1367),
    .B(_0885_),
    .C(_0886_),
    .Y(_0086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6367_ (.A(net1484),
    .B(net323),
    .X(_0087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6368_ (.Y(_0893_),
    .A(net1235),
    .B(net420),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6369_ (.A0(\s0.data_out[16][2] ),
    .A1(\s0.data_out[15][2] ),
    .S(net1232),
    .X(_0894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6370_ (.A(net1225),
    .B_N(net1164),
    .Y(_0895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6371_ (.A2(_0894_),
    .A1(net1225),
    .B1(_0895_),
    .X(_0896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6372_ (.Y(_0897_),
    .B(net420),
    .A_N(net1248),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6373_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0781_),
    .A2(_0897_),
    .Y(_0898_),
    .B1(net1242));
 sg13g2_a21oi_1 _6374_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1242),
    .A2(_0896_),
    .Y(_0899_),
    .B1(_0898_));
 sg13g2_or2_1 _6375_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0900_),
    .B(_0899_),
    .A(net1446));
 sg13g2_nand2_1 _6376_ (.Y(_0901_),
    .A(net1232),
    .B(net530),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6377_ (.B1(_0901_),
    .VDD(VPWR),
    .Y(_0902_),
    .VSS(VGND),
    .A1(net1232),
    .A2(_2813_));
 sg13g2_nor2b_1 _6378_ (.A(net1226),
    .B_N(net1168),
    .Y(_0903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6379_ (.A2(_0902_),
    .A1(net1226),
    .B1(_0903_),
    .X(_0904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6380_ (.Y(_0905_),
    .B(\s0.data_out[15][1] ),
    .A_N(net1248),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6381_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0790_),
    .A2(_0905_),
    .Y(_0906_),
    .B1(net1239));
 sg13g2_a21oi_1 _6382_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1242),
    .A2(_0904_),
    .Y(_0907_),
    .B1(_0906_));
 sg13g2_mux2_1 _6383_ (.A0(\s0.data_out[16][0] ),
    .A1(\s0.data_out[15][0] ),
    .S(net1232),
    .X(_0908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6384_ (.A(net1226),
    .B_N(net1171),
    .Y(_0909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6385_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1225),
    .A2(_0908_),
    .Y(_0910_),
    .B1(_0909_));
 sg13g2_nand2b_1 _6386_ (.Y(_0911_),
    .B(net1243),
    .A_N(_0910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6387_ (.A0(\s0.data_out[15][0] ),
    .A1(\s0.data_out[16][0] ),
    .S(net1248),
    .X(_0912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6388_ (.Y(_0913_),
    .B(_0912_),
    .A_N(net1243),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _6389_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0913_),
    .C1(net1459),
    .B1(_0911_),
    .A1(net1456),
    .Y(_0914_),
    .A2(_0907_));
 sg13g2_o21ai_1 _6390_ (.B1(_0900_),
    .VDD(VPWR),
    .Y(_0915_),
    .VSS(VGND),
    .A1(net1456),
    .A2(_0907_));
 sg13g2_nand2_1 _6391_ (.Y(_0916_),
    .A(net1232),
    .B(net553),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6392_ (.B1(_0916_),
    .VDD(VPWR),
    .Y(_0917_),
    .VSS(VGND),
    .A1(net1232),
    .A2(_2811_));
 sg13g2_nor2_1 _6393_ (.A(net1226),
    .B(net994),
    .Y(_0918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6394_ (.A2(_0917_),
    .A1(net1225),
    .B1(_0918_),
    .X(_0919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6395_ (.Y(_0920_),
    .B(\s0.data_out[15][3] ),
    .A_N(net1248),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6396_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0804_),
    .A2(_0920_),
    .Y(_0921_),
    .B1(net1242));
 sg13g2_a21oi_1 _6397_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1242),
    .A2(_0919_),
    .Y(_0922_),
    .B1(_0921_));
 sg13g2_a22oi_1 _6398_ (.Y(_0923_),
    .B1(_0922_),
    .B2(net1440),
    .A2(_0899_),
    .A1(net1446),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6399_ (.B1(_0923_),
    .VDD(VPWR),
    .Y(_0924_),
    .VSS(VGND),
    .A1(_0914_),
    .A2(_0915_));
 sg13g2_nand2_1 _6400_ (.Y(_0925_),
    .A(net1234),
    .B(\s0.data_out[15][6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6401_ (.A0(\s0.data_out[16][6] ),
    .A1(\s0.data_out[15][6] ),
    .S(net1233),
    .X(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6402_ (.A(net1223),
    .B_N(net1149),
    .Y(_0927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6403_ (.A2(_0926_),
    .A1(net1223),
    .B1(_0927_),
    .X(_0928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6404_ (.Y(_0929_),
    .B(\s0.data_out[15][6] ),
    .A_N(net1247),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6405_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0820_),
    .A2(_0929_),
    .Y(_0930_),
    .B1(net1240));
 sg13g2_a21oi_1 _6406_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1240),
    .A2(_0928_),
    .Y(_0931_),
    .B1(_0930_));
 sg13g2_nand2_1 _6407_ (.Y(_0932_),
    .A(net1234),
    .B(net561),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6408_ (.A0(\s0.data_out[16][7] ),
    .A1(\s0.data_out[15][7] ),
    .S(net1233),
    .X(_0933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6409_ (.A(net1224),
    .B_N(net1144),
    .Y(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6410_ (.A2(_0933_),
    .A1(net1224),
    .B1(_0934_),
    .X(_0935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6411_ (.Y(_0936_),
    .B(\s0.data_out[15][7] ),
    .A_N(net1247),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6412_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0813_),
    .A2(_0936_),
    .Y(_0937_),
    .B1(net1241));
 sg13g2_a21oi_1 _6413_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1241),
    .A2(_0935_),
    .Y(_0938_),
    .B1(_0937_));
 sg13g2_a22oi_1 _6414_ (.Y(_0939_),
    .B1(_0938_),
    .B2(net1402),
    .A2(_0931_),
    .A1(net1411),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _6415_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0940_),
    .B(_0931_),
    .A(net1411));
 sg13g2_or2_1 _6416_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0941_),
    .B(_0938_),
    .A(net1402));
 sg13g2_inv_1 _6417_ (.VDD(VPWR),
    .Y(_0942_),
    .A(_0941_),
    .VSS(VGND));
 sg13g2_and3_1 _6418_ (.X(_0943_),
    .A(_0939_),
    .B(_0940_),
    .C(_0941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _6419_ (.B(_0940_),
    .C(_0941_),
    .A(_0939_),
    .Y(_0944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6420_ (.Y(_0945_),
    .A(net1233),
    .B(\s0.data_out[15][4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6421_ (.B1(_0945_),
    .VDD(VPWR),
    .Y(_0946_),
    .VSS(VGND),
    .A1(net1233),
    .A2(_2810_));
 sg13g2_nor2b_1 _6422_ (.A(net1223),
    .B_N(net1158),
    .Y(_0947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6423_ (.A2(_0946_),
    .A1(net1223),
    .B1(_0947_),
    .X(_0948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6424_ (.Y(_0949_),
    .B(\s0.data_out[15][4] ),
    .A_N(net1247),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6425_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0842_),
    .A2(_0949_),
    .Y(_0950_),
    .B1(net1240));
 sg13g2_a21oi_1 _6426_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1240),
    .A2(_0948_),
    .Y(_0951_),
    .B1(_0950_));
 sg13g2_nand2_1 _6427_ (.Y(_0952_),
    .A(net1430),
    .B(_0951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6428_ (.Y(_0953_),
    .A(net1234),
    .B(net430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _6429_ (.A0(\s0.data_out[16][5] ),
    .A1(\s0.data_out[15][5] ),
    .S(net1233),
    .X(_0954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _6430_ (.A(net1224),
    .B_N(net1154),
    .Y(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _6431_ (.A2(_0954_),
    .A1(net1224),
    .B1(_0955_),
    .X(_0956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _6432_ (.Y(_0957_),
    .B(net430),
    .A_N(net1248),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6433_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0833_),
    .A2(_0957_),
    .Y(_0958_),
    .B1(net1241));
 sg13g2_a21oi_1 _6434_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1241),
    .A2(_0956_),
    .Y(_0959_),
    .B1(_0958_));
 sg13g2_nor2_1 _6435_ (.A(net1421),
    .B(_0959_),
    .Y(_0960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _6436_ (.Y(_0961_),
    .A(net1421),
    .B(_0959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6437_ (.B1(_0961_),
    .VDD(VPWR),
    .Y(_0962_),
    .VSS(VGND),
    .A1(net1440),
    .A2(_0922_));
 sg13g2_xnor2_1 _6438_ (.Y(_0963_),
    .A(net1430),
    .B(_0951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _6439_ (.A(_0944_),
    .B(_0960_),
    .C(_0962_),
    .D(_0963_),
    .Y(_0964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6440_ (.B1(_0961_),
    .VDD(VPWR),
    .Y(_0965_),
    .VSS(VGND),
    .A1(_0952_),
    .A2(_0960_));
 sg13g2_o21ai_1 _6441_ (.B1(_0887_),
    .VDD(VPWR),
    .Y(_0966_),
    .VSS(VGND),
    .A1(_0939_),
    .A2(_0942_));
 sg13g2_a221oi_1 _6442_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0943_),
    .C1(_0966_),
    .B1(_0965_),
    .A1(_0924_),
    .Y(_0967_),
    .A2(_0964_));
 sg13g2_nor3_1 _6443_ (.A(net326),
    .B(net1331),
    .C(_0967_),
    .Y(_0088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6444_ (.A(net1226),
    .B(\s0.data_out[15][0] ),
    .X(_0968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6445_ (.B1(net1243),
    .VDD(VPWR),
    .Y(_0969_),
    .VSS(VGND),
    .A1(_0909_),
    .A2(_0968_));
 sg13g2_nand3_1 _6446_ (.B(_0913_),
    .C(_0969_),
    .A(net1477),
    .Y(_0970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6447_ (.B1(_0970_),
    .VDD(VPWR),
    .Y(_0971_),
    .VSS(VGND),
    .A1(net1483),
    .A2(net662));
 sg13g2_inv_1 _6448_ (.VDD(VPWR),
    .Y(_0089_),
    .A(_0971_),
    .VSS(VGND));
 sg13g2_and2_1 _6449_ (.A(net1225),
    .B(\s0.data_out[15][1] ),
    .X(_0972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6450_ (.B1(net1242),
    .VDD(VPWR),
    .Y(_0973_),
    .VSS(VGND),
    .A1(_0903_),
    .A2(_0972_));
 sg13g2_nor2_1 _6451_ (.A(net1369),
    .B(_0906_),
    .Y(_0974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6452_ (.Y(_0090_),
    .B1(_0973_),
    .B2(_0974_),
    .A2(_2813_),
    .A1(net1369),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6453_ (.A(net1225),
    .B(net420),
    .X(_0975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6454_ (.B1(net1242),
    .VDD(VPWR),
    .Y(_0976_),
    .VSS(VGND),
    .A1(_0895_),
    .A2(_0975_));
 sg13g2_nor2_1 _6455_ (.A(net1367),
    .B(_0898_),
    .Y(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6456_ (.Y(_0091_),
    .B1(_0976_),
    .B2(_0977_),
    .A2(_2812_),
    .A1(net1367),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6457_ (.A(net1225),
    .B(\s0.data_out[15][3] ),
    .X(_0978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6458_ (.B1(net1242),
    .VDD(VPWR),
    .Y(_0979_),
    .VSS(VGND),
    .A1(_0918_),
    .A2(_0978_));
 sg13g2_nor2_1 _6459_ (.A(net1369),
    .B(_0921_),
    .Y(_0980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6460_ (.Y(_0092_),
    .B1(_0979_),
    .B2(_0980_),
    .A2(_2811_),
    .A1(net1369),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6461_ (.A(net1223),
    .B(\s0.data_out[15][4] ),
    .X(_0981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6462_ (.B1(net1240),
    .VDD(VPWR),
    .Y(_0982_),
    .VSS(VGND),
    .A1(_0947_),
    .A2(_0981_));
 sg13g2_nor2_1 _6463_ (.A(net1367),
    .B(_0950_),
    .Y(_0983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6464_ (.Y(_0093_),
    .B1(_0982_),
    .B2(_0983_),
    .A2(_2810_),
    .A1(net1367),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6465_ (.A(net1224),
    .B(net430),
    .X(_0984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6466_ (.B1(net1241),
    .VDD(VPWR),
    .Y(_0985_),
    .VSS(VGND),
    .A1(_0955_),
    .A2(_0984_));
 sg13g2_nor2_1 _6467_ (.A(net1368),
    .B(_0958_),
    .Y(_0986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6468_ (.Y(_0094_),
    .B1(_0985_),
    .B2(_0986_),
    .A2(_2809_),
    .A1(net1368),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _6469_ (.A(net1223),
    .B(\s0.data_out[15][6] ),
    .X(_0987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6470_ (.B1(net1240),
    .VDD(VPWR),
    .Y(_0988_),
    .VSS(VGND),
    .A1(_0927_),
    .A2(_0987_));
 sg13g2_nand3b_1 _6471_ (.B(_0988_),
    .C(net1477),
    .Y(_0989_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0930_));
 sg13g2_o21ai_1 _6472_ (.B1(_0989_),
    .VDD(VPWR),
    .Y(_0990_),
    .VSS(VGND),
    .A1(net1477),
    .A2(net599));
 sg13g2_inv_1 _6473_ (.VDD(VPWR),
    .Y(_0095_),
    .A(_0990_),
    .VSS(VGND));
 sg13g2_and2_1 _6474_ (.A(net1224),
    .B(\s0.data_out[15][7] ),
    .X(_0991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6475_ (.B1(net1241),
    .VDD(VPWR),
    .Y(_0992_),
    .VSS(VGND),
    .A1(_0934_),
    .A2(_0991_));
 sg13g2_nor2_1 _6476_ (.A(net1368),
    .B(_0937_),
    .Y(_0993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _6477_ (.Y(_0096_),
    .B1(_0992_),
    .B2(_0993_),
    .A2(_2808_),
    .A1(net1368),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6478_ (.B1(net1229),
    .VDD(VPWR),
    .Y(_0994_),
    .VSS(VGND),
    .A1(net1217),
    .A2(net1395));
 sg13g2_nor2b_1 _6479_ (.A(net1395),
    .B_N(net1221),
    .Y(_0995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6480_ (.A(_0994_),
    .B(_0995_),
    .Y(_0996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _6481_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1337),
    .A2(net1235),
    .Y(_0997_),
    .B1(net1229));
 sg13g2_nor2_1 _6482_ (.A(_0996_),
    .B(_0997_),
    .Y(_0998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6483_ (.B1(_0996_),
    .VDD(VPWR),
    .Y(_0999_),
    .VSS(VGND),
    .A1(\s0.was_valid_out[14] [0]),
    .A2(net1221));
 sg13g2_nor2_1 _6484_ (.A(net1217),
    .B(_0994_),
    .Y(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _6485_ (.A(\s0.was_valid_out[14] [0]),
    .B(net1234),
    .Y(_1001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _6486_ (.B1(_0999_),
    .VDD(VPWR),
    .Y(_1002_),
    .VSS(VGND),
    .A1(net1229),
    .A2(_1001_));
 sg13g2_o21ai_1 _6487_ (.B1(net1484),
    .VDD(VPWR),
    .Y(_1003_),
    .VSS(VGND),
    .A1(_1000_),
    .A2(_1002_));
 sg13g2_a21oi_1 _6488_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2735_),
    .A2(_0998_),
    .Y(_0097_),
    .B1(_1003_));
 sg13g2_nor3_1 _6489_ (.A(net1380),
    .B(_0996_),
    .C(_0997_),
    .Y(_0098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _6490_ (.RESET_B(net215),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0000_),
    .Q(\s0.module0.bubble ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6491_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0001_),
    .Q(\s0.was_valid_out[23] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6492_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0002_),
    .Q(\s0.valid_out[23] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6493_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0003_),
    .Q(\s0.genblk1[22].modules.bubble ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _6494_ (.RESET_B(net59),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0004_),
    .Q(\s0.shift_out[23] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6495_ (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net380),
    .Q(\s0.data_out[23][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6496_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net382),
    .Q(\s0.data_out[23][1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6497_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net413),
    .Q(\s0.data_out[23][2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6498_ (.RESET_B(net55),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0008_),
    .Q(\s0.data_out[23][3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6499_ (.RESET_B(net54),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net417),
    .Q(\s0.data_out[23][4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6500_ (.RESET_B(net53),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net460),
    .Q(\s0.data_out[23][5] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6501_ (.RESET_B(net52),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net456),
    .Q(\s0.data_out[23][6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6502_ (.RESET_B(net51),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net439),
    .Q(\s0.data_out[23][7] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6503_ (.RESET_B(net50),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net393),
    .Q(\s0.was_valid_out[22] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6504_ (.RESET_B(net48),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0014_),
    .Q(\s0.valid_out[22] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6505_ (.RESET_B(net47),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0015_),
    .Q(\s0.genblk1[21].modules.bubble ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6506_ (.RESET_B(net46),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0016_),
    .Q(\s0.shift_out[22] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6507_ (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net604),
    .Q(\s0.data_out[22][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6508_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net641),
    .Q(\s0.data_out[22][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6509_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0019_),
    .Q(\s0.data_out[22][2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6510_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net587),
    .Q(\s0.data_out[22][3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6511_ (.RESET_B(net41),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0021_),
    .Q(\s0.data_out[22][4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _6512_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0022_),
    .Q(\s0.data_out[22][5] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _6513_ (.RESET_B(net39),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net594),
    .Q(\s0.data_out[22][6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _6514_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0024_),
    .Q(\s0.data_out[22][7] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6515_ (.RESET_B(net37),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0025_),
    .Q(\s0.was_valid_out[21] [0]),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6516_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0026_),
    .Q(\s0.valid_out[21] [0]),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6517_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0027_),
    .Q(\s0.genblk1[20].modules.bubble ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6518_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0028_),
    .Q(\s0.shift_out[21] [0]),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6519_ (.RESET_B(net32),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0029_),
    .Q(\s0.data_out[21][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6520_ (.RESET_B(net31),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net558),
    .Q(\s0.data_out[21][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6521_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0031_),
    .Q(\s0.data_out[21][2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6522_ (.RESET_B(net29),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net520),
    .Q(\s0.data_out[21][3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6523_ (.RESET_B(net28),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0033_),
    .Q(\s0.data_out[21][4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6524_ (.RESET_B(net27),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0034_),
    .Q(\s0.data_out[21][5] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6525_ (.RESET_B(net26),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0035_),
    .Q(\s0.data_out[21][6] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6526_ (.RESET_B(net25),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0036_),
    .Q(\s0.data_out[21][7] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6527_ (.RESET_B(net24),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0037_),
    .Q(\s0.was_valid_out[20] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6528_ (.RESET_B(net318),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0038_),
    .Q(\s0.valid_out[20] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6529_ (.RESET_B(net317),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0039_),
    .Q(\s0.genblk1[1].modules.bubble ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6530_ (.RESET_B(net316),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0040_),
    .Q(\s0.shift_out[20] [0]),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6531_ (.RESET_B(net315),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0041_),
    .Q(\s0.data_out[20][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6532_ (.RESET_B(net314),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net634),
    .Q(\s0.data_out[20][1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6533_ (.RESET_B(net313),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net425),
    .Q(\s0.data_out[20][2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6534_ (.RESET_B(net312),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net629),
    .Q(\s0.data_out[20][3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6535_ (.RESET_B(net311),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net497),
    .Q(\s0.data_out[20][4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6536_ (.RESET_B(net310),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net469),
    .Q(\s0.data_out[20][5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6537_ (.RESET_B(net309),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net433),
    .Q(\s0.data_out[20][6] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6538_ (.RESET_B(net308),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net474),
    .Q(\s0.data_out[20][7] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6539_ (.RESET_B(net307),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net367),
    .Q(\s0.was_valid_out[19] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6540_ (.RESET_B(net305),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0050_),
    .Q(\s0.valid_out[19] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6541_ (.RESET_B(net304),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0051_),
    .Q(\s0.genblk1[18].modules.bubble ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6542_ (.RESET_B(net303),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0052_),
    .Q(\s0.shift_out[19] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6543_ (.RESET_B(net302),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0053_),
    .Q(\s0.data_out[19][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6544_ (.RESET_B(net301),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net696),
    .Q(\s0.data_out[19][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6545_ (.RESET_B(net300),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net658),
    .Q(\s0.data_out[19][2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6546_ (.RESET_B(net299),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net691),
    .Q(\s0.data_out[19][3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6547_ (.RESET_B(net298),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net487),
    .Q(\s0.data_out[19][4] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6548_ (.RESET_B(net297),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0058_),
    .Q(\s0.data_out[19][5] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6549_ (.RESET_B(net296),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0059_),
    .Q(\s0.data_out[19][6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6550_ (.RESET_B(net295),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0060_),
    .Q(\s0.data_out[19][7] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6551_ (.RESET_B(net294),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net544),
    .Q(\s0.was_valid_out[18] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6552_ (.RESET_B(net292),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0062_),
    .Q(\s0.valid_out[18] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6553_ (.RESET_B(net291),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0063_),
    .Q(\s0.genblk1[17].modules.bubble ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6554_ (.RESET_B(net290),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0064_),
    .Q(\s0.shift_out[18] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6555_ (.RESET_B(net289),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0065_),
    .Q(\s0.data_out[18][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6556_ (.RESET_B(net288),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net419),
    .Q(\s0.data_out[18][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6557_ (.RESET_B(net287),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net429),
    .Q(\s0.data_out[18][2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6558_ (.RESET_B(net286),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net411),
    .Q(\s0.data_out[18][3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6559_ (.RESET_B(net285),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net441),
    .Q(\s0.data_out[18][4] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6560_ (.RESET_B(net284),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0070_),
    .Q(\s0.data_out[18][5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6561_ (.RESET_B(net283),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0071_),
    .Q(\s0.data_out[18][6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6562_ (.RESET_B(net282),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net500),
    .Q(\s0.data_out[18][7] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6563_ (.RESET_B(net281),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0073_),
    .Q(\s0.was_valid_out[17] [0]),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6564_ (.RESET_B(net279),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0074_),
    .Q(\s0.valid_out[17] [0]),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6565_ (.RESET_B(net278),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0075_),
    .Q(\s0.genblk1[16].modules.bubble ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6566_ (.RESET_B(net277),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0076_),
    .Q(\s0.shift_out[17] [0]),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6567_ (.RESET_B(net276),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0077_),
    .Q(\s0.data_out[17][0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6568_ (.RESET_B(net275),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0078_),
    .Q(\s0.data_out[17][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6569_ (.RESET_B(net274),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0079_),
    .Q(\s0.data_out[17][2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6570_ (.RESET_B(net273),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0080_),
    .Q(\s0.data_out[17][3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6571_ (.RESET_B(net272),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0081_),
    .Q(\s0.data_out[17][4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6572_ (.RESET_B(net271),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\s0.data_out[17][5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6573_ (.RESET_B(net270),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0083_),
    .Q(\s0.data_out[17][6] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6574_ (.RESET_B(net269),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0084_),
    .Q(\s0.data_out[17][7] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6575_ (.RESET_B(net268),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0085_),
    .Q(\s0.was_valid_out[16] [0]),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6576_ (.RESET_B(net266),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0086_),
    .Q(\s0.valid_out[16] [0]),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6577_ (.RESET_B(net265),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0087_),
    .Q(\s0.genblk1[15].modules.bubble ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6578_ (.RESET_B(net264),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0088_),
    .Q(\s0.shift_out[16] [0]),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6579_ (.RESET_B(net263),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0089_),
    .Q(\s0.data_out[16][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6580_ (.RESET_B(net262),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net480),
    .Q(\s0.data_out[16][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6581_ (.RESET_B(net261),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0091_),
    .Q(\s0.data_out[16][2] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6582_ (.RESET_B(net260),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net483),
    .Q(\s0.data_out[16][3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6583_ (.RESET_B(net259),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net526),
    .Q(\s0.data_out[16][4] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6584_ (.RESET_B(net258),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net476),
    .Q(\s0.data_out[16][5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6585_ (.RESET_B(net257),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0095_),
    .Q(\s0.data_out[16][6] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6586_ (.RESET_B(net256),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net504),
    .Q(\s0.data_out[16][7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6587_ (.RESET_B(net255),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net363),
    .Q(\s0.was_valid_out[15] [0]),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6588_ (.RESET_B(net253),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0098_),
    .Q(\s0.valid_out[15] [0]),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6589_ (.RESET_B(net252),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0099_),
    .Q(\s0.genblk1[14].modules.bubble ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6590_ (.RESET_B(net251),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0100_),
    .Q(\s0.shift_out[15] [0]),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6591_ (.RESET_B(net250),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0101_),
    .Q(\s0.data_out[15][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6592_ (.RESET_B(net249),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net531),
    .Q(\s0.data_out[15][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6593_ (.RESET_B(net248),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net421),
    .Q(\s0.data_out[15][2] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6594_ (.RESET_B(net247),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net554),
    .Q(\s0.data_out[15][3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6595_ (.RESET_B(net246),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0105_),
    .Q(\s0.data_out[15][4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6596_ (.RESET_B(net245),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net431),
    .Q(\s0.data_out[15][5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6597_ (.RESET_B(net244),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0107_),
    .Q(\s0.data_out[15][6] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6598_ (.RESET_B(net243),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net562),
    .Q(\s0.data_out[15][7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6599_ (.RESET_B(net242),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0109_),
    .Q(\s0.was_valid_out[14] [0]),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6600_ (.RESET_B(net240),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0110_),
    .Q(\s0.valid_out[14] [0]),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6601_ (.RESET_B(net239),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0111_),
    .Q(\s0.genblk1[13].modules.bubble ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6602_ (.RESET_B(net238),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0112_),
    .Q(\s0.shift_out[14] [0]),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6603_ (.RESET_B(net237),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0113_),
    .Q(\s0.data_out[14][0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6604_ (.RESET_B(net236),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0114_),
    .Q(\s0.data_out[14][1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6605_ (.RESET_B(net235),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0115_),
    .Q(\s0.data_out[14][2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6606_ (.RESET_B(net234),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0116_),
    .Q(\s0.data_out[14][3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6607_ (.RESET_B(net233),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0117_),
    .Q(\s0.data_out[14][4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6608_ (.RESET_B(net232),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0118_),
    .Q(\s0.data_out[14][5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6609_ (.RESET_B(net231),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net546),
    .Q(\s0.data_out[14][6] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6610_ (.RESET_B(net230),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0120_),
    .Q(\s0.data_out[14][7] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6611_ (.RESET_B(net229),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net567),
    .Q(\s0.was_valid_out[13] [0]),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6612_ (.RESET_B(net227),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0122_),
    .Q(\s0.valid_out[13] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6613_ (.RESET_B(net226),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0123_),
    .Q(\s0.genblk1[12].modules.bubble ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6614_ (.RESET_B(net225),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0124_),
    .Q(\s0.shift_out[13] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6615_ (.RESET_B(net224),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0125_),
    .Q(\s0.data_out[13][0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6616_ (.RESET_B(net223),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0126_),
    .Q(\s0.data_out[13][1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6617_ (.RESET_B(net222),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net458),
    .Q(\s0.data_out[13][2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6618_ (.RESET_B(net221),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net533),
    .Q(\s0.data_out[13][3] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6619_ (.RESET_B(net220),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0129_),
    .Q(\s0.data_out[13][4] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6620_ (.RESET_B(net219),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0130_),
    .Q(\s0.data_out[13][5] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6621_ (.RESET_B(net218),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\s0.data_out[13][6] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6622_ (.RESET_B(net217),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net407),
    .Q(\s0.data_out[13][7] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6623_ (.RESET_B(net216),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net349),
    .Q(\s0.was_valid_out[12] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6624_ (.RESET_B(net214),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0134_),
    .Q(\s0.valid_out[12] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6625_ (.RESET_B(net213),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0135_),
    .Q(\s0.shift_out[12] [0]),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6626_ (.RESET_B(net212),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0136_),
    .Q(\s0.data_out[12][0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6627_ (.RESET_B(net211),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net443),
    .Q(\s0.data_out[12][1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6628_ (.RESET_B(net210),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0138_),
    .Q(\s0.data_out[12][2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6629_ (.RESET_B(net209),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0139_),
    .Q(\s0.data_out[12][3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6630_ (.RESET_B(net208),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0140_),
    .Q(\s0.data_out[12][4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6631_ (.RESET_B(net207),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0141_),
    .Q(\s0.data_out[12][5] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6632_ (.RESET_B(net206),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net620),
    .Q(\s0.data_out[12][6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6633_ (.RESET_B(net205),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0143_),
    .Q(\s0.data_out[12][7] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6634_ (.RESET_B(net204),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net645),
    .Q(\s0.was_valid_out[11] [0]),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6635_ (.RESET_B(net202),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0145_),
    .Q(\s0.valid_out[11] [0]),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6636_ (.RESET_B(net201),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0146_),
    .Q(\s0.genblk1[11].modules.bubble ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6637_ (.RESET_B(net200),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0147_),
    .Q(\s0.genblk1[10].modules.bubble ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6638_ (.RESET_B(net199),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0148_),
    .Q(\s0.shift_out[11] [0]),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6639_ (.RESET_B(net198),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0149_),
    .Q(\s0.data_out[11][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6640_ (.RESET_B(net197),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0150_),
    .Q(\s0.data_out[11][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6641_ (.RESET_B(net196),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net423),
    .Q(\s0.data_out[11][2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6642_ (.RESET_B(net195),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net462),
    .Q(\s0.data_out[11][3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6643_ (.RESET_B(net194),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0153_),
    .Q(\s0.data_out[11][4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6644_ (.RESET_B(net193),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0154_),
    .Q(\s0.data_out[11][5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6645_ (.RESET_B(net192),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0155_),
    .Q(\s0.data_out[11][6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6646_ (.RESET_B(net191),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net452),
    .Q(\s0.data_out[11][7] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6647_ (.RESET_B(net190),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net351),
    .Q(\s0.was_valid_out[10] [0]),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6648_ (.RESET_B(net188),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0158_),
    .Q(\s0.valid_out[10] [0]),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6649_ (.RESET_B(net187),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0159_),
    .Q(\s0.data_new_delayed[0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6650_ (.RESET_B(net186),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0160_),
    .Q(\s0.data_new_delayed[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6651_ (.RESET_B(net185),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0161_),
    .Q(\s0.data_new_delayed[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6652_ (.RESET_B(net184),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0162_),
    .Q(\s0.data_new_delayed[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6653_ (.RESET_B(net183),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0163_),
    .Q(\s0.data_new_delayed[4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6654_ (.RESET_B(net182),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0164_),
    .Q(\s0.data_new_delayed[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6655_ (.RESET_B(net181),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0165_),
    .Q(\s0.data_new_delayed[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6656_ (.RESET_B(net180),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0166_),
    .Q(\s0.data_new_delayed[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6657_ (.RESET_B(net179),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0167_),
    .Q(\s0.shift_out[10] [0]),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6658_ (.RESET_B(net178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0168_),
    .Q(\s0.data_out[10][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6659_ (.RESET_B(net177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net490),
    .Q(\s0.data_out[10][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6660_ (.RESET_B(net176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0170_),
    .Q(\s0.data_out[10][2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6661_ (.RESET_B(net175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net478),
    .Q(\s0.data_out[10][3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6662_ (.RESET_B(net174),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0172_),
    .Q(\s0.data_out[10][4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6663_ (.RESET_B(net173),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0173_),
    .Q(\s0.data_out[10][5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6664_ (.RESET_B(net172),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0174_),
    .Q(\s0.data_out[10][6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6665_ (.RESET_B(net171),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0175_),
    .Q(\s0.data_out[10][7] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6666_ (.RESET_B(net170),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net667),
    .Q(\s0.was_valid_out[9] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6667_ (.RESET_B(net168),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0177_),
    .Q(\s0.valid_out[9] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6668_ (.RESET_B(net167),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0178_),
    .Q(\s0.genblk1[8].modules.bubble ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6669_ (.RESET_B(net166),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0179_),
    .Q(\s0.shift_out[9] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6670_ (.RESET_B(net165),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0180_),
    .Q(\s0.data_out[9][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6671_ (.RESET_B(net164),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net573),
    .Q(\s0.data_out[9][1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6672_ (.RESET_B(net163),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net466),
    .Q(\s0.data_out[9][2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6673_ (.RESET_B(net162),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net590),
    .Q(\s0.data_out[9][3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6674_ (.RESET_B(net161),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0184_),
    .Q(\s0.data_out[9][4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6675_ (.RESET_B(net160),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0185_),
    .Q(\s0.data_out[9][5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6676_ (.RESET_B(net159),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net510),
    .Q(\s0.data_out[9][6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6677_ (.RESET_B(net158),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0187_),
    .Q(\s0.data_out[9][7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6678_ (.RESET_B(net157),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net359),
    .Q(\s0.was_valid_out[8] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6679_ (.RESET_B(net155),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0189_),
    .Q(\s0.valid_out[8] [0]),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6680_ (.RESET_B(net154),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0190_),
    .Q(\s0.genblk1[7].modules.bubble ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6681_ (.RESET_B(net153),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0191_),
    .Q(\s0.shift_out[8] [0]),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6682_ (.RESET_B(net152),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\s0.data_out[8][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6683_ (.RESET_B(net151),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0193_),
    .Q(\s0.data_out[8][1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6684_ (.RESET_B(net150),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0194_),
    .Q(\s0.data_out[8][2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6685_ (.RESET_B(net149),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net638),
    .Q(\s0.data_out[8][3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6686_ (.RESET_B(net148),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net671),
    .Q(\s0.data_out[8][4] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6687_ (.RESET_B(net147),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net688),
    .Q(\s0.data_out[8][5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6688_ (.RESET_B(net146),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0198_),
    .Q(\s0.data_out[8][6] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6689_ (.RESET_B(net145),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0199_),
    .Q(\s0.data_out[8][7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6690_ (.RESET_B(net144),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0200_),
    .Q(\s0.was_valid_out[7] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6691_ (.RESET_B(net142),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0201_),
    .Q(\s0.valid_out[7] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6692_ (.RESET_B(net141),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0202_),
    .Q(\s0.genblk1[6].modules.bubble ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6693_ (.RESET_B(net140),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0203_),
    .Q(\s0.shift_out[7] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6694_ (.RESET_B(net139),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0204_),
    .Q(\s0.data_out[7][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6695_ (.RESET_B(net138),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net409),
    .Q(\s0.data_out[7][1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6696_ (.RESET_B(net137),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net454),
    .Q(\s0.data_out[7][2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6697_ (.RESET_B(net136),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0207_),
    .Q(\s0.data_out[7][3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6698_ (.RESET_B(net135),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0208_),
    .Q(\s0.data_out[7][4] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6699_ (.RESET_B(net134),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net471),
    .Q(\s0.data_out[7][5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6700_ (.RESET_B(net133),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0210_),
    .Q(\s0.data_out[7][6] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6701_ (.RESET_B(net132),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0211_),
    .Q(\s0.data_out[7][7] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6702_ (.RESET_B(net131),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0212_),
    .Q(\s0.was_valid_out[6] [0]),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6703_ (.RESET_B(net129),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0213_),
    .Q(\s0.valid_out[6] [0]),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6704_ (.RESET_B(net128),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0214_),
    .Q(\s0.genblk1[5].modules.bubble ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6705_ (.RESET_B(net127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0215_),
    .Q(\s0.shift_out[6] [0]),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6706_ (.RESET_B(net126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0216_),
    .Q(\s0.data_out[6][0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6707_ (.RESET_B(net125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net502),
    .Q(\s0.data_out[6][1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6708_ (.RESET_B(net124),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0218_),
    .Q(\s0.data_out[6][2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6709_ (.RESET_B(net123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net448),
    .Q(\s0.data_out[6][3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6710_ (.RESET_B(net122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0220_),
    .Q(\s0.data_out[6][4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6711_ (.RESET_B(net121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0221_),
    .Q(\s0.data_out[6][5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6712_ (.RESET_B(net120),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0222_),
    .Q(\s0.data_out[6][6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6713_ (.RESET_B(net119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0223_),
    .Q(\s0.data_out[6][7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6714_ (.RESET_B(net118),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net346),
    .Q(\s0.was_valid_out[5] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6715_ (.RESET_B(net116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0225_),
    .Q(\s0.valid_out[5] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6716_ (.RESET_B(net115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0226_),
    .Q(\s0.genblk1[4].modules.bubble ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6717_ (.RESET_B(net114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0227_),
    .Q(\s0.shift_out[5] [0]),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6718_ (.RESET_B(net113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0228_),
    .Q(\s0.data_out[5][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6719_ (.RESET_B(net112),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0229_),
    .Q(\s0.data_out[5][1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6720_ (.RESET_B(net111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0230_),
    .Q(\s0.data_out[5][2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6721_ (.RESET_B(net110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0231_),
    .Q(\s0.data_out[5][3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6722_ (.RESET_B(net109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0232_),
    .Q(\s0.data_out[5][4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6723_ (.RESET_B(net108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0233_),
    .Q(\s0.data_out[5][5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6724_ (.RESET_B(net107),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net450),
    .Q(\s0.data_out[5][6] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6725_ (.RESET_B(net106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0235_),
    .Q(\s0.data_out[5][7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6726_ (.RESET_B(net105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0236_),
    .Q(\s0.was_valid_out[4] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6727_ (.RESET_B(net103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0237_),
    .Q(\s0.valid_out[4] [0]),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6728_ (.RESET_B(net102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0238_),
    .Q(\s0.genblk1[3].modules.bubble ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6729_ (.RESET_B(net101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0239_),
    .Q(\s0.shift_out[4] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6730_ (.RESET_B(net100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0240_),
    .Q(\s0.data_out[4][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6731_ (.RESET_B(net99),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0241_),
    .Q(\s0.data_out[4][1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6732_ (.RESET_B(net98),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0242_),
    .Q(\s0.data_out[4][2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6733_ (.RESET_B(net97),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net445),
    .Q(\s0.data_out[4][3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6734_ (.RESET_B(net96),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0244_),
    .Q(\s0.data_out[4][4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6735_ (.RESET_B(net95),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0245_),
    .Q(\s0.data_out[4][5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6736_ (.RESET_B(net94),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net508),
    .Q(\s0.data_out[4][6] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6737_ (.RESET_B(net93),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net493),
    .Q(\s0.data_out[4][7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6738_ (.RESET_B(net92),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0248_),
    .Q(\s0.was_valid_out[3] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6739_ (.RESET_B(net90),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0249_),
    .Q(\s0.valid_out[3] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6740_ (.RESET_B(net89),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0250_),
    .Q(\s0.genblk1[2].modules.bubble ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6741_ (.RESET_B(net88),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0251_),
    .Q(\s0.shift_out[3] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6742_ (.RESET_B(net87),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0252_),
    .Q(\s0.data_out[3][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6743_ (.RESET_B(net86),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net401),
    .Q(\s0.data_out[3][1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6744_ (.RESET_B(net85),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net435),
    .Q(\s0.data_out[3][2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6745_ (.RESET_B(net84),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net575),
    .Q(\s0.data_out[3][3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6746_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0256_),
    .Q(\s0.data_out[3][4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6747_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0257_),
    .Q(\s0.data_out[3][5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6748_ (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0258_),
    .Q(\s0.data_out[3][6] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _6749_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net485),
    .Q(\s0.data_out[3][7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6750_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net357),
    .Q(\s0.was_valid_out[2] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6751_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0261_),
    .Q(\s0.valid_out[2] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6752_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0262_),
    .Q(\s0.genblk1[23].modules.bubble ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6753_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0263_),
    .Q(\s0.shift_out[2] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6754_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0264_),
    .Q(\s0.data_out[2][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6755_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net515),
    .Q(\s0.data_out[2][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6756_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0266_),
    .Q(\s0.data_out[2][2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6757_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net464),
    .Q(\s0.data_out[2][3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6758_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0268_),
    .Q(\s0.data_out[2][4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6759_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0269_),
    .Q(\s0.data_out[2][5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6760_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net581),
    .Q(\s0.data_out[2][6] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _6761_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net513),
    .Q(\s0.data_out[2][7] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6762_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net517),
    .Q(\s0.was_valid_out[1] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6763_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0273_),
    .Q(\s0.valid_out[1] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6764_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0274_),
    .Q(\s0.genblk1[19].modules.bubble ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6765_ (.RESET_B(net49),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0275_),
    .Q(\s0.shift_out[1] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _6766_ (.RESET_B(net36),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0276_),
    .Q(\s0.data_out[1][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6767_ (.RESET_B(net23),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net495),
    .Q(\s0.data_out[1][1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6768_ (.RESET_B(net306),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0278_),
    .Q(\s0.data_out[1][2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6769_ (.RESET_B(net293),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0279_),
    .Q(\s0.data_out[1][3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6770_ (.RESET_B(net280),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0280_),
    .Q(\s0.data_out[1][4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6771_ (.RESET_B(net267),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0281_),
    .Q(\s0.data_out[1][5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6772_ (.RESET_B(net254),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0282_),
    .Q(\s0.data_out[1][6] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _6773_ (.RESET_B(net241),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0283_),
    .Q(\s0.data_out[1][7] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6774_ (.RESET_B(net228),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0284_),
    .Q(\s0.was_valid_out[0] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6775_ (.RESET_B(net203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0285_),
    .Q(\s0.valid_out[0] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6776_ (.RESET_B(net189),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0286_),
    .Q(\s0.genblk1[9].modules.bubble ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6777_ (.RESET_B(net169),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0287_),
    .Q(\s0.shift_out[0] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6778_ (.RESET_B(net156),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0288_),
    .Q(\s0.data_out[0][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6779_ (.RESET_B(net143),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net376),
    .Q(\s0.data_out[0][1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6780_ (.RESET_B(net130),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0290_),
    .Q(\s0.data_out[0][2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6781_ (.RESET_B(net117),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net403),
    .Q(\s0.data_out[0][3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6782_ (.RESET_B(net104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0292_),
    .Q(\s0.data_out[0][4] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6783_ (.RESET_B(net91),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0293_),
    .Q(\s0.data_out[0][5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6784_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0294_),
    .Q(\s0.data_out[0][6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6785_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0295_),
    .Q(\s0.data_out[0][7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_tiehi _6527__24 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net24));
 sg13g2_tiehi _6526__25 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net25));
 sg13g2_tiehi _6525__26 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net26));
 sg13g2_tiehi _6524__27 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net27));
 sg13g2_tiehi _6523__28 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net28));
 sg13g2_tiehi _6522__29 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net29));
 sg13g2_tiehi _6521__30 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net30));
 sg13g2_tiehi _6520__31 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net31));
 sg13g2_tiehi _6519__32 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net32));
 sg13g2_tiehi _6518__33 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net33));
 sg13g2_tiehi _6517__34 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net34));
 sg13g2_tiehi _6516__35 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net35));
 sg13g2_tiehi _6766__36 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net36));
 sg13g2_tiehi _6515__37 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net37));
 sg13g2_tiehi _6514__38 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_tiehi _6513__39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi _6512__40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_tiehi _6511__41 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net41));
 sg13g2_tiehi _6510__42 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net42));
 sg13g2_tiehi _6509__43 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net43));
 sg13g2_tiehi _6508__44 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net44));
 sg13g2_tiehi _6507__45 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net45));
 sg13g2_tiehi _6506__46 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net46));
 sg13g2_tiehi _6505__47 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net47));
 sg13g2_tiehi _6504__48 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net48));
 sg13g2_tiehi _6765__49 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net49));
 sg13g2_tiehi _6503__50 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net50));
 sg13g2_tiehi _6502__51 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net51));
 sg13g2_tiehi _6501__52 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net52));
 sg13g2_tiehi _6500__53 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net53));
 sg13g2_tiehi _6499__54 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net54));
 sg13g2_tiehi _6498__55 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net55));
 sg13g2_tiehi _6497__56 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net56));
 sg13g2_tiehi _6496__57 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net57));
 sg13g2_tiehi _6495__58 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net58));
 sg13g2_tiehi _6494__59 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net59));
 sg13g2_tiehi _6493__60 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net60));
 sg13g2_tiehi _6492__61 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net61));
 sg13g2_tiehi _6764__62 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net62));
 sg13g2_tiehi _6491__63 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net63));
 sg13g2_tiehi _6763__64 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net64));
 sg13g2_tiehi _6785__65 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net65));
 sg13g2_tiehi _6762__66 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net66));
 sg13g2_tiehi _6761__67 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net67));
 sg13g2_tiehi _6760__68 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net68));
 sg13g2_tiehi _6759__69 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net69));
 sg13g2_tiehi _6758__70 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net70));
 sg13g2_tiehi _6757__71 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net71));
 sg13g2_tiehi _6756__72 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net72));
 sg13g2_tiehi _6755__73 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net73));
 sg13g2_tiehi _6754__74 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net74));
 sg13g2_tiehi _6753__75 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net75));
 sg13g2_tiehi _6752__76 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net76));
 sg13g2_tiehi _6751__77 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net77));
 sg13g2_tiehi _6784__78 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net78));
 sg13g2_tiehi _6750__79 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net79));
 sg13g2_tiehi _6749__80 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net80));
 sg13g2_tiehi _6748__81 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net81));
 sg13g2_tiehi _6747__82 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net82));
 sg13g2_tiehi _6746__83 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net83));
 sg13g2_tiehi _6745__84 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net84));
 sg13g2_tiehi _6744__85 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net85));
 sg13g2_tiehi _6743__86 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net86));
 sg13g2_tiehi _6742__87 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net87));
 sg13g2_tiehi _6741__88 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net88));
 sg13g2_tiehi _6740__89 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net89));
 sg13g2_tiehi _6739__90 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net90));
 sg13g2_tiehi _6783__91 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net91));
 sg13g2_tiehi _6738__92 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net92));
 sg13g2_tiehi _6737__93 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net93));
 sg13g2_tiehi _6736__94 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net94));
 sg13g2_tiehi _6735__95 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net95));
 sg13g2_tiehi _6734__96 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net96));
 sg13g2_tiehi _6733__97 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net97));
 sg13g2_tiehi _6732__98 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net98));
 sg13g2_tiehi _6731__99 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net99));
 sg13g2_tiehi _6730__100 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net100));
 sg13g2_tiehi _6729__101 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net101));
 sg13g2_tiehi _6728__102 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net102));
 sg13g2_tiehi _6727__103 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net103));
 sg13g2_tiehi _6782__104 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net104));
 sg13g2_tiehi _6726__105 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net105));
 sg13g2_tiehi _6725__106 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net106));
 sg13g2_tiehi _6724__107 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net107));
 sg13g2_tiehi _6723__108 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net108));
 sg13g2_tiehi _6722__109 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net109));
 sg13g2_tiehi _6721__110 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net110));
 sg13g2_tiehi _6720__111 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net111));
 sg13g2_tiehi _6719__112 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net112));
 sg13g2_tiehi _6718__113 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net113));
 sg13g2_tiehi _6717__114 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net114));
 sg13g2_tiehi _6716__115 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net115));
 sg13g2_tiehi _6715__116 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net116));
 sg13g2_tiehi _6781__117 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net117));
 sg13g2_tiehi _6714__118 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net118));
 sg13g2_tiehi _6713__119 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net119));
 sg13g2_tiehi _6712__120 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net120));
 sg13g2_tiehi _6711__121 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net121));
 sg13g2_tiehi _6710__122 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net122));
 sg13g2_tiehi _6709__123 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net123));
 sg13g2_tiehi _6708__124 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net124));
 sg13g2_tiehi _6707__125 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net125));
 sg13g2_tiehi _6706__126 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net126));
 sg13g2_tiehi _6705__127 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net127));
 sg13g2_tiehi _6704__128 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net128));
 sg13g2_tiehi _6703__129 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net129));
 sg13g2_tiehi _6780__130 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net130));
 sg13g2_tiehi _6702__131 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net131));
 sg13g2_tiehi _6701__132 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net132));
 sg13g2_tiehi _6700__133 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net133));
 sg13g2_tiehi _6699__134 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net134));
 sg13g2_tiehi _6698__135 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net135));
 sg13g2_tiehi _6697__136 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net136));
 sg13g2_tiehi _6696__137 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net137));
 sg13g2_tiehi _6695__138 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net138));
 sg13g2_tiehi _6694__139 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net139));
 sg13g2_tiehi _6693__140 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net140));
 sg13g2_tiehi _6692__141 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net141));
 sg13g2_tiehi _6691__142 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net142));
 sg13g2_tiehi _6779__143 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net143));
 sg13g2_tiehi _6690__144 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net144));
 sg13g2_tiehi _6689__145 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net145));
 sg13g2_tiehi _6688__146 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net146));
 sg13g2_tiehi _6687__147 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net147));
 sg13g2_tiehi _6686__148 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net148));
 sg13g2_tiehi _6685__149 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net149));
 sg13g2_tiehi _6684__150 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net150));
 sg13g2_tiehi _6683__151 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net151));
 sg13g2_tiehi _6682__152 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net152));
 sg13g2_tiehi _6681__153 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net153));
 sg13g2_tiehi _6680__154 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net154));
 sg13g2_tiehi _6679__155 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net155));
 sg13g2_tiehi _6778__156 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net156));
 sg13g2_tiehi _6678__157 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net157));
 sg13g2_tiehi _6677__158 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net158));
 sg13g2_tiehi _6676__159 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net159));
 sg13g2_tiehi _6675__160 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net160));
 sg13g2_tiehi _6674__161 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net161));
 sg13g2_tiehi _6673__162 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net162));
 sg13g2_tiehi _6672__163 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net163));
 sg13g2_tiehi _6671__164 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net164));
 sg13g2_tiehi _6670__165 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net165));
 sg13g2_tiehi _6669__166 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net166));
 sg13g2_tiehi _6668__167 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net167));
 sg13g2_tiehi _6667__168 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net168));
 sg13g2_tiehi _6777__169 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net169));
 sg13g2_tiehi _6666__170 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net170));
 sg13g2_tiehi _6665__171 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net171));
 sg13g2_tiehi _6664__172 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net172));
 sg13g2_tiehi _6663__173 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net173));
 sg13g2_tiehi _6662__174 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net174));
 sg13g2_tiehi _6661__175 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net175));
 sg13g2_tiehi _6660__176 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net176));
 sg13g2_tiehi _6659__177 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net177));
 sg13g2_tiehi _6658__178 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net178));
 sg13g2_tiehi _6657__179 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net179));
 sg13g2_tiehi _6656__180 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net180));
 sg13g2_tiehi _6655__181 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net181));
 sg13g2_tiehi _6654__182 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net182));
 sg13g2_tiehi _6653__183 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net183));
 sg13g2_tiehi _6652__184 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net184));
 sg13g2_tiehi _6651__185 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net185));
 sg13g2_tiehi _6650__186 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net186));
 sg13g2_tiehi _6649__187 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net187));
 sg13g2_tiehi _6648__188 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net188));
 sg13g2_tiehi _6776__189 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net189));
 sg13g2_tiehi _6647__190 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net190));
 sg13g2_tiehi _6646__191 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net191));
 sg13g2_tiehi _6645__192 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net192));
 sg13g2_tiehi _6644__193 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net193));
 sg13g2_tiehi _6643__194 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net194));
 sg13g2_tiehi _6642__195 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net195));
 sg13g2_tiehi _6641__196 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net196));
 sg13g2_tiehi _6640__197 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net197));
 sg13g2_tiehi _6639__198 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net198));
 sg13g2_tiehi _6638__199 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net199));
 sg13g2_tiehi _6637__200 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net200));
 sg13g2_tiehi _6636__201 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net201));
 sg13g2_tiehi _6635__202 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net202));
 sg13g2_tiehi _6775__203 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net203));
 sg13g2_tiehi _6634__204 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net204));
 sg13g2_tiehi _6633__205 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net205));
 sg13g2_tiehi _6632__206 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net206));
 sg13g2_tiehi _6631__207 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net207));
 sg13g2_tiehi _6630__208 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net208));
 sg13g2_tiehi _6629__209 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net209));
 sg13g2_tiehi _6628__210 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net210));
 sg13g2_tiehi _6627__211 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net211));
 sg13g2_tiehi _6626__212 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net212));
 sg13g2_tiehi _6625__213 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net213));
 sg13g2_tiehi _6624__214 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net214));
 sg13g2_tiehi _6490__215 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net215));
 sg13g2_tiehi _6623__216 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net216));
 sg13g2_tiehi _6622__217 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net217));
 sg13g2_tiehi _6621__218 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net218));
 sg13g2_tiehi _6620__219 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net219));
 sg13g2_tiehi _6619__220 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net220));
 sg13g2_tiehi _6618__221 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net221));
 sg13g2_tiehi _6617__222 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net222));
 sg13g2_tiehi _6616__223 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net223));
 sg13g2_tiehi _6615__224 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net224));
 sg13g2_tiehi _6614__225 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net225));
 sg13g2_tiehi _6613__226 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net226));
 sg13g2_tiehi _6612__227 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net227));
 sg13g2_tiehi _6774__228 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net228));
 sg13g2_tiehi _6611__229 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net229));
 sg13g2_tiehi _6610__230 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net230));
 sg13g2_tiehi _6609__231 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net231));
 sg13g2_tiehi _6608__232 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net232));
 sg13g2_tiehi _6607__233 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net233));
 sg13g2_tiehi _6606__234 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net234));
 sg13g2_tiehi _6605__235 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net235));
 sg13g2_tiehi _6604__236 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net236));
 sg13g2_tiehi _6603__237 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net237));
 sg13g2_tiehi _6602__238 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net238));
 sg13g2_tiehi _6601__239 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net239));
 sg13g2_tiehi _6600__240 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net240));
 sg13g2_tiehi _6773__241 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net241));
 sg13g2_tiehi _6599__242 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net242));
 sg13g2_tiehi _6598__243 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net243));
 sg13g2_tiehi _6597__244 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net244));
 sg13g2_tiehi _6596__245 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net245));
 sg13g2_tiehi _6595__246 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net246));
 sg13g2_tiehi _6594__247 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net247));
 sg13g2_tiehi _6593__248 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net248));
 sg13g2_tiehi _6592__249 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net249));
 sg13g2_tiehi _6591__250 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net250));
 sg13g2_tiehi _6590__251 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net251));
 sg13g2_tiehi _6589__252 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net252));
 sg13g2_tiehi _6588__253 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net253));
 sg13g2_tiehi _6772__254 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net254));
 sg13g2_tiehi _6587__255 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net255));
 sg13g2_tiehi _6586__256 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net256));
 sg13g2_tiehi _6585__257 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net257));
 sg13g2_tiehi _6584__258 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net258));
 sg13g2_tiehi _6583__259 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net259));
 sg13g2_tiehi _6582__260 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net260));
 sg13g2_tiehi _6581__261 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net261));
 sg13g2_tiehi _6580__262 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net262));
 sg13g2_tiehi _6579__263 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net263));
 sg13g2_tiehi _6578__264 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net264));
 sg13g2_tiehi _6577__265 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net265));
 sg13g2_tiehi _6576__266 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net266));
 sg13g2_tiehi _6771__267 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net267));
 sg13g2_tiehi _6575__268 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net268));
 sg13g2_tiehi _6574__269 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net269));
 sg13g2_tiehi _6573__270 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net270));
 sg13g2_tiehi _6572__271 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net271));
 sg13g2_tiehi _6571__272 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net272));
 sg13g2_tiehi _6570__273 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net273));
 sg13g2_tiehi _6569__274 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net274));
 sg13g2_tiehi _6568__275 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net275));
 sg13g2_tiehi _6567__276 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net276));
 sg13g2_tiehi _6566__277 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net277));
 sg13g2_tiehi _6565__278 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net278));
 sg13g2_tiehi _6564__279 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net279));
 sg13g2_tiehi _6770__280 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net280));
 sg13g2_tiehi _6563__281 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net281));
 sg13g2_tiehi _6562__282 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net282));
 sg13g2_tiehi _6561__283 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net283));
 sg13g2_tiehi _6560__284 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net284));
 sg13g2_tiehi _6559__285 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net285));
 sg13g2_tiehi _6558__286 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net286));
 sg13g2_tiehi _6557__287 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net287));
 sg13g2_tiehi _6556__288 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net288));
 sg13g2_tiehi _6555__289 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net289));
 sg13g2_tiehi _6554__290 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net290));
 sg13g2_tiehi _6553__291 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net291));
 sg13g2_tiehi _6552__292 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net292));
 sg13g2_tiehi _6769__293 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net293));
 sg13g2_tiehi _6551__294 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net294));
 sg13g2_tiehi _6550__295 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net295));
 sg13g2_tiehi _6549__296 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net296));
 sg13g2_tiehi _6548__297 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net297));
 sg13g2_tiehi _6547__298 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net298));
 sg13g2_tiehi _6546__299 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net299));
 sg13g2_tiehi _6545__300 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net300));
 sg13g2_tiehi _6544__301 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net301));
 sg13g2_tiehi _6543__302 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net302));
 sg13g2_tiehi _6542__303 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net303));
 sg13g2_tiehi _6541__304 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net304));
 sg13g2_tiehi _6540__305 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net305));
 sg13g2_tiehi _6768__306 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net306));
 sg13g2_tiehi _6539__307 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net307));
 sg13g2_tiehi _6538__308 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net308));
 sg13g2_tiehi _6537__309 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net309));
 sg13g2_tiehi _6536__310 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net310));
 sg13g2_tiehi _6535__311 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net311));
 sg13g2_tiehi _6534__312 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net312));
 sg13g2_tiehi _6533__313 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net313));
 sg13g2_tiehi _6532__314 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net314));
 sg13g2_tiehi _6531__315 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net315));
 sg13g2_tiehi _6530__316 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net316));
 sg13g2_tiehi _6529__317 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net317));
 sg13g2_tiehi _6528__318 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net318));
 sg13g2_tiehi heichips25_top_sorter_319 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net319));
 sg13g2_tiehi heichips25_top_sorter_320 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net320));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_top_sorter_11 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net11));
 sg13g2_tielo heichips25_top_sorter_12 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net12));
 sg13g2_tielo heichips25_top_sorter_13 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net13));
 sg13g2_tielo heichips25_top_sorter_14 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net14));
 sg13g2_tielo heichips25_top_sorter_15 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net15));
 sg13g2_tielo heichips25_top_sorter_16 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net16));
 sg13g2_tielo heichips25_top_sorter_17 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net17));
 sg13g2_tielo heichips25_top_sorter_18 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net18));
 sg13g2_tielo heichips25_top_sorter_19 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net19));
 sg13g2_tielo heichips25_top_sorter_20 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net20));
 sg13g2_tielo heichips25_top_sorter_21 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net21));
 sg13g2_tielo heichips25_top_sorter_22 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net22));
 sg13g2_tiehi _6767__23 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net23));
 sg13g2_buf_1 _7097_ (.A(\s0.was_valid_out[23] [0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout991 (.A(net992),
    .X(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout992 (.A(_2885_),
    .X(net992),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout993 (.A(_2772_),
    .X(net993),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout994 (.A(_2772_),
    .X(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout995 (.A(_2762_),
    .X(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout996 (.A(_2762_),
    .X(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout997 (.A(net998),
    .X(net997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout998 (.A(_2761_),
    .X(net998),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout999 (.A(_2761_),
    .X(net999),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1000 (.A(_2759_),
    .X(net1000),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1001 (.A(_2758_),
    .X(net1001),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1002 (.A(_2757_),
    .X(net1002),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1003 (.A(_2755_),
    .X(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1004 (.A(net1006),
    .X(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1005 (.A(net1006),
    .X(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1006 (.A(_2754_),
    .X(net1006),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1007 (.A(net1008),
    .X(net1007),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1008 (.A(_2752_),
    .X(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1009 (.A(net1010),
    .X(net1009),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1010 (.A(_2751_),
    .X(net1010),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1011 (.A(_2749_),
    .X(net1011),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1012 (.A(_2749_),
    .X(net1012),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1013 (.A(_2746_),
    .X(net1013),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1014 (.A(_2746_),
    .X(net1014),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1015 (.A(net1016),
    .X(net1015),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1016 (.A(_2744_),
    .X(net1016),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1017 (.A(_2741_),
    .X(net1017),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1018 (.A(_2741_),
    .X(net1018),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1019 (.A(net1021),
    .X(net1019),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1020 (.A(net1021),
    .X(net1020),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1021 (.A(net397),
    .X(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1022 (.A(net1023),
    .X(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1023 (.A(net397),
    .X(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1024 (.A(net1026),
    .X(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1025 (.A(net1026),
    .X(net1025),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1026 (.A(\s0.valid_out[0] [0]),
    .X(net1026),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1027 (.A(net1029),
    .X(net1027),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1028 (.A(net1029),
    .X(net1028),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1029 (.A(\s0.shift_out[1] [0]),
    .X(net1029),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1030 (.A(net1032),
    .X(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1031 (.A(net710),
    .X(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1032 (.A(\s0.shift_out[1] [0]),
    .X(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1033 (.A(net1035),
    .X(net1033),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1034 (.A(net1035),
    .X(net1034),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1035 (.A(\s0.valid_out[1] [0]),
    .X(net1035),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1036 (.A(net1042),
    .X(net1036),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1037 (.A(net1042),
    .X(net1037),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1038 (.A(net1042),
    .X(net1038),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1039 (.A(net1041),
    .X(net1039),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1040 (.A(net1041),
    .X(net1040),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1041 (.A(net1042),
    .X(net1041),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1042 (.A(\s0.shift_out[2] [0]),
    .X(net1042),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1043 (.A(net1046),
    .X(net1043),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1044 (.A(net1046),
    .X(net1044),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1045 (.A(net1046),
    .X(net1045),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1046 (.A(net396),
    .X(net1046),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1047 (.A(net1055),
    .X(net1047),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1048 (.A(net1055),
    .X(net1048),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1049 (.A(net1050),
    .X(net1049),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1050 (.A(net1055),
    .X(net1050),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1051 (.A(net1054),
    .X(net1051),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1052 (.A(net1054),
    .X(net1052),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1053 (.A(net1054),
    .X(net1053),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1054 (.A(net1055),
    .X(net1054),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1055 (.A(net585),
    .X(net1055),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1056 (.A(net1059),
    .X(net1056),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1057 (.A(net1059),
    .X(net1057),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1058 (.A(net1059),
    .X(net1058),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1059 (.A(\s0.valid_out[3] [0]),
    .X(net1059),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1060 (.A(net1063),
    .X(net1060),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1061 (.A(net1063),
    .X(net1061),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1062 (.A(net1063),
    .X(net1062),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1063 (.A(net608),
    .X(net1063),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1064 (.A(net1066),
    .X(net1064),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1065 (.A(net1066),
    .X(net1065),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1066 (.A(net608),
    .X(net1066),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1067 (.A(net1071),
    .X(net1067),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1068 (.A(net1071),
    .X(net1068),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1069 (.A(net1071),
    .X(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1070 (.A(net1071),
    .X(net1070),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1071 (.A(net706),
    .X(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1072 (.A(net1073),
    .X(net1072),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1073 (.A(net384),
    .X(net1073),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1074 (.A(net1075),
    .X(net1074),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1075 (.A(net384),
    .X(net1075),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1076 (.A(net1077),
    .X(net1076),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1077 (.A(net1079),
    .X(net1077),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1078 (.A(net1079),
    .X(net1078),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1079 (.A(\s0.shift_out[5] [0]),
    .X(net1079),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1080 (.A(net1084),
    .X(net1080),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1081 (.A(net1084),
    .X(net1081),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1082 (.A(net1084),
    .X(net1082),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1083 (.A(net1084),
    .X(net1083),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1084 (.A(net711),
    .X(net1084),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1085 (.A(net1087),
    .X(net1085),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1086 (.A(net1087),
    .X(net1086),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1087 (.A(net1091),
    .X(net1087),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1088 (.A(net1090),
    .X(net1088),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1089 (.A(net1090),
    .X(net1089),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1090 (.A(net1091),
    .X(net1090),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1091 (.A(net446),
    .X(net1091),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1092 (.A(\s0.valid_out[6] [0]),
    .X(net1092),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1093 (.A(\s0.valid_out[6] [0]),
    .X(net1093),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1094 (.A(net1095),
    .X(net1094),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1095 (.A(\s0.valid_out[6] [0]),
    .X(net1095),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1096 (.A(net1097),
    .X(net1096),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1097 (.A(net1104),
    .X(net1097),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1098 (.A(net1099),
    .X(net1098),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1099 (.A(net1104),
    .X(net1099),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1100 (.A(net1101),
    .X(net1100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1101 (.A(net1104),
    .X(net1101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1102 (.A(net1104),
    .X(net1102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1103 (.A(net1104),
    .X(net1103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1104 (.A(net563),
    .X(net1104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1105 (.A(net1109),
    .X(net1105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1106 (.A(net1109),
    .X(net1106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1107 (.A(net1109),
    .X(net1107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1108 (.A(net1109),
    .X(net1108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1109 (.A(\s0.valid_out[7] [0]),
    .X(net1109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1110 (.A(net1112),
    .X(net1110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1111 (.A(net1112),
    .X(net1111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1112 (.A(net1113),
    .X(net1112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1113 (.A(\s0.shift_out[8] [0]),
    .X(net1113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1114 (.A(net1117),
    .X(net1114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1115 (.A(net1117),
    .X(net1115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1116 (.A(net1117),
    .X(net1116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1117 (.A(\s0.shift_out[8] [0]),
    .X(net1117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1118 (.A(net1119),
    .X(net1118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1119 (.A(\s0.valid_out[8] [0]),
    .X(net1119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1120 (.A(\s0.valid_out[8] [0]),
    .X(net1120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1121 (.A(\s0.valid_out[8] [0]),
    .X(net1121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1122 (.A(net1123),
    .X(net1122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1123 (.A(net1127),
    .X(net1123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1124 (.A(net1127),
    .X(net1124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1125 (.A(net1126),
    .X(net1125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1126 (.A(net1127),
    .X(net1126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1127 (.A(\s0.shift_out[9] [0]),
    .X(net1127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1128 (.A(net1129),
    .X(net1128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1129 (.A(net1130),
    .X(net1129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1130 (.A(\s0.shift_out[9] [0]),
    .X(net1130),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1131 (.A(net1133),
    .X(net1131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1132 (.A(net1133),
    .X(net1132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1133 (.A(net1134),
    .X(net1133),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1134 (.A(\s0.valid_out[9] [0]),
    .X(net1134),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1135 (.A(net1136),
    .X(net1135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1136 (.A(net1137),
    .X(net1136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1137 (.A(net1141),
    .X(net1137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1138 (.A(net1141),
    .X(net1138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1139 (.A(net1141),
    .X(net1139),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1140 (.A(net1141),
    .X(net1140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1141 (.A(net360),
    .X(net1141),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1142 (.A(net1146),
    .X(net1142),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1143 (.A(net1146),
    .X(net1143),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1144 (.A(net1146),
    .X(net1144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1145 (.A(net1146),
    .X(net1145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1146 (.A(net707),
    .X(net1146),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1147 (.A(net1150),
    .X(net1147),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1148 (.A(net1150),
    .X(net1148),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1149 (.A(net1150),
    .X(net1149),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1150 (.A(net709),
    .X(net1150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1151 (.A(net1155),
    .X(net1151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1152 (.A(net1155),
    .X(net1152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1153 (.A(net1155),
    .X(net1153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1154 (.A(net1155),
    .X(net1154),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1155 (.A(net708),
    .X(net1155),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1156 (.A(net1160),
    .X(net1156),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1157 (.A(net1160),
    .X(net1157),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1158 (.A(net1160),
    .X(net1158),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1159 (.A(net1160),
    .X(net1159),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1160 (.A(net704),
    .X(net1160),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1161 (.A(\s0.data_new_delayed[3] ),
    .X(net1161),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1162 (.A(net700),
    .X(net1162),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1163 (.A(\s0.data_new_delayed[2] ),
    .X(net1163),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1164 (.A(net1165),
    .X(net1164),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1165 (.A(\s0.data_new_delayed[2] ),
    .X(net1165),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1166 (.A(net702),
    .X(net1166),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1167 (.A(\s0.data_new_delayed[1] ),
    .X(net1167),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1168 (.A(net1169),
    .X(net1168),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1169 (.A(\s0.data_new_delayed[1] ),
    .X(net1169),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1170 (.A(net1173),
    .X(net1170),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1171 (.A(net1172),
    .X(net1171),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1172 (.A(net1173),
    .X(net1172),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1173 (.A(net705),
    .X(net1173),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1174 (.A(net1177),
    .X(net1174),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1175 (.A(net1176),
    .X(net1175),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1176 (.A(net1177),
    .X(net1176),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1177 (.A(\s0.valid_out[10] [0]),
    .X(net1177),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1178 (.A(net1180),
    .X(net1178),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1179 (.A(net1180),
    .X(net1179),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1180 (.A(net1181),
    .X(net1180),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1181 (.A(net1186),
    .X(net1181),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1182 (.A(net1183),
    .X(net1182),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1183 (.A(net1186),
    .X(net1183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1184 (.A(net1185),
    .X(net1184),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1185 (.A(net1186),
    .X(net1185),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1186 (.A(\s0.shift_out[11] [0]),
    .X(net1186),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1187 (.A(net1190),
    .X(net1187),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1188 (.A(net1190),
    .X(net1188),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1189 (.A(net1190),
    .X(net1189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1190 (.A(\s0.valid_out[11] [0]),
    .X(net1190),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1191 (.A(net1192),
    .X(net1191),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1192 (.A(net1193),
    .X(net1192),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1193 (.A(net391),
    .X(net1193),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1194 (.A(net391),
    .X(net1194),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1195 (.A(net1196),
    .X(net1195),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1196 (.A(net391),
    .X(net1196),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1197 (.A(net1200),
    .X(net1197),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1198 (.A(net1200),
    .X(net1198),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1199 (.A(net1200),
    .X(net1199),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1200 (.A(\s0.valid_out[12] [0]),
    .X(net1200),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1201 (.A(net1202),
    .X(net1201),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1202 (.A(net1203),
    .X(net1202),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1203 (.A(net1209),
    .X(net1203),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1204 (.A(net1209),
    .X(net1204),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1205 (.A(net1208),
    .X(net1205),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1206 (.A(net1208),
    .X(net1206),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1207 (.A(net1208),
    .X(net1207),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1208 (.A(net1209),
    .X(net1208),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1209 (.A(\s0.shift_out[13] [0]),
    .X(net1209),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1210 (.A(net1212),
    .X(net1210),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1211 (.A(net1212),
    .X(net1211),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1212 (.A(\s0.valid_out[13] [0]),
    .X(net1212),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1213 (.A(net1215),
    .X(net1213),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1214 (.A(net1215),
    .X(net1214),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1215 (.A(net1216),
    .X(net1215),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1216 (.A(net365),
    .X(net1216),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1217 (.A(net1218),
    .X(net1217),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1218 (.A(net365),
    .X(net1218),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1219 (.A(net1220),
    .X(net1219),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1220 (.A(\s0.valid_out[14] [0]),
    .X(net1220),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1221 (.A(\s0.valid_out[14] [0]),
    .X(net1221),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1222 (.A(\s0.valid_out[14] [0]),
    .X(net1222),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1223 (.A(net1231),
    .X(net1223),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1224 (.A(net1231),
    .X(net1224),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1225 (.A(net1228),
    .X(net1225),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1226 (.A(net1228),
    .X(net1226),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1227 (.A(net1228),
    .X(net1227),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1228 (.A(net1231),
    .X(net1228),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1229 (.A(net1230),
    .X(net1229),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1230 (.A(net1231),
    .X(net1230),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1231 (.A(\s0.shift_out[15] [0]),
    .X(net1231),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1232 (.A(net1233),
    .X(net1232),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1233 (.A(net1235),
    .X(net1233),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1234 (.A(net1235),
    .X(net1234),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1235 (.A(net701),
    .X(net1235),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1236 (.A(net1244),
    .X(net1236),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1237 (.A(net1244),
    .X(net1237),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1238 (.A(net1239),
    .X(net1238),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1239 (.A(net1244),
    .X(net1239),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1240 (.A(net1244),
    .X(net1240),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1241 (.A(net1244),
    .X(net1241),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1242 (.A(net1243),
    .X(net1242),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1243 (.A(net1244),
    .X(net1243),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1244 (.A(net703),
    .X(net1244),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1245 (.A(\s0.valid_out[16] [0]),
    .X(net1245),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1246 (.A(\s0.valid_out[16] [0]),
    .X(net1246),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1247 (.A(net1248),
    .X(net1247),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1248 (.A(\s0.valid_out[16] [0]),
    .X(net1248),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1249 (.A(net1251),
    .X(net1249),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1250 (.A(net1251),
    .X(net1250),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1251 (.A(net498),
    .X(net1251),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1252 (.A(net1256),
    .X(net1252),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1253 (.A(net1256),
    .X(net1253),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1254 (.A(net1256),
    .X(net1254),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1255 (.A(net1256),
    .X(net1255),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1256 (.A(net498),
    .X(net1256),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1257 (.A(net1258),
    .X(net1257),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1258 (.A(\s0.valid_out[17] [0]),
    .X(net1258),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1259 (.A(\s0.valid_out[17] [0]),
    .X(net1259),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1260 (.A(\s0.valid_out[17] [0]),
    .X(net1260),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1261 (.A(net1264),
    .X(net1261),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1262 (.A(net1263),
    .X(net1262),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1263 (.A(net1264),
    .X(net1263),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1264 (.A(\s0.shift_out[18] [0]),
    .X(net1264),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1265 (.A(net1266),
    .X(net1265),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1266 (.A(net472),
    .X(net1266),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1267 (.A(net1268),
    .X(net1267),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1268 (.A(\s0.shift_out[18] [0]),
    .X(net1268),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1269 (.A(net1272),
    .X(net1269),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1270 (.A(net1272),
    .X(net1270),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1271 (.A(net1272),
    .X(net1271),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1272 (.A(\s0.valid_out[18] [0]),
    .X(net1272),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1273 (.A(net1275),
    .X(net1273),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1274 (.A(net1275),
    .X(net1274),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1275 (.A(net1280),
    .X(net1275),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1276 (.A(net1277),
    .X(net1276),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1277 (.A(net1280),
    .X(net1277),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1278 (.A(net1280),
    .X(net1278),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1279 (.A(net1280),
    .X(net1279),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1280 (.A(\s0.shift_out[19] [0]),
    .X(net1280),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1281 (.A(net1285),
    .X(net1281),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1282 (.A(net1285),
    .X(net1282),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1283 (.A(net1285),
    .X(net1283),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1284 (.A(net1285),
    .X(net1284),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1285 (.A(\s0.valid_out[19] [0]),
    .X(net1285),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1286 (.A(net1289),
    .X(net1286),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1287 (.A(net1289),
    .X(net1287),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1288 (.A(net1289),
    .X(net1288),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1289 (.A(\s0.shift_out[20] [0]),
    .X(net1289),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1290 (.A(net1292),
    .X(net1290),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1291 (.A(net1292),
    .X(net1291),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1292 (.A(\s0.shift_out[20] [0]),
    .X(net1292),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1293 (.A(net1295),
    .X(net1293),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1294 (.A(net1295),
    .X(net1294),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1295 (.A(\s0.shift_out[20] [0]),
    .X(net1295),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1296 (.A(net1299),
    .X(net1296),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1297 (.A(net1299),
    .X(net1297),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1298 (.A(net1299),
    .X(net1298),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1299 (.A(\s0.valid_out[20] [0]),
    .X(net1299),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1300 (.A(net1302),
    .X(net1300),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1301 (.A(net1302),
    .X(net1301),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1302 (.A(net347),
    .X(net1302),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1303 (.A(net1304),
    .X(net1303),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1304 (.A(net1306),
    .X(net1304),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1305 (.A(net1306),
    .X(net1305),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1306 (.A(net347),
    .X(net1306),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1307 (.A(net1310),
    .X(net1307),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1308 (.A(net1310),
    .X(net1308),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1309 (.A(net1310),
    .X(net1309),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1310 (.A(net539),
    .X(net1310),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1311 (.A(net1314),
    .X(net1311),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1312 (.A(net1314),
    .X(net1312),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1313 (.A(net1314),
    .X(net1313),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1314 (.A(\s0.shift_out[22] [0]),
    .X(net1314),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1315 (.A(net1317),
    .X(net1315),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1316 (.A(net1317),
    .X(net1316),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1317 (.A(\s0.shift_out[22] [0]),
    .X(net1317),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1318 (.A(net1322),
    .X(net1318),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1319 (.A(net1322),
    .X(net1319),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1320 (.A(net1322),
    .X(net1320),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1321 (.A(net1322),
    .X(net1321),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1322 (.A(\s0.valid_out[22] [0]),
    .X(net1322),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1323 (.A(net1324),
    .X(net1323),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1324 (.A(net398),
    .X(net1324),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1325 (.A(net1326),
    .X(net1325),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1326 (.A(net398),
    .X(net1326),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1327 (.A(\s0.valid_out[23] [0]),
    .X(net1327),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1328 (.A(\s0.valid_out[23] [0]),
    .X(net1328),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1329 (.A(net1333),
    .X(net1329),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1330 (.A(net1333),
    .X(net1330),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1331 (.A(net1333),
    .X(net1331),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1332 (.A(net1333),
    .X(net1332),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1333 (.A(_2983_),
    .X(net1333),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1334 (.A(_2774_),
    .X(net1334),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1335 (.A(_2774_),
    .X(net1335),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1336 (.A(net1338),
    .X(net1336),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1337 (.A(net1338),
    .X(net1337),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1338 (.A(_2743_),
    .X(net1338),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1339 (.A(net1340),
    .X(net1339),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1340 (.A(net1343),
    .X(net1340),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1341 (.A(net1343),
    .X(net1341),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1342 (.A(net1343),
    .X(net1342),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1343 (.A(net1351),
    .X(net1343),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1344 (.A(net1351),
    .X(net1344),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1345 (.A(net1351),
    .X(net1345),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1346 (.A(net1350),
    .X(net1346),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1347 (.A(net1350),
    .X(net1347),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1348 (.A(net1350),
    .X(net1348),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1349 (.A(net1350),
    .X(net1349),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1350 (.A(net1351),
    .X(net1350),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1351 (.A(net1389),
    .X(net1351),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1352 (.A(net1354),
    .X(net1352),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1353 (.A(net1354),
    .X(net1353),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1354 (.A(net1357),
    .X(net1354),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1355 (.A(net1356),
    .X(net1355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1356 (.A(net1357),
    .X(net1356),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1357 (.A(net1364),
    .X(net1357),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1358 (.A(net1362),
    .X(net1358),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1359 (.A(net1362),
    .X(net1359),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1360 (.A(net1362),
    .X(net1360),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1361 (.A(net1362),
    .X(net1361),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1362 (.A(net1364),
    .X(net1362),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1363 (.A(net1364),
    .X(net1363),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1364 (.A(net1389),
    .X(net1364),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1365 (.A(net1377),
    .X(net1365),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1366 (.A(net1377),
    .X(net1366),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1367 (.A(net1369),
    .X(net1367),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1368 (.A(net1369),
    .X(net1368),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1369 (.A(net1377),
    .X(net1369),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1370 (.A(net1373),
    .X(net1370),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1371 (.A(net1373),
    .X(net1371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1372 (.A(net1373),
    .X(net1372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1373 (.A(net1377),
    .X(net1373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1374 (.A(net1376),
    .X(net1374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1375 (.A(net1376),
    .X(net1375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1376 (.A(net1377),
    .X(net1376),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1377 (.A(net1389),
    .X(net1377),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1378 (.A(net1383),
    .X(net1378),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1379 (.A(net1383),
    .X(net1379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1380 (.A(net1383),
    .X(net1380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1381 (.A(net1383),
    .X(net1381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1382 (.A(net1383),
    .X(net1382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1383 (.A(net1389),
    .X(net1383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1384 (.A(net1388),
    .X(net1384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1385 (.A(net1388),
    .X(net1385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1386 (.A(net1388),
    .X(net1386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1387 (.A(net1388),
    .X(net1387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1388 (.A(net1389),
    .X(net1388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1389 (.A(_2742_),
    .X(net1389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1390 (.A(uio_in[1]),
    .X(net1390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1391 (.A(uio_in[1]),
    .X(net1391),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1392 (.A(net1393),
    .X(net1392),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1393 (.A(net1397),
    .X(net1393),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1394 (.A(net1396),
    .X(net1394),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1395 (.A(net1396),
    .X(net1395),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1396 (.A(net1397),
    .X(net1396),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1397 (.A(uio_in[0]),
    .X(net1397),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1398 (.A(net1401),
    .X(net1398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1399 (.A(net1401),
    .X(net1399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1400 (.A(net1401),
    .X(net1400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1401 (.A(ui_in[7]),
    .X(net1401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1402 (.A(net1406),
    .X(net1402),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1403 (.A(net1406),
    .X(net1403),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1404 (.A(net1406),
    .X(net1404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1405 (.A(net1406),
    .X(net1405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1406 (.A(ui_in[7]),
    .X(net1406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1407 (.A(net1410),
    .X(net1407),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1408 (.A(net1410),
    .X(net1408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1409 (.A(net1410),
    .X(net1409),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1410 (.A(ui_in[6]),
    .X(net1410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1411 (.A(net1415),
    .X(net1411),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1412 (.A(net1415),
    .X(net1412),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1413 (.A(net1415),
    .X(net1413),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1414 (.A(net1415),
    .X(net1414),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1415 (.A(ui_in[6]),
    .X(net1415),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1416 (.A(net1420),
    .X(net1416),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1417 (.A(net1420),
    .X(net1417),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1418 (.A(net1420),
    .X(net1418),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1419 (.A(net1420),
    .X(net1419),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1420 (.A(ui_in[5]),
    .X(net1420),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1421 (.A(net1425),
    .X(net1421),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1422 (.A(net1425),
    .X(net1422),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1423 (.A(net1425),
    .X(net1423),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1424 (.A(net1425),
    .X(net1424),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1425 (.A(ui_in[5]),
    .X(net1425),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1426 (.A(net1429),
    .X(net1426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1427 (.A(net1429),
    .X(net1427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1428 (.A(net1429),
    .X(net1428),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1429 (.A(ui_in[4]),
    .X(net1429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1430 (.A(net1434),
    .X(net1430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1431 (.A(net1434),
    .X(net1431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1432 (.A(net1434),
    .X(net1432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1433 (.A(net1434),
    .X(net1433),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1434 (.A(ui_in[4]),
    .X(net1434),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1435 (.A(net1438),
    .X(net1435),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1436 (.A(net1438),
    .X(net1436),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1437 (.A(net1438),
    .X(net1437),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1438 (.A(ui_in[3]),
    .X(net1438),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1439 (.A(net1442),
    .X(net1439),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1440 (.A(net1441),
    .X(net1440),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1441 (.A(net1442),
    .X(net1441),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1442 (.A(ui_in[3]),
    .X(net1442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1443 (.A(net1448),
    .X(net1443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1444 (.A(net1448),
    .X(net1444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1445 (.A(net1446),
    .X(net1445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1446 (.A(net1448),
    .X(net1446),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1447 (.A(net1448),
    .X(net1447),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1448 (.A(ui_in[2]),
    .X(net1448),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1449 (.A(net1451),
    .X(net1449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1450 (.A(net1451),
    .X(net1450),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1451 (.A(net1457),
    .X(net1451),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1452 (.A(net1457),
    .X(net1452),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1453 (.A(net1457),
    .X(net1453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1454 (.A(net1456),
    .X(net1454),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1455 (.A(net1456),
    .X(net1455),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1456 (.A(net1457),
    .X(net1456),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1457 (.A(ui_in[1]),
    .X(net1457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1458 (.A(net1461),
    .X(net1458),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1459 (.A(net1460),
    .X(net1459),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1460 (.A(net1461),
    .X(net1460),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1461 (.A(ui_in[0]),
    .X(net1461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1462 (.A(net1463),
    .X(net1462),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1463 (.A(net1476),
    .X(net1463),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1464 (.A(net1465),
    .X(net1464),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1465 (.A(net1469),
    .X(net1465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1466 (.A(net1467),
    .X(net1466),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1467 (.A(net1469),
    .X(net1467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1468 (.A(net1469),
    .X(net1468),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1469 (.A(net1476),
    .X(net1469),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1470 (.A(net1472),
    .X(net1470),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1471 (.A(net1472),
    .X(net1471),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1472 (.A(net1476),
    .X(net1472),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1473 (.A(net1475),
    .X(net1473),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1474 (.A(net1475),
    .X(net1474),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1475 (.A(net1476),
    .X(net1475),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1476 (.A(net1493),
    .X(net1476),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1477 (.A(net1483),
    .X(net1477),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1478 (.A(net1483),
    .X(net1478),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1479 (.A(net1482),
    .X(net1479),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1480 (.A(net1482),
    .X(net1480),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1481 (.A(net1482),
    .X(net1481),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1482 (.A(net1483),
    .X(net1482),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1483 (.A(net1493),
    .X(net1483),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1484 (.A(net1487),
    .X(net1484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1485 (.A(net1487),
    .X(net1485),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1486 (.A(net1487),
    .X(net1486),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1487 (.A(net1493),
    .X(net1487),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1488 (.A(net1492),
    .X(net1488),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1489 (.A(net1492),
    .X(net1489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1490 (.A(net1492),
    .X(net1490),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1491 (.A(net1492),
    .X(net1491),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1492 (.A(net1493),
    .X(net1492),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1493 (.A(rst_n),
    .X(net1493),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output1 (.A(net1),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_top_sorter_10 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net10));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_14_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_25_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload0 (.A(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload1 (.VDD(VPWR),
    .A(clknet_leaf_4_clk),
    .VSS(VGND));
 sg13g2_buf_8 clkload2 (.A(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload3 (.VDD(VPWR),
    .A(clknet_leaf_6_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload4 (.VDD(VPWR),
    .A(clknet_leaf_14_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload7 (.VDD(VPWR),
    .A(clknet_leaf_16_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload8 (.VDD(VPWR),
    .A(clknet_leaf_26_clk),
    .VSS(VGND));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\s0.genblk1[4].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold2 (.A(\s0.genblk1[17].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold3 (.A(\s0.genblk1[15].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold4 (.A(\s0.genblk1[8].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold5 (.A(\s0.genblk1[1].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold6 (.A(\s0.genblk1[16].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold7 (.A(\s0.genblk1[19].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold8 (.A(\s0.genblk1[14].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold9 (.A(\s0.genblk1[10].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold10 (.A(\s0.genblk1[22].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold11 (.A(\s0.genblk1[5].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold12 (.A(\s0.genblk1[21].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold13 (.A(\s0.module0.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold14 (.A(\s0.genblk1[2].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold15 (.A(\s0.genblk1[23].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold16 (.A(\s0.genblk1[9].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold17 (.A(\s0.genblk1[18].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold18 (.A(\s0.genblk1[20].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold19 (.A(\s0.genblk1[6].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold20 (.A(\s0.genblk1[3].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold21 (.A(\s0.genblk1[11].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold22 (.A(\s0.genblk1[12].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold23 (.A(\s0.genblk1[13].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold24 (.A(\s0.genblk1[7].modules.bubble ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold25 (.A(\s0.was_valid_out[5] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0224_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold27 (.A(\s0.shift_out[21] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold28 (.A(\s0.was_valid_out[12] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0133_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold30 (.A(\s0.was_valid_out[10] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0157_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold32 (.A(\s0.data_out[19][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0517_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold34 (.A(\s0.data_out[23][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold35 (.A(_2932_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold36 (.A(\s0.was_valid_out[2] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0260_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold38 (.A(\s0.was_valid_out[8] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0188_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold40 (.A(\s0.shift_out[10] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold41 (.A(\s0.data_out[0][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold42 (.A(\s0.was_valid_out[15] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0097_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold44 (.A(\s0.was_valid_out[6] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold45 (.A(\s0.shift_out[14] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold46 (.A(\s0.was_valid_out[19] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0049_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold48 (.A(\s0.data_out[17][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0734_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold50 (.A(\s0.was_valid_out[16] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold51 (.A(\s0.data_out[8][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold52 (.A(_1731_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold53 (.A(\s0.data_out[11][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold54 (.A(_1515_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold55 (.A(\s0.data_out[0][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0289_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold57 (.A(\s0.data_out[22][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold58 (.A(_3057_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold59 (.A(\s0.data_out[23][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold61 (.A(\s0.data_out[23][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold63 (.A(\s0.was_valid_out[17] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold64 (.A(\s0.shift_out[5] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold65 (.A(\s0.data_out[0][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold66 (.A(\s0.data_out[0][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold67 (.A(\s0.data_out[3][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold68 (.A(_2426_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold69 (.A(\s0.data_out[6][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold70 (.A(_1939_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold71 (.A(\s0.shift_out[12] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold72 (.A(\s0.was_valid_out[22] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0013_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold74 (.A(\s0.data_out[0][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold75 (.A(\s0.data_out[0][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold76 (.A(\s0.valid_out[2] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold77 (.A(\s0.shift_out[0] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold78 (.A(\s0.shift_out[23] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold79 (.A(_2995_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold80 (.A(\s0.data_out[3][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0253_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold82 (.A(\s0.data_out[0][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0291_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold84 (.A(\s0.data_out[6][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold85 (.A(_2061_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold86 (.A(\s0.data_out[13][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0132_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold88 (.A(\s0.data_out[7][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0205_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold90 (.A(\s0.data_out[18][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0068_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold92 (.A(\s0.data_out[23][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold94 (.A(\s0.data_out[12][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold95 (.A(_1288_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold96 (.A(\s0.data_out[23][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0009_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold98 (.A(\s0.data_out[18][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0066_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold100 (.A(\s0.data_out[15][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0103_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold102 (.A(\s0.data_out[11][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0151_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold104 (.A(\s0.data_out[20][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold106 (.A(\s0.data_out[16][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold107 (.A(\s0.was_valid_out[0] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold108 (.A(\s0.data_out[18][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0067_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold110 (.A(\s0.data_out[15][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0106_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold112 (.A(\s0.data_out[20][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0047_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold114 (.A(\s0.data_out[3][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0254_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold116 (.A(\s0.data_out[18][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0653_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold118 (.A(\s0.data_out[23][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0012_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold120 (.A(\s0.data_out[18][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0069_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold122 (.A(\s0.data_out[12][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0137_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold124 (.A(\s0.data_out[4][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0243_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold126 (.A(\s0.shift_out[6] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold127 (.A(_2109_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0219_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold129 (.A(\s0.data_out[5][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0234_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold131 (.A(\s0.data_out[11][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0156_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold133 (.A(\s0.data_out[7][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0206_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold135 (.A(\s0.data_out[23][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold137 (.A(\s0.data_out[13][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0127_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold139 (.A(\s0.data_out[23][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0010_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold141 (.A(\s0.data_out[11][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0152_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold143 (.A(\s0.data_out[2][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0267_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold145 (.A(\s0.data_out[9][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0182_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold147 (.A(\s0.data_out[12][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold148 (.A(\s0.data_out[20][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0046_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold150 (.A(\s0.data_out[7][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0209_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold152 (.A(\s0.shift_out[18] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold153 (.A(\s0.data_out[20][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0048_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold155 (.A(\s0.data_out[16][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0094_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold157 (.A(\s0.data_out[10][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0171_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold159 (.A(\s0.data_out[16][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0090_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold161 (.A(\s0.data_out[13][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold162 (.A(\s0.data_out[16][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0092_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold164 (.A(\s0.data_out[3][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0259_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold166 (.A(\s0.data_out[19][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0057_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold168 (.A(\s0.data_out[5][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold169 (.A(\s0.data_out[10][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0169_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold171 (.A(\s0.data_out[13][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold172 (.A(\s0.data_out[4][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0247_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold174 (.A(\s0.data_out[1][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0277_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold176 (.A(\s0.data_out[20][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0045_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold178 (.A(\s0.shift_out[17] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold179 (.A(\s0.data_out[18][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0072_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold181 (.A(\s0.data_out[6][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0217_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold183 (.A(\s0.data_out[16][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0096_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold185 (.A(\s0.data_out[9][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold186 (.A(\s0.data_out[19][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold187 (.A(\s0.data_out[4][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0246_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold189 (.A(\s0.data_out[9][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0186_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold191 (.A(\s0.data_out[17][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold192 (.A(\s0.data_out[2][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0271_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold194 (.A(\s0.data_out[2][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0265_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold196 (.A(\s0.was_valid_out[1] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0272_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold198 (.A(\s0.data_out[8][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold199 (.A(\s0.data_out[21][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0032_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold201 (.A(\s0.data_out[7][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold202 (.A(\s0.data_out[14][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold203 (.A(_1206_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold204 (.A(\s0.was_valid_out[3] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold205 (.A(\s0.data_out[16][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0093_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold207 (.A(\s0.data_out[21][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0324_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold209 (.A(\s0.data_out[17][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold210 (.A(\s0.data_out[15][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0102_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold212 (.A(\s0.data_out[13][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0128_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold214 (.A(\s0.data_out[18][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0769_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold216 (.A(\s0.data_out[10][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold217 (.A(\s0.data_out[8][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1878_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold219 (.A(\s0.valid_out[21] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold220 (.A(\s0.data_out[3][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold221 (.A(\s0.data_out[1][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold222 (.A(_2668_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold223 (.A(\s0.was_valid_out[18] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0061_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold225 (.A(\s0.data_out[14][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0119_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold227 (.A(\s0.data_out[0][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold228 (.A(\s0.data_out[14][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold229 (.A(\s0.data_out[5][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold230 (.A(\s0.data_out[13][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold231 (.A(_1325_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold232 (.A(\s0.was_valid_out[7] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold233 (.A(\s0.data_out[15][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0104_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold235 (.A(\s0.data_out[7][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold236 (.A(_1899_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold237 (.A(\s0.data_out[21][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0030_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold239 (.A(\s0.was_valid_out[23] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold240 (.A(\s0.data_out[17][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold241 (.A(\s0.data_out[15][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0108_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold243 (.A(\s0.shift_out[7] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold244 (.A(\s0.data_out[22][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0319_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold246 (.A(\s0.was_valid_out[13] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0121_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold248 (.A(\s0.data_out[5][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold249 (.A(\s0.data_out[4][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold250 (.A(\s0.data_out[5][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold251 (.A(\s0.data_out[5][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold252 (.A(\s0.data_out[9][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0181_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold254 (.A(\s0.data_out[3][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0255_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold256 (.A(\s0.data_out[2][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold257 (.A(_2567_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold258 (.A(\s0.data_out[6][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold259 (.A(\s0.data_out[1][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold260 (.A(\s0.data_out[2][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0270_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold262 (.A(\s0.data_out[2][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold263 (.A(\s0.data_out[2][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold264 (.A(_2563_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold265 (.A(\s0.shift_out[3] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold266 (.A(\s0.data_out[22][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold268 (.A(\s0.data_out[11][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold269 (.A(\s0.data_out[9][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0183_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold271 (.A(\s0.data_out[14][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold272 (.A(_1193_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold273 (.A(\s0.data_out[22][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0023_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold275 (.A(\s0.data_out[12][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold276 (.A(\s0.data_out[9][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold277 (.A(\s0.data_out[19][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0639_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold279 (.A(\s0.data_out[16][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold280 (.A(\s0.data_out[4][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold281 (.A(\s0.data_out[3][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold282 (.A(\s0.data_out[14][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold283 (.A(\s0.data_out[22][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0017_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold285 (.A(\s0.data_out[1][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold286 (.A(\s0.data_out[5][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold287 (.A(\s0.data_out[15][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold288 (.A(\s0.shift_out[4] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold289 (.A(\s0.data_out[21][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold290 (.A(\s0.data_out[10][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold291 (.A(_1543_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold292 (.A(\s0.data_out[14][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold293 (.A(\s0.data_out[10][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold294 (.A(_1670_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold295 (.A(\s0.was_valid_out[14] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold296 (.A(\s0.data_out[12][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold297 (.A(_1438_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold298 (.A(\s0.data_out[11][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold299 (.A(\s0.data_out[12][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0142_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold301 (.A(\s0.data_out[12][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold302 (.A(\s0.data_out[19][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0658_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold304 (.A(\s0.data_out[21][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold305 (.A(\s0.data_out[1][7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold306 (.A(\s0.data_out[10][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold307 (.A(\s0.data_out[7][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold308 (.A(\s0.data_out[20][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0044_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold310 (.A(\s0.data_out[6][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold311 (.A(\s0.data_out[12][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold312 (.A(\s0.data_out[7][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold313 (.A(\s0.data_out[20][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0042_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold315 (.A(\s0.data_out[22][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold316 (.A(\s0.data_out[10][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold317 (.A(\s0.data_out[8][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0195_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold319 (.A(\s0.data_out[7][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold320 (.A(\s0.data_out[22][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold322 (.A(\s0.data_out[4][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold323 (.A(\s0.data_out[15][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold324 (.A(\s0.was_valid_out[11] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0144_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold326 (.A(\s0.data_out[22][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold327 (.A(\s0.data_out[14][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold328 (.A(\s0.data_out[21][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold329 (.A(\s0.was_valid_out[20] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold330 (.A(\s0.data_out[21][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold331 (.A(\s0.data_out[12][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold332 (.A(\s0.data_out[1][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold333 (.A(\s0.data_out[17][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold334 (.A(\s0.data_out[8][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold335 (.A(_1897_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold336 (.A(\s0.data_out[5][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold337 (.A(\s0.data_out[19][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0055_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold339 (.A(\s0.data_out[21][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold340 (.A(\s0.data_out[18][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold341 (.A(\s0.data_out[11][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold342 (.A(\s0.data_out[16][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold343 (.A(\s0.data_out[2][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold344 (.A(\s0.data_out[17][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0880_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold346 (.A(\s0.was_valid_out[9] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0176_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold348 (.A(\s0.data_out[17][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold349 (.A(\s0.data_out[6][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold350 (.A(\s0.data_out[8][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0196_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold352 (.A(\s0.data_out[20][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold353 (.A(\s0.data_out[8][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold354 (.A(\s0.data_out[10][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold355 (.A(\s0.data_out[9][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold356 (.A(\s0.data_out[4][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold357 (.A(\s0.data_out[1][4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold358 (.A(\s0.data_out[3][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold359 (.A(\s0.data_out[13][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold360 (.A(\s0.data_out[9][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold361 (.A(\s0.data_out[4][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold362 (.A(\s0.data_out[6][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold363 (.A(\s0.data_out[1][2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold364 (.A(\s0.data_out[14][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold365 (.A(_1210_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold366 (.A(\s0.data_out[13][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold367 (.A(\s0.data_out[8][5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0197_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold369 (.A(\s0.data_out[17][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold370 (.A(\s0.data_out[19][3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0056_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold372 (.A(\s0.data_out[6][0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold373 (.A(\s0.data_out[15][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold374 (.A(_1102_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold375 (.A(\s0.data_out[19][1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0054_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold377 (.A(\s0.data_out[11][6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold378 (.A(\s0.was_valid_out[21] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold379 (.A(\s0.was_valid_out[4] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold380 (.A(\s0.data_new_delayed[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold381 (.A(\s0.valid_out[15] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold382 (.A(\s0.data_new_delayed[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold383 (.A(\s0.shift_out[16] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold384 (.A(\s0.data_new_delayed[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold385 (.A(\s0.data_new_delayed[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold386 (.A(\s0.valid_out[4] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold387 (.A(\s0.data_new_delayed[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold388 (.A(\s0.data_new_delayed[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold389 (.A(\s0.data_new_delayed[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold390 (.A(\s0.shift_out[1] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold391 (.A(\s0.valid_out[5] [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold392 (.A(\s0.data_new_delayed[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net712));
 sg13g2_decap_8 FILLER_0_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net10;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net319;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net320;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
endmodule
