module heichips25_template (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net36;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire \sap_3_inst.alu.clk_regs ;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire clk_div_out;
 wire mem_mar_we;
 wire mem_ram_we;
 wire regFile_serial;
 wire regFile_serial_start;
 wire \sap_3_inst.alu.acc[0] ;
 wire \sap_3_inst.alu.acc[1] ;
 wire \sap_3_inst.alu.acc[2] ;
 wire \sap_3_inst.alu.acc[3] ;
 wire \sap_3_inst.alu.acc[4] ;
 wire \sap_3_inst.alu.acc[5] ;
 wire \sap_3_inst.alu.acc[6] ;
 wire \sap_3_inst.alu.acc[7] ;
 wire \sap_3_inst.alu.act[0] ;
 wire \sap_3_inst.alu.act[1] ;
 wire \sap_3_inst.alu.act[2] ;
 wire \sap_3_inst.alu.act[3] ;
 wire \sap_3_inst.alu.act[4] ;
 wire \sap_3_inst.alu.act[5] ;
 wire \sap_3_inst.alu.act[6] ;
 wire \sap_3_inst.alu.act[7] ;
 wire \sap_3_inst.alu.carry ;
 wire \sap_3_inst.alu.clk ;
 wire \sap_3_inst.alu.flags[0] ;
 wire \sap_3_inst.alu.flags[1] ;
 wire \sap_3_inst.alu.flags[2] ;
 wire \sap_3_inst.alu.flags[3] ;
 wire \sap_3_inst.alu.flags[4] ;
 wire \sap_3_inst.alu.flags[5] ;
 wire \sap_3_inst.alu.flags[6] ;
 wire \sap_3_inst.alu.flags[7] ;
 wire \sap_3_inst.alu.tmp[0] ;
 wire \sap_3_inst.alu.tmp[1] ;
 wire \sap_3_inst.alu.tmp[2] ;
 wire \sap_3_inst.alu.tmp[3] ;
 wire \sap_3_inst.alu.tmp[4] ;
 wire \sap_3_inst.alu.tmp[5] ;
 wire \sap_3_inst.alu.tmp[6] ;
 wire \sap_3_inst.alu.tmp[7] ;
 wire \sap_3_inst.controller.opcode[0] ;
 wire \sap_3_inst.controller.opcode[1] ;
 wire \sap_3_inst.controller.opcode[2] ;
 wire \sap_3_inst.controller.opcode[3] ;
 wire \sap_3_inst.controller.opcode[4] ;
 wire \sap_3_inst.controller.opcode[5] ;
 wire \sap_3_inst.controller.opcode[6] ;
 wire \sap_3_inst.controller.opcode[7] ;
 wire \sap_3_inst.controller.stage[0] ;
 wire \sap_3_inst.controller.stage[1] ;
 wire \sap_3_inst.controller.stage[2] ;
 wire \sap_3_inst.controller.stage[3] ;
 wire \sap_3_inst.out[0] ;
 wire \sap_3_inst.out[1] ;
 wire \sap_3_inst.out[2] ;
 wire \sap_3_inst.out[3] ;
 wire \sap_3_inst.out[4] ;
 wire \sap_3_inst.out[5] ;
 wire \sap_3_inst.out[6] ;
 wire \sap_3_inst.out[7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.bit_pos[0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[0][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[10][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[11][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[1][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[2][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[3][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[4][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[5][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[6][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[7][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[8][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.data[9][7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[3] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[4] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[5] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[6] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.shadow_reg[7] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.state[0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.state[1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.word_index[0] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.word_index[1] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.word_index[2] ;
 wire \sap_3_inst.reg_file.array_serializer_inst.word_index[3] ;
 wire sap_3_outputReg_serial;
 wire sap_3_outputReg_start_sync;
 wire \u_ser.bit_pos[0] ;
 wire \u_ser.bit_pos[1] ;
 wire \u_ser.bit_pos[2] ;
 wire \u_ser.shadow_reg[0] ;
 wire \u_ser.shadow_reg[1] ;
 wire \u_ser.shadow_reg[2] ;
 wire \u_ser.shadow_reg[3] ;
 wire \u_ser.shadow_reg[4] ;
 wire \u_ser.shadow_reg[5] ;
 wire \u_ser.shadow_reg[6] ;
 wire \u_ser.shadow_reg[7] ;
 wire \u_ser.state[0] ;
 wire \u_ser.state[1] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net34;
 wire net35;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net31;
 wire net32;
 wire net33;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_0_clk_div_out;
 wire clknet_1_0__leaf_clk_div_out;
 wire clknet_1_1__leaf_clk_div_out;
 wire \clknet_leaf_0_sap_3_inst.alu.clk ;
 wire \clknet_leaf_1_sap_3_inst.alu.clk ;
 wire \clknet_leaf_2_sap_3_inst.alu.clk ;
 wire \clknet_leaf_3_sap_3_inst.alu.clk ;
 wire \clknet_0_sap_3_inst.alu.clk ;
 wire \clknet_1_0__leaf_sap_3_inst.alu.clk ;
 wire \clknet_1_1__leaf_sap_3_inst.alu.clk ;
 wire \clknet_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_0_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_1_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_2_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_3_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_4_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_5_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_6_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_7_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_8_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_9_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_10_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_11_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_12_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_13_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_14_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_4_15_0_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_0__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_1__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_2__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_3__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_4__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_5__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_6__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_7__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_8__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_9__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_10__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_11__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_12__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_13__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_14__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_15__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_16__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_17__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_18__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_19__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_20__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_21__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_22__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_23__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_24__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_25__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_26__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_27__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_28__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_29__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_30__leaf_sap_3_inst.alu.clk_regs ;
 wire \clknet_5_31__leaf_sap_3_inst.alu.clk_regs ;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;

 sg13g2_inv_1 _2009_ (.Y(_1432_),
    .A(\u_ser.state[0] ));
 sg13g2_inv_1 _2010_ (.Y(_1433_),
    .A(\u_ser.state[1] ));
 sg13g2_inv_1 _2011_ (.Y(_1434_),
    .A(\u_ser.bit_pos[2] ));
 sg13g2_inv_1 _2012_ (.Y(_1435_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ));
 sg13g2_inv_4 _2013_ (.A(net738),
    .Y(_1436_));
 sg13g2_inv_2 _2014_ (.Y(_1437_),
    .A(net732));
 sg13g2_inv_2 _2015_ (.Y(_1438_),
    .A(net729));
 sg13g2_inv_1 _2016_ (.Y(_1439_),
    .A(net725));
 sg13g2_inv_2 _2017_ (.Y(_1440_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][3] ));
 sg13g2_inv_1 _2018_ (.Y(_1441_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ));
 sg13g2_inv_1 _2019_ (.Y(_1442_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ));
 sg13g2_inv_1 _2020_ (.Y(_1443_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ));
 sg13g2_inv_1 _2021_ (.Y(_1444_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][2] ));
 sg13g2_inv_1 _2022_ (.Y(_1445_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ));
 sg13g2_inv_1 _2023_ (.Y(_1446_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ));
 sg13g2_inv_1 _2024_ (.Y(_1447_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ));
 sg13g2_inv_1 _2025_ (.Y(_1448_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ));
 sg13g2_inv_1 _2026_ (.Y(_1449_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ));
 sg13g2_inv_1 _2027_ (.Y(_1450_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ));
 sg13g2_inv_1 _2028_ (.Y(_1451_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ));
 sg13g2_inv_2 _2029_ (.Y(_1452_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ));
 sg13g2_inv_1 _2030_ (.Y(_1453_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ));
 sg13g2_inv_2 _2031_ (.Y(_1454_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ));
 sg13g2_inv_2 _2032_ (.Y(_1455_),
    .A(net757));
 sg13g2_inv_1 _2033_ (.Y(_1456_),
    .A(net760));
 sg13g2_inv_2 _2034_ (.Y(_1457_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][1] ));
 sg13g2_inv_1 _2035_ (.Y(_1458_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ));
 sg13g2_inv_1 _2036_ (.Y(_1459_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ));
 sg13g2_inv_2 _2037_ (.Y(_1460_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][0] ));
 sg13g2_inv_1 _2038_ (.Y(_1461_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ));
 sg13g2_inv_1 _2039_ (.Y(_1462_),
    .A(\sap_3_inst.alu.act[0] ));
 sg13g2_inv_2 _2040_ (.Y(_1463_),
    .A(\sap_3_inst.alu.tmp[1] ));
 sg13g2_inv_1 _2041_ (.Y(_1464_),
    .A(\sap_3_inst.alu.tmp[2] ));
 sg13g2_inv_1 _2042_ (.Y(_1465_),
    .A(\sap_3_inst.alu.tmp[3] ));
 sg13g2_inv_1 _2043_ (.Y(_1466_),
    .A(\sap_3_inst.alu.tmp[5] ));
 sg13g2_inv_1 _2044_ (.Y(_1467_),
    .A(\sap_3_inst.alu.tmp[6] ));
 sg13g2_inv_2 _2045_ (.Y(_1468_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][4] ));
 sg13g2_inv_1 _2046_ (.Y(_1469_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ));
 sg13g2_inv_1 _2047_ (.Y(_1470_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ));
 sg13g2_inv_1 _2048_ (.Y(_1471_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ));
 sg13g2_inv_1 _2049_ (.Y(_1472_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ));
 sg13g2_inv_1 _2050_ (.Y(_1473_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ));
 sg13g2_inv_1 _2051_ (.Y(_1474_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ));
 sg13g2_inv_2 _2052_ (.Y(_1475_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][5] ));
 sg13g2_inv_1 _2053_ (.Y(_1476_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ));
 sg13g2_inv_1 _2054_ (.Y(_1477_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ));
 sg13g2_inv_1 _2055_ (.Y(_1478_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ));
 sg13g2_inv_2 _2056_ (.Y(_1479_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][6] ));
 sg13g2_inv_1 _2057_ (.Y(_1480_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ));
 sg13g2_inv_1 _2058_ (.Y(_1481_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ));
 sg13g2_inv_1 _2059_ (.Y(_1482_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ));
 sg13g2_inv_1 _2060_ (.Y(_1483_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ));
 sg13g2_inv_1 _2061_ (.Y(_1484_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ));
 sg13g2_inv_1 _2062_ (.Y(_1485_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ));
 sg13g2_inv_1 _2063_ (.Y(_1486_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ));
 sg13g2_inv_1 _2064_ (.Y(_1487_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ));
 sg13g2_inv_1 _2065_ (.Y(_1488_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ));
 sg13g2_inv_1 _2066_ (.Y(_1489_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ));
 sg13g2_inv_2 _2067_ (.Y(_1490_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][7] ));
 sg13g2_inv_1 _2068_ (.Y(_1491_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ));
 sg13g2_inv_1 _2069_ (.Y(_1492_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ));
 sg13g2_inv_1 _2070_ (.Y(_1493_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ));
 sg13g2_inv_1 _2071_ (.Y(_1494_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ));
 sg13g2_inv_1 _2072_ (.Y(_1495_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ));
 sg13g2_inv_1 _2073_ (.Y(_1496_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ));
 sg13g2_inv_4 _2074_ (.A(net82),
    .Y(_1497_));
 sg13g2_inv_1 _2075_ (.Y(_1498_),
    .A(net768));
 sg13g2_inv_1 _2077__2 (.Y(net36),
    .A(\clknet_leaf_2_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4025__3 (.Y(net37),
    .A(\clknet_leaf_2_sap_3_inst.alu.clk ));
 sg13g2_nor2_2 _2078_ (.A(net717),
    .B(net716),
    .Y(_1499_));
 sg13g2_or2_1 _2079_ (.X(_1500_),
    .B(net716),
    .A(net717));
 sg13g2_nor2_1 _2080_ (.A(net719),
    .B(net718),
    .Y(_1501_));
 sg13g2_nor2_1 _2081_ (.A(net718),
    .B(_1500_),
    .Y(_1502_));
 sg13g2_nand2_1 _2082_ (.Y(_1503_),
    .A(_1499_),
    .B(net715));
 sg13g2_and2_1 _2083_ (.A(net731),
    .B(net729),
    .X(_1504_));
 sg13g2_nand2_1 _2084_ (.Y(_1505_),
    .A(\sap_3_inst.controller.opcode[4] ),
    .B(net730));
 sg13g2_nor2b_2 _2085_ (.A(net742),
    .B_N(net739),
    .Y(_1506_));
 sg13g2_nand2b_2 _2086_ (.Y(_1507_),
    .B(net739),
    .A_N(net742));
 sg13g2_nor2_2 _2087_ (.A(_1436_),
    .B(_1507_),
    .Y(_1508_));
 sg13g2_nand3b_1 _2088_ (.B(net737),
    .C(net740),
    .Y(_1509_),
    .A_N(net742));
 sg13g2_nor2b_2 _2089_ (.A(net725),
    .B_N(net727),
    .Y(_1510_));
 sg13g2_nand2b_2 _2090_ (.Y(_1511_),
    .B(net727),
    .A_N(net725));
 sg13g2_nor2_1 _2091_ (.A(_1509_),
    .B(_1511_),
    .Y(_1512_));
 sg13g2_nand2_1 _2092_ (.Y(_1513_),
    .A(_1508_),
    .B(_1510_));
 sg13g2_nor3_2 _2093_ (.A(net736),
    .B(net724),
    .C(_1511_),
    .Y(_1514_));
 sg13g2_nand3b_1 _2094_ (.B(_1504_),
    .C(_1510_),
    .Y(_1515_),
    .A_N(net733));
 sg13g2_nor2_1 _2095_ (.A(net740),
    .B(net741),
    .Y(_1516_));
 sg13g2_or2_1 _2096_ (.X(_1517_),
    .B(net741),
    .A(net739));
 sg13g2_nor2_2 _2097_ (.A(\sap_3_inst.controller.opcode[4] ),
    .B(net730),
    .Y(_1518_));
 sg13g2_or2_1 _2098_ (.X(_1519_),
    .B(net729),
    .A(net732));
 sg13g2_nor2_2 _2099_ (.A(net726),
    .B(net727),
    .Y(_1520_));
 sg13g2_or2_1 _2100_ (.X(_1521_),
    .B(net728),
    .A(net726));
 sg13g2_nor2_2 _2101_ (.A(net735),
    .B(net737),
    .Y(_1522_));
 sg13g2_nor3_1 _2102_ (.A(net738),
    .B(net725),
    .C(net727),
    .Y(_1523_));
 sg13g2_or3_1 _2103_ (.A(net738),
    .B(net725),
    .C(net727),
    .X(_1524_));
 sg13g2_nand4_1 _2104_ (.B(_1518_),
    .C(_1520_),
    .A(_1516_),
    .Y(_1525_),
    .D(_1522_));
 sg13g2_o21ai_1 _2105_ (.B1(_1525_),
    .Y(_1526_),
    .A1(_1509_),
    .A2(_1515_));
 sg13g2_and2_1 _2106_ (.A(net719),
    .B(net718),
    .X(_1527_));
 sg13g2_nand2_2 _2107_ (.Y(_1528_),
    .A(net719),
    .B(\sap_3_inst.controller.stage[1] ));
 sg13g2_nor2_1 _2108_ (.A(_1500_),
    .B(_1528_),
    .Y(_1529_));
 sg13g2_nand2_2 _2109_ (.Y(_1530_),
    .A(_1499_),
    .B(_1527_));
 sg13g2_nor2b_2 _2110_ (.A(net718),
    .B_N(net719),
    .Y(_1531_));
 sg13g2_nand2_1 _2111_ (.Y(_1532_),
    .A(_1499_),
    .B(_1531_));
 sg13g2_nor2b_2 _2112_ (.A(\sap_3_inst.controller.stage[0] ),
    .B_N(net718),
    .Y(_1533_));
 sg13g2_nand2_1 _2113_ (.Y(_1534_),
    .A(_1499_),
    .B(_1533_));
 sg13g2_xnor2_1 _2114_ (.Y(_1535_),
    .A(net719),
    .B(net718));
 sg13g2_xor2_1 _2115_ (.B(\sap_3_inst.controller.stage[1] ),
    .A(net719),
    .X(_1536_));
 sg13g2_a221oi_1 _2116_ (.B2(_1499_),
    .C1(_1526_),
    .B1(_1536_),
    .A1(net713),
    .Y(_1537_),
    .A2(net694));
 sg13g2_nand2_2 _2117_ (.Y(_1538_),
    .A(net712),
    .B(net694));
 sg13g2_nand2b_1 _2118_ (.Y(_1539_),
    .B(net737),
    .A_N(net736));
 sg13g2_nor4_2 _2119_ (.A(net723),
    .B(_1517_),
    .C(_1521_),
    .Y(_1540_),
    .D(_1539_));
 sg13g2_a21o_1 _2120_ (.A2(_1540_),
    .A1(net698),
    .B1(net712),
    .X(_1541_));
 sg13g2_nor2_1 _2121_ (.A(_1439_),
    .B(net727),
    .Y(_1542_));
 sg13g2_nand2b_1 _2122_ (.Y(_1543_),
    .B(net725),
    .A_N(net727));
 sg13g2_nor3_1 _2123_ (.A(_1500_),
    .B(_1528_),
    .C(_1543_),
    .Y(_1544_));
 sg13g2_nand2_1 _2124_ (.Y(_1545_),
    .A(net698),
    .B(_1542_));
 sg13g2_nor2_2 _2125_ (.A(_1509_),
    .B(_1543_),
    .Y(_1546_));
 sg13g2_nand2_1 _2126_ (.Y(_1547_),
    .A(net698),
    .B(_1546_));
 sg13g2_nand2b_1 _2127_ (.Y(_1548_),
    .B(_1547_),
    .A_N(_1541_));
 sg13g2_nor3_2 _2128_ (.A(net739),
    .B(_1436_),
    .C(_1521_),
    .Y(_1549_));
 sg13g2_nand3b_1 _2129_ (.B(net737),
    .C(_1520_),
    .Y(_1550_),
    .A_N(net739));
 sg13g2_nor2_2 _2130_ (.A(_1546_),
    .B(_1549_),
    .Y(_1551_));
 sg13g2_nand2b_1 _2131_ (.Y(_1552_),
    .B(_1550_),
    .A_N(_1546_));
 sg13g2_nor2_2 _2132_ (.A(_1509_),
    .B(_1521_),
    .Y(_1553_));
 sg13g2_nand2b_2 _2133_ (.Y(_1554_),
    .B(_1520_),
    .A_N(_1509_));
 sg13g2_nor4_2 _2134_ (.A(net735),
    .B(net723),
    .C(_1509_),
    .Y(_1555_),
    .D(_1521_));
 sg13g2_nor2b_2 _2135_ (.A(\sap_3_inst.controller.stage[3] ),
    .B_N(net717),
    .Y(_1556_));
 sg13g2_nand2b_2 _2136_ (.Y(_1557_),
    .B(net717),
    .A_N(\sap_3_inst.controller.stage[3] ));
 sg13g2_and2_1 _2137_ (.A(net711),
    .B(net710),
    .X(_1558_));
 sg13g2_nand2_2 _2138_ (.Y(_1559_),
    .A(net711),
    .B(net710));
 sg13g2_o21ai_1 _2139_ (.B1(_1555_),
    .Y(_1560_),
    .A1(net699),
    .A2(_1558_));
 sg13g2_and2_1 _2140_ (.A(net726),
    .B(net728),
    .X(_1561_));
 sg13g2_nand2_2 _2141_ (.Y(_1562_),
    .A(net726),
    .B(net728));
 sg13g2_and2_1 _2142_ (.A(net740),
    .B(net741),
    .X(_1563_));
 sg13g2_nand2_1 _2143_ (.Y(_1564_),
    .A(net740),
    .B(net741));
 sg13g2_nand2_2 _2144_ (.Y(_1565_),
    .A(net737),
    .B(_1563_));
 sg13g2_nor2_1 _2145_ (.A(_1521_),
    .B(net709),
    .Y(_1566_));
 sg13g2_nand3_1 _2146_ (.B(net726),
    .C(net728),
    .A(net738),
    .Y(_1567_));
 sg13g2_nor2_2 _2147_ (.A(_1509_),
    .B(_1562_),
    .Y(_1568_));
 sg13g2_nor4_2 _2148_ (.A(_1542_),
    .B(_1555_),
    .C(_1566_),
    .Y(_1569_),
    .D(_1568_));
 sg13g2_nand2_1 _2149_ (.Y(_1570_),
    .A(net699),
    .B(_1568_));
 sg13g2_nand2_1 _2150_ (.Y(_1571_),
    .A(_1560_),
    .B(_1570_));
 sg13g2_o21ai_1 _2151_ (.B1(_1551_),
    .Y(_1572_),
    .A1(_1569_),
    .A2(_1571_));
 sg13g2_nor2b_2 _2152_ (.A(net740),
    .B_N(net741),
    .Y(_1573_));
 sg13g2_nand2b_2 _2153_ (.Y(_1574_),
    .B(net741),
    .A_N(net740));
 sg13g2_nor4_2 _2154_ (.A(net735),
    .B(net737),
    .C(_1562_),
    .Y(_1575_),
    .D(_1574_));
 sg13g2_nand3_1 _2155_ (.B(_1561_),
    .C(_1573_),
    .A(_1522_),
    .Y(_1576_));
 sg13g2_and2_1 _2156_ (.A(_1533_),
    .B(_1556_),
    .X(_1577_));
 sg13g2_nand2_2 _2157_ (.Y(_1578_),
    .A(_1533_),
    .B(net710));
 sg13g2_a22oi_1 _2158_ (.Y(_1579_),
    .B1(_1533_),
    .B2(net710),
    .A2(_1527_),
    .A1(_1499_));
 sg13g2_nand2_1 _2159_ (.Y(_1580_),
    .A(net694),
    .B(_1578_));
 sg13g2_nor2_2 _2160_ (.A(_1536_),
    .B(_1557_),
    .Y(_1581_));
 sg13g2_nand2_2 _2161_ (.Y(_1582_),
    .A(_1535_),
    .B(net710));
 sg13g2_nor2_2 _2162_ (.A(_1567_),
    .B(_1574_),
    .Y(_1583_));
 sg13g2_nand2b_2 _2163_ (.Y(_1584_),
    .B(_1573_),
    .A_N(_1567_));
 sg13g2_nand2_1 _2164_ (.Y(_1585_),
    .A(_1581_),
    .B(_1583_));
 sg13g2_o21ai_1 _2165_ (.B1(_1585_),
    .Y(_1586_),
    .A1(_1576_),
    .A2(_1579_));
 sg13g2_nor3_2 _2166_ (.A(net738),
    .B(_1507_),
    .C(_1562_),
    .Y(_1587_));
 sg13g2_nand3_1 _2167_ (.B(_1506_),
    .C(_1561_),
    .A(_1436_),
    .Y(_1588_));
 sg13g2_nor4_2 _2168_ (.A(net735),
    .B(net737),
    .C(_1521_),
    .Y(_1589_),
    .D(_1574_));
 sg13g2_nand3_1 _2169_ (.B(_1522_),
    .C(_1573_),
    .A(_1520_),
    .Y(_1590_));
 sg13g2_and2_1 _2170_ (.A(_1522_),
    .B(_1563_),
    .X(_1591_));
 sg13g2_and4_1 _2171_ (.A(_1518_),
    .B(_1522_),
    .C(_1561_),
    .D(_1563_),
    .X(_1592_));
 sg13g2_nand4_1 _2172_ (.B(_1522_),
    .C(_1561_),
    .A(_1518_),
    .Y(_1593_),
    .D(_1563_));
 sg13g2_nand3_1 _2173_ (.B(_1590_),
    .C(_1593_),
    .A(_1588_),
    .Y(_1594_));
 sg13g2_nand3b_1 _2174_ (.B(net741),
    .C(net736),
    .Y(_1595_),
    .A_N(net739));
 sg13g2_nor4_2 _2175_ (.A(net738),
    .B(_1519_),
    .C(_1562_),
    .Y(_1596_),
    .D(_1595_));
 sg13g2_or4_1 _2176_ (.A(net737),
    .B(_1519_),
    .C(_1562_),
    .D(_1595_),
    .X(_1597_));
 sg13g2_nand2_1 _2177_ (.Y(_1598_),
    .A(_1516_),
    .B(_1561_));
 sg13g2_nor3_2 _2178_ (.A(net738),
    .B(_1517_),
    .C(_1562_),
    .Y(_1599_));
 sg13g2_inv_1 _2179_ (.Y(_1600_),
    .A(_1599_));
 sg13g2_or2_1 _2180_ (.X(_1601_),
    .B(_1599_),
    .A(_1596_));
 sg13g2_or2_1 _2181_ (.X(_1602_),
    .B(_1601_),
    .A(_1594_));
 sg13g2_nor3_1 _2182_ (.A(_1519_),
    .B(_1567_),
    .C(_1595_),
    .Y(_1603_));
 sg13g2_or3_1 _2183_ (.A(_1519_),
    .B(_1567_),
    .C(_1595_),
    .X(_1604_));
 sg13g2_nor2_2 _2184_ (.A(_1517_),
    .B(_1567_),
    .Y(_1605_));
 sg13g2_or2_1 _2185_ (.X(_1606_),
    .B(_1567_),
    .A(_1517_));
 sg13g2_nor2_2 _2186_ (.A(net707),
    .B(_1605_),
    .Y(_1607_));
 sg13g2_nand2_1 _2187_ (.Y(_1608_),
    .A(_1604_),
    .B(_1606_));
 sg13g2_nor2_2 _2188_ (.A(_1507_),
    .B(net722),
    .Y(_1609_));
 sg13g2_nand2_1 _2189_ (.Y(_1610_),
    .A(_1506_),
    .B(_1523_));
 sg13g2_nor2_1 _2190_ (.A(net722),
    .B(_1595_),
    .Y(_1611_));
 sg13g2_or2_1 _2191_ (.X(_1612_),
    .B(_1595_),
    .A(_1524_));
 sg13g2_nand4_1 _2192_ (.B(_1590_),
    .C(_1610_),
    .A(_1554_),
    .Y(_1613_),
    .D(_1612_));
 sg13g2_nor2b_2 _2193_ (.A(net731),
    .B_N(net729),
    .Y(_1614_));
 sg13g2_and2_1 _2194_ (.A(_1609_),
    .B(_1614_),
    .X(_1615_));
 sg13g2_nand3_1 _2195_ (.B(_1523_),
    .C(_1614_),
    .A(_1506_),
    .Y(_1616_));
 sg13g2_nor4_1 _2196_ (.A(_1594_),
    .B(_1601_),
    .C(_1608_),
    .D(_1613_),
    .Y(_1617_));
 sg13g2_nor2b_1 _2197_ (.A(_1586_),
    .B_N(net680),
    .Y(_1618_));
 sg13g2_nand2b_1 _2198_ (.Y(_1619_),
    .B(net680),
    .A_N(_1586_));
 sg13g2_nor2_2 _2199_ (.A(_1437_),
    .B(net730),
    .Y(_1620_));
 sg13g2_mux4_1 _2200_ (.S0(net732),
    .A0(\sap_3_inst.alu.flags[0] ),
    .A1(net720),
    .A2(\sap_3_inst.alu.flags[2] ),
    .A3(\sap_3_inst.alu.flags[3] ),
    .S1(net730),
    .X(_1621_));
 sg13g2_xnor2_1 _2201_ (.Y(_1622_),
    .A(net735),
    .B(_1621_));
 sg13g2_nand2_2 _2202_ (.Y(_1623_),
    .A(net700),
    .B(_1622_));
 sg13g2_nor2b_1 _2203_ (.A(net717),
    .B_N(net716),
    .Y(_1624_));
 sg13g2_nand2b_1 _2204_ (.Y(_1625_),
    .B(net716),
    .A_N(net717));
 sg13g2_and2_1 _2205_ (.A(net711),
    .B(net704),
    .X(_1626_));
 sg13g2_nand2_2 _2206_ (.Y(_1627_),
    .A(net711),
    .B(net704));
 sg13g2_nor2_1 _2207_ (.A(_1577_),
    .B(_1626_),
    .Y(_1628_));
 sg13g2_a21oi_1 _2208_ (.A1(_1623_),
    .A2(_1628_),
    .Y(_1629_),
    .B1(_1600_));
 sg13g2_a21oi_1 _2209_ (.A1(_1579_),
    .A2(_1627_),
    .Y(_1630_),
    .B1(_1597_));
 sg13g2_nor3_1 _2210_ (.A(net680),
    .B(_1629_),
    .C(_1630_),
    .Y(_1631_));
 sg13g2_or3_1 _2211_ (.A(net680),
    .B(_1629_),
    .C(_1630_),
    .X(_1632_));
 sg13g2_and2_1 _2212_ (.A(net717),
    .B(net716),
    .X(_1633_));
 sg13g2_nand2_1 _2213_ (.Y(_1634_),
    .A(net717),
    .B(net716));
 sg13g2_and3_2 _2214_ (.X(_1635_),
    .A(\sap_3_inst.controller.stage[2] ),
    .B(net719),
    .C(net718));
 sg13g2_nand2_2 _2215_ (.Y(_1636_),
    .A(net716),
    .B(_1635_));
 sg13g2_inv_2 _2216_ (.Y(_1637_),
    .A(_1636_));
 sg13g2_and2_1 _2217_ (.A(net718),
    .B(net705),
    .X(_1638_));
 sg13g2_and2_1 _2218_ (.A(_1533_),
    .B(net705),
    .X(_1639_));
 sg13g2_nand2_1 _2219_ (.Y(_1640_),
    .A(_1533_),
    .B(net705));
 sg13g2_and2_1 _2220_ (.A(net711),
    .B(_1633_),
    .X(_1641_));
 sg13g2_a22oi_1 _2221_ (.Y(_1642_),
    .B1(_1633_),
    .B2(net711),
    .A2(net704),
    .A1(_1533_));
 sg13g2_nand2_1 _2222_ (.Y(_1643_),
    .A(_1578_),
    .B(_1642_));
 sg13g2_nand4_1 _2223_ (.B(_1623_),
    .C(_1636_),
    .A(_1578_),
    .Y(_1644_),
    .D(_1642_));
 sg13g2_nand2_1 _2224_ (.Y(_1645_),
    .A(_1605_),
    .B(_1644_));
 sg13g2_and2_1 _2225_ (.A(net714),
    .B(net704),
    .X(_1646_));
 sg13g2_nand2_2 _2226_ (.Y(_1647_),
    .A(net714),
    .B(net705));
 sg13g2_nand2_1 _2227_ (.Y(_1648_),
    .A(_1578_),
    .B(_1647_));
 sg13g2_nand2b_1 _2228_ (.Y(_1649_),
    .B(_1623_),
    .A_N(_1648_));
 sg13g2_nand2_1 _2229_ (.Y(_1650_),
    .A(_1587_),
    .B(_1649_));
 sg13g2_a22oi_1 _2230_ (.Y(_1651_),
    .B1(_1633_),
    .B2(net714),
    .A2(net704),
    .A1(net711));
 sg13g2_nand2_1 _2231_ (.Y(_1652_),
    .A(_1579_),
    .B(_1651_));
 sg13g2_a22oi_1 _2232_ (.Y(_1653_),
    .B1(_1652_),
    .B2(_1615_),
    .A2(_1643_),
    .A1(net707));
 sg13g2_a22oi_1 _2233_ (.Y(_1654_),
    .B1(_1647_),
    .B2(_1579_),
    .A2(_1593_),
    .A1(_1590_));
 sg13g2_nor3_2 _2234_ (.A(net729),
    .B(_1507_),
    .C(net722),
    .Y(_1655_));
 sg13g2_nor3_1 _2235_ (.A(net722),
    .B(_1528_),
    .C(_1595_),
    .Y(_1656_));
 sg13g2_nor4_1 _2236_ (.A(net722),
    .B(_1528_),
    .C(_1595_),
    .D(_1625_),
    .Y(_1657_));
 sg13g2_nand2_2 _2237_ (.Y(_1658_),
    .A(_1527_),
    .B(net705));
 sg13g2_or2_1 _2238_ (.X(_1659_),
    .B(_1658_),
    .A(_1612_));
 sg13g2_a21o_1 _2239_ (.A2(_1655_),
    .A1(net687),
    .B1(_1657_),
    .X(_1660_));
 sg13g2_nor3_1 _2240_ (.A(net723),
    .B(_1507_),
    .C(net722),
    .Y(_1661_));
 sg13g2_nand3_1 _2241_ (.B(_1506_),
    .C(_1523_),
    .A(_1504_),
    .Y(_1662_));
 sg13g2_a21oi_1 _2242_ (.A1(_1579_),
    .A2(_1627_),
    .Y(_1663_),
    .B1(_1662_));
 sg13g2_nor2_1 _2243_ (.A(net694),
    .B(_1554_),
    .Y(_1664_));
 sg13g2_nand2_1 _2244_ (.Y(_1665_),
    .A(net696),
    .B(_1553_));
 sg13g2_a22oi_1 _2245_ (.Y(_1666_),
    .B1(_1665_),
    .B2(_1604_),
    .A2(_1636_),
    .A1(net694));
 sg13g2_nor4_1 _2246_ (.A(_1654_),
    .B(_1660_),
    .C(_1663_),
    .D(_1666_),
    .Y(_1667_));
 sg13g2_nand4_1 _2247_ (.B(_1650_),
    .C(_1653_),
    .A(_1645_),
    .Y(_1668_),
    .D(_1667_));
 sg13g2_o21ai_1 _2248_ (.B1(_1619_),
    .Y(_1669_),
    .A1(_1632_),
    .A2(_1668_));
 sg13g2_a21oi_1 _2249_ (.A1(_1569_),
    .A2(_1669_),
    .Y(_1670_),
    .B1(_1572_));
 sg13g2_o21ai_1 _2250_ (.B1(_1538_),
    .Y(_1671_),
    .A1(_1548_),
    .A2(_1670_));
 sg13g2_nand2_1 _2251_ (.Y(_1672_),
    .A(net703),
    .B(_1671_));
 sg13g2_a22oi_1 _2252_ (.Y(_1673_),
    .B1(_1537_),
    .B2(_1672_),
    .A2(net715),
    .A1(_1499_));
 sg13g2_and2_1 _2253_ (.A(net715),
    .B(_1556_),
    .X(_1674_));
 sg13g2_nand2_2 _2254_ (.Y(_1675_),
    .A(net715),
    .B(net710));
 sg13g2_a21oi_1 _2255_ (.A1(net709),
    .A2(net685),
    .Y(_1676_),
    .B1(_1538_));
 sg13g2_o21ai_1 _2256_ (.B1(_1604_),
    .Y(_1677_),
    .A1(_1438_),
    .A2(_1610_));
 sg13g2_nand2_1 _2257_ (.Y(_1678_),
    .A(_1593_),
    .B(_1597_));
 sg13g2_nor4_1 _2258_ (.A(net707),
    .B(_1609_),
    .C(net706),
    .D(_1678_),
    .Y(_1679_));
 sg13g2_o21ai_1 _2259_ (.B1(_1589_),
    .Y(_1680_),
    .A1(_1580_),
    .A2(_1646_));
 sg13g2_o21ai_1 _2260_ (.B1(_1648_),
    .Y(_1681_),
    .A1(_1592_),
    .A2(_1679_));
 sg13g2_o21ai_1 _2261_ (.B1(net684),
    .Y(_1682_),
    .A1(net706),
    .A2(_1655_));
 sg13g2_o21ai_1 _2262_ (.B1(_1682_),
    .Y(_1683_),
    .A1(_1578_),
    .A2(_1616_));
 sg13g2_or2_1 _2263_ (.X(_1684_),
    .B(_1630_),
    .A(net700));
 sg13g2_or2_1 _2264_ (.X(_1685_),
    .B(_1651_),
    .A(_1616_));
 sg13g2_or3_1 _2265_ (.A(net733),
    .B(_1616_),
    .C(_1642_),
    .X(_1686_));
 sg13g2_nor2_1 _2266_ (.A(net714),
    .B(_1634_),
    .Y(_1687_));
 sg13g2_or2_1 _2267_ (.X(_1688_),
    .B(_1638_),
    .A(_1577_));
 sg13g2_o21ai_1 _2268_ (.B1(net707),
    .Y(_1689_),
    .A1(_1687_),
    .A2(_1688_));
 sg13g2_nor2_2 _2269_ (.A(_1528_),
    .B(_1557_),
    .Y(_1690_));
 sg13g2_nor2_1 _2270_ (.A(_1536_),
    .B(_1625_),
    .Y(_1691_));
 sg13g2_or2_1 _2271_ (.X(_1692_),
    .B(_1691_),
    .A(_1690_));
 sg13g2_a22oi_1 _2272_ (.Y(_1693_),
    .B1(_1692_),
    .B2(net706),
    .A2(_1655_),
    .A1(net687));
 sg13g2_nand4_1 _2273_ (.B(_1686_),
    .C(_1689_),
    .A(_1685_),
    .Y(_1694_),
    .D(_1693_));
 sg13g2_nor4_1 _2274_ (.A(_1663_),
    .B(_1683_),
    .C(_1684_),
    .D(_1694_),
    .Y(_1695_));
 sg13g2_a22oi_1 _2275_ (.Y(_1696_),
    .B1(_1681_),
    .B2(_1695_),
    .A2(_1680_),
    .A1(_1679_));
 sg13g2_inv_1 _2276_ (.Y(_1697_),
    .A(_1696_));
 sg13g2_a21oi_2 _2277_ (.B1(_1584_),
    .Y(_1698_),
    .A2(_1647_),
    .A1(_1559_));
 sg13g2_nand2_2 _2278_ (.Y(_1699_),
    .A(_1555_),
    .B(_1577_));
 sg13g2_inv_1 _2279_ (.Y(_1700_),
    .A(_1699_));
 sg13g2_and2_1 _2280_ (.A(_1544_),
    .B(net709),
    .X(_1701_));
 sg13g2_nor4_1 _2281_ (.A(net689),
    .B(_1664_),
    .C(_1700_),
    .D(_1701_),
    .Y(_1702_));
 sg13g2_a22oi_1 _2282_ (.Y(_1703_),
    .B1(net704),
    .B2(net714),
    .A2(net710),
    .A1(net711));
 sg13g2_nand2_1 _2283_ (.Y(_1704_),
    .A(_1559_),
    .B(_1647_));
 sg13g2_nor3_1 _2284_ (.A(_1584_),
    .B(net708),
    .C(_1703_),
    .Y(_1705_));
 sg13g2_a221oi_1 _2285_ (.B2(net724),
    .C1(_1571_),
    .B1(_1705_),
    .A1(_1586_),
    .Y(_1706_),
    .A2(_1604_));
 sg13g2_or3_1 _2286_ (.A(net696),
    .B(_1687_),
    .C(_1688_),
    .X(_1707_));
 sg13g2_nor2_1 _2287_ (.A(net695),
    .B(_1622_),
    .Y(_1708_));
 sg13g2_nor2_1 _2288_ (.A(_1606_),
    .B(_1708_),
    .Y(_1709_));
 sg13g2_a21oi_1 _2289_ (.A1(_1707_),
    .A2(_1709_),
    .Y(_1710_),
    .B1(_1629_));
 sg13g2_and4_1 _2290_ (.A(_1650_),
    .B(_1702_),
    .C(_1706_),
    .D(_1710_),
    .X(_1711_));
 sg13g2_nor2_1 _2291_ (.A(net722),
    .B(_1564_),
    .Y(_1712_));
 sg13g2_o21ai_1 _2292_ (.B1(_1511_),
    .Y(_1713_),
    .A1(net722),
    .A2(_1564_));
 sg13g2_nor2_1 _2293_ (.A(_1540_),
    .B(_1713_),
    .Y(_1714_));
 sg13g2_or2_1 _2294_ (.X(_1715_),
    .B(_1713_),
    .A(_1540_));
 sg13g2_nand2_2 _2295_ (.Y(_1716_),
    .A(net734),
    .B(_1504_));
 sg13g2_and2_1 _2296_ (.A(net698),
    .B(_1716_),
    .X(_1717_));
 sg13g2_nor2_1 _2297_ (.A(_1551_),
    .B(_1717_),
    .Y(_1718_));
 sg13g2_a221oi_1 _2298_ (.B2(_1547_),
    .C1(_1715_),
    .B1(_1718_),
    .A1(_1697_),
    .Y(_1719_),
    .A2(_1711_));
 sg13g2_and3_1 _2299_ (.X(_1720_),
    .A(_1510_),
    .B(net698),
    .C(net709));
 sg13g2_nor3_1 _2300_ (.A(_1541_),
    .B(_1719_),
    .C(_1720_),
    .Y(_1721_));
 sg13g2_o21ai_1 _2301_ (.B1(net703),
    .Y(_1722_),
    .A1(_1676_),
    .A2(_1721_));
 sg13g2_and3_2 _2302_ (.X(_1723_),
    .A(_1537_),
    .B(net567),
    .C(_1722_));
 sg13g2_nand2_1 _2303_ (.Y(_1724_),
    .A(_1620_),
    .B(_1698_));
 sg13g2_nor2_1 _2304_ (.A(_1627_),
    .B(_1662_),
    .Y(_1725_));
 sg13g2_a221oi_1 _2305_ (.B2(_1594_),
    .C1(_1725_),
    .B1(_1646_),
    .A1(_1608_),
    .Y(_1726_),
    .A2(_1637_));
 sg13g2_o21ai_1 _2306_ (.B1(net714),
    .Y(_1727_),
    .A1(net710),
    .A2(net705));
 sg13g2_nor2_1 _2307_ (.A(_1612_),
    .B(_1727_),
    .Y(_1728_));
 sg13g2_nand2b_1 _2308_ (.Y(_1729_),
    .B(net706),
    .A_N(_1727_));
 sg13g2_o21ai_1 _2309_ (.B1(_1655_),
    .Y(_1730_),
    .A1(net697),
    .A2(net684));
 sg13g2_a21o_1 _2310_ (.A2(_1730_),
    .A1(_1729_),
    .B1(_1437_),
    .X(_1731_));
 sg13g2_a21oi_1 _2311_ (.A1(_1604_),
    .A2(_1606_),
    .Y(_1732_),
    .B1(_1642_));
 sg13g2_nor2_1 _2312_ (.A(_1660_),
    .B(_1732_),
    .Y(_1733_));
 sg13g2_and4_1 _2313_ (.A(_1685_),
    .B(_1726_),
    .C(_1731_),
    .D(_1733_),
    .X(_1734_));
 sg13g2_a22oi_1 _2314_ (.Y(_1735_),
    .B1(_1734_),
    .B2(_1631_),
    .A2(_1724_),
    .A1(_1618_));
 sg13g2_nand3_1 _2315_ (.B(net689),
    .C(_1717_),
    .A(net732),
    .Y(_1736_));
 sg13g2_nand2_1 _2316_ (.Y(_1737_),
    .A(net739),
    .B(_1701_));
 sg13g2_nand3_1 _2317_ (.B(_1736_),
    .C(_1737_),
    .A(_1699_),
    .Y(_1738_));
 sg13g2_o21ai_1 _2318_ (.B1(net683),
    .Y(_1739_),
    .A1(_1509_),
    .A2(_1545_));
 sg13g2_inv_1 _2319_ (.Y(_1740_),
    .A(_1739_));
 sg13g2_o21ai_1 _2320_ (.B1(_1740_),
    .Y(_1741_),
    .A1(_1735_),
    .A2(_1738_));
 sg13g2_a21oi_1 _2321_ (.A1(net739),
    .A2(_1720_),
    .Y(_1742_),
    .B1(net712));
 sg13g2_nand3_1 _2322_ (.B(net709),
    .C(net684),
    .A(net740),
    .Y(_1743_));
 sg13g2_nor2_1 _2323_ (.A(\sap_3_inst.controller.stage[2] ),
    .B(_1527_),
    .Y(_1744_));
 sg13g2_o21ai_1 _2324_ (.B1(net702),
    .Y(_1745_),
    .A1(_1500_),
    .A2(_1527_));
 sg13g2_a221oi_1 _2325_ (.B2(net712),
    .C1(_1745_),
    .B1(_1743_),
    .A1(_1741_),
    .Y(_1746_),
    .A2(_1742_));
 sg13g2_nand3_1 _2326_ (.B(net709),
    .C(net684),
    .A(net741),
    .Y(_1747_));
 sg13g2_and2_1 _2327_ (.A(_1514_),
    .B(_1747_),
    .X(_1748_));
 sg13g2_nor2b_1 _2328_ (.A(_1616_),
    .B_N(_1641_),
    .Y(_1749_));
 sg13g2_nand2_1 _2329_ (.Y(_1750_),
    .A(_1615_),
    .B(_1641_));
 sg13g2_nor2_1 _2330_ (.A(net733),
    .B(_1750_),
    .Y(_1751_));
 sg13g2_nand4_1 _2331_ (.B(net724),
    .C(net698),
    .A(net735),
    .Y(_1752_),
    .D(_1549_));
 sg13g2_nor2_1 _2332_ (.A(_1607_),
    .B(_1658_),
    .Y(_1753_));
 sg13g2_nand2_1 _2333_ (.Y(_1754_),
    .A(_1511_),
    .B(_1569_));
 sg13g2_nand4_1 _2334_ (.B(net699),
    .C(_1565_),
    .A(net742),
    .Y(_1755_),
    .D(_1754_));
 sg13g2_nand4_1 _2335_ (.B(_1583_),
    .C(net681),
    .A(net723),
    .Y(_1756_),
    .D(_1646_));
 sg13g2_nand2_1 _2336_ (.Y(_1757_),
    .A(net696),
    .B(net706));
 sg13g2_nand2_1 _2337_ (.Y(_1758_),
    .A(_1682_),
    .B(_1757_));
 sg13g2_nor3_1 _2338_ (.A(_1751_),
    .B(net679),
    .C(_1758_),
    .Y(_1759_));
 sg13g2_and4_1 _2339_ (.A(_1752_),
    .B(_1755_),
    .C(_1756_),
    .D(_1759_),
    .X(_1760_));
 sg13g2_a21oi_2 _2340_ (.B1(_1748_),
    .Y(_1761_),
    .A2(_1760_),
    .A1(_1515_));
 sg13g2_a21o_2 _2341_ (.A2(_1760_),
    .A1(_1515_),
    .B1(_1748_),
    .X(_1762_));
 sg13g2_a22oi_1 _2342_ (.Y(_1763_),
    .B1(_1623_),
    .B2(_1578_),
    .A2(_1598_),
    .A1(_1588_));
 sg13g2_nand3_1 _2343_ (.B(_1593_),
    .C(_1597_),
    .A(_1590_),
    .Y(_1764_));
 sg13g2_o21ai_1 _2344_ (.B1(_1580_),
    .Y(_1765_),
    .A1(_1677_),
    .A2(_1764_));
 sg13g2_nor3_1 _2345_ (.A(net723),
    .B(_1612_),
    .C(_1727_),
    .Y(_1766_));
 sg13g2_nand2_1 _2346_ (.Y(_1767_),
    .A(_1533_),
    .B(_1633_));
 sg13g2_a22oi_1 _2347_ (.Y(_1768_),
    .B1(_1658_),
    .B2(_1767_),
    .A2(_1606_),
    .A1(_1604_));
 sg13g2_nor4_1 _2348_ (.A(_1664_),
    .B(_1732_),
    .C(_1766_),
    .D(_1768_),
    .Y(_1769_));
 sg13g2_nand3b_1 _2349_ (.B(_1765_),
    .C(_1769_),
    .Y(_1770_),
    .A_N(net681));
 sg13g2_o21ai_1 _2350_ (.B1(_1619_),
    .Y(_1771_),
    .A1(_1763_),
    .A2(_1770_));
 sg13g2_nand3_1 _2351_ (.B(_1570_),
    .C(_1771_),
    .A(_1503_),
    .Y(_1772_));
 sg13g2_inv_1 _2352_ (.Y(_1773_),
    .A(_1772_));
 sg13g2_nor2_2 _2353_ (.A(_1436_),
    .B(_1563_),
    .Y(_1774_));
 sg13g2_a21o_1 _2354_ (.A2(_1774_),
    .A1(net697),
    .B1(net682),
    .X(_1775_));
 sg13g2_o21ai_1 _2355_ (.B1(_1614_),
    .Y(_1776_),
    .A1(_1698_),
    .A2(_1728_));
 sg13g2_a22oi_1 _2356_ (.Y(_1777_),
    .B1(_1774_),
    .B2(_1544_),
    .A2(_1655_),
    .A1(net687));
 sg13g2_a22oi_1 _2357_ (.Y(_1778_),
    .B1(_1634_),
    .B2(_1656_),
    .A2(net688),
    .A1(_1555_));
 sg13g2_and4_1 _2358_ (.A(_1685_),
    .B(_1686_),
    .C(_1777_),
    .D(_1778_),
    .X(_1779_));
 sg13g2_o21ai_1 _2359_ (.B1(_1626_),
    .Y(_1780_),
    .A1(_1596_),
    .A2(_1599_));
 sg13g2_and2_1 _2360_ (.A(net734),
    .B(net731),
    .X(_1781_));
 sg13g2_nor2_1 _2361_ (.A(_1438_),
    .B(_1781_),
    .Y(_1782_));
 sg13g2_nor4_1 _2362_ (.A(_1438_),
    .B(_1500_),
    .C(_1528_),
    .D(_1781_),
    .Y(_1783_));
 sg13g2_o21ai_1 _2363_ (.B1(_1783_),
    .Y(_1784_),
    .A1(_1546_),
    .A2(_1549_));
 sg13g2_and4_1 _2364_ (.A(_1699_),
    .B(net682),
    .C(_1780_),
    .D(_1784_),
    .X(_1785_));
 sg13g2_nor2_1 _2365_ (.A(_1554_),
    .B(_1559_),
    .Y(_1786_));
 sg13g2_nand4_1 _2366_ (.B(_1776_),
    .C(_1779_),
    .A(_1726_),
    .Y(_1787_),
    .D(_1785_));
 sg13g2_a21oi_1 _2367_ (.A1(_1775_),
    .A2(_1787_),
    .Y(_1788_),
    .B1(net712));
 sg13g2_a21oi_1 _2368_ (.A1(net684),
    .A2(_1774_),
    .Y(_1789_),
    .B1(_1538_));
 sg13g2_nor4_2 _2369_ (.A(_1502_),
    .B(_1526_),
    .C(_1788_),
    .Y(_1790_),
    .D(_1789_));
 sg13g2_inv_1 _2370_ (.Y(_1791_),
    .A(_1790_));
 sg13g2_nor2_1 _2371_ (.A(_1772_),
    .B(_1790_),
    .Y(_1792_));
 sg13g2_or2_1 _2372_ (.X(_1793_),
    .B(_1790_),
    .A(_1772_));
 sg13g2_nor3_2 _2373_ (.A(_1746_),
    .B(_1761_),
    .C(_1793_),
    .Y(_1794_));
 sg13g2_and3_2 _2374_ (.X(_1795_),
    .A(_1746_),
    .B(_1762_),
    .C(_1792_));
 sg13g2_nor3_2 _2375_ (.A(net662),
    .B(_1761_),
    .C(_1791_),
    .Y(_1796_));
 sg13g2_and3_2 _2376_ (.X(_1797_),
    .A(net662),
    .B(_1762_),
    .C(_1772_));
 sg13g2_nor3_2 _2377_ (.A(net662),
    .B(_1762_),
    .C(_1793_),
    .Y(_1798_));
 sg13g2_and3_2 _2378_ (.X(_1799_),
    .A(net662),
    .B(_1762_),
    .C(_1790_));
 sg13g2_and3_2 _2379_ (.X(_1800_),
    .A(net662),
    .B(_1761_),
    .C(_1792_));
 sg13g2_nor3_2 _2380_ (.A(net662),
    .B(_1762_),
    .C(_1791_),
    .Y(_1801_));
 sg13g2_and3_2 _2381_ (.X(_1802_),
    .A(net662),
    .B(_1761_),
    .C(_1772_));
 sg13g2_nor3_2 _2382_ (.A(net662),
    .B(_1761_),
    .C(_1773_),
    .Y(_1803_));
 sg13g2_a221oi_1 _2383_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .C1(net638),
    .B1(net623),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .Y(_1804_),
    .A2(net625));
 sg13g2_a22oi_1 _2384_ (.Y(_1805_),
    .B1(net627),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .A2(net635),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ));
 sg13g2_a22oi_1 _2385_ (.Y(_1806_),
    .B1(net619),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .A2(net633),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ));
 sg13g2_a22oi_1 _2386_ (.Y(_1807_),
    .B1(net629),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .A2(net677),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ));
 sg13g2_nand3_1 _2387_ (.B(_1806_),
    .C(_1807_),
    .A(_1805_),
    .Y(_1808_));
 sg13g2_a221oi_1 _2388_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .C1(_1808_),
    .B1(net621),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ),
    .Y(_1809_),
    .A2(net631));
 sg13g2_a22oi_1 _2389_ (.Y(_1810_),
    .B1(_1804_),
    .B2(_1809_),
    .A2(net638),
    .A1(_1490_));
 sg13g2_and2_1 _2390_ (.A(_1723_),
    .B(_1810_),
    .X(_1811_));
 sg13g2_nand2_1 _2391_ (.Y(_1812_),
    .A(net712),
    .B(net685));
 sg13g2_nor2_1 _2392_ (.A(net709),
    .B(_1812_),
    .Y(_1813_));
 sg13g2_nor2_2 _2393_ (.A(_1550_),
    .B(_1559_),
    .Y(_1814_));
 sg13g2_a22oi_1 _2394_ (.Y(_1815_),
    .B1(_1690_),
    .B2(_1655_),
    .A2(_1661_),
    .A1(_1639_));
 sg13g2_nor2_1 _2395_ (.A(net736),
    .B(_1815_),
    .Y(_1816_));
 sg13g2_nor3_1 _2396_ (.A(net724),
    .B(_1559_),
    .C(_1584_),
    .Y(_1817_));
 sg13g2_a21oi_1 _2397_ (.A1(_1578_),
    .A2(_1640_),
    .Y(_1818_),
    .B1(_1612_));
 sg13g2_or4_1 _2398_ (.A(net689),
    .B(_1816_),
    .C(_1817_),
    .D(_1818_),
    .X(_1819_));
 sg13g2_o21ai_1 _2399_ (.B1(_1819_),
    .Y(_1820_),
    .A1(_1551_),
    .A2(_1814_));
 sg13g2_nor2_1 _2400_ (.A(net695),
    .B(_1565_),
    .Y(_1821_));
 sg13g2_nand2_1 _2401_ (.Y(_1822_),
    .A(_1540_),
    .B(_1577_));
 sg13g2_nand2_1 _2402_ (.Y(_1823_),
    .A(_1715_),
    .B(_1822_));
 sg13g2_a21oi_1 _2403_ (.A1(_1510_),
    .A2(_1821_),
    .Y(_1824_),
    .B1(_1823_));
 sg13g2_a21oi_1 _2404_ (.A1(net683),
    .A2(_1820_),
    .Y(_1825_),
    .B1(_1824_));
 sg13g2_a21oi_1 _2405_ (.A1(_1515_),
    .A2(_1825_),
    .Y(_1826_),
    .B1(_1813_));
 sg13g2_inv_4 _2406_ (.A(_1826_),
    .Y(_1827_));
 sg13g2_nor3_2 _2407_ (.A(net723),
    .B(_1584_),
    .C(_1647_),
    .Y(_1828_));
 sg13g2_a22oi_1 _2408_ (.Y(_1829_),
    .B1(_1828_),
    .B2(\sap_3_inst.alu.flags[7] ),
    .A2(_1827_),
    .A1(net743));
 sg13g2_a21oi_1 _2409_ (.A1(net713),
    .A2(_1675_),
    .Y(_1830_),
    .B1(_1526_));
 sg13g2_a21o_1 _2410_ (.A2(_1675_),
    .A1(net713),
    .B1(_1526_),
    .X(_1831_));
 sg13g2_nand3_1 _2411_ (.B(_1639_),
    .C(_1661_),
    .A(net733),
    .Y(_1832_));
 sg13g2_nand2_1 _2412_ (.Y(_1833_),
    .A(net686),
    .B(_1832_));
 sg13g2_nand2b_1 _2413_ (.Y(_1834_),
    .B(net734),
    .A_N(_1642_));
 sg13g2_a21oi_1 _2414_ (.A1(_1582_),
    .A2(_1834_),
    .Y(_1835_),
    .B1(_1616_));
 sg13g2_a21o_1 _2415_ (.A2(net685),
    .A1(_1568_),
    .B1(net689),
    .X(_1836_));
 sg13g2_and3_1 _2416_ (.X(_1837_),
    .A(net736),
    .B(_1655_),
    .C(_1690_));
 sg13g2_nor2_1 _2417_ (.A(_1576_),
    .B(net686),
    .Y(_1838_));
 sg13g2_nor2_1 _2418_ (.A(_1554_),
    .B(_1675_),
    .Y(_1839_));
 sg13g2_nand3b_1 _2419_ (.B(_1607_),
    .C(_1662_),
    .Y(_1840_),
    .A_N(_1838_));
 sg13g2_o21ai_1 _2420_ (.B1(_1833_),
    .Y(_1841_),
    .A1(_1602_),
    .A2(_1840_));
 sg13g2_nor4_1 _2421_ (.A(_1835_),
    .B(_1836_),
    .C(_1837_),
    .D(_1839_),
    .Y(_1842_));
 sg13g2_nand2_1 _2422_ (.Y(_1843_),
    .A(net689),
    .B(_1743_));
 sg13g2_a221oi_1 _2423_ (.B2(_1842_),
    .C1(_1715_),
    .B1(_1841_),
    .A1(net689),
    .Y(_1844_),
    .A2(_1743_));
 sg13g2_and2_1 _2424_ (.A(_1540_),
    .B(net685),
    .X(_1845_));
 sg13g2_nor3_1 _2425_ (.A(_1512_),
    .B(_1844_),
    .C(_1845_),
    .Y(_1846_));
 sg13g2_o21ai_1 _2426_ (.B1(net693),
    .Y(_1847_),
    .A1(_1831_),
    .A2(_1846_));
 sg13g2_nand2_1 _2427_ (.Y(_1848_),
    .A(net8),
    .B(_1847_));
 sg13g2_nand2_1 _2428_ (.Y(_1849_),
    .A(_1829_),
    .B(_1848_));
 sg13g2_a22oi_1 _2429_ (.Y(_1850_),
    .B1(net619),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ),
    .A2(net631),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ));
 sg13g2_a22oi_1 _2430_ (.Y(_1851_),
    .B1(net625),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .A2(net627),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ));
 sg13g2_a221oi_1 _2431_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .C1(net621),
    .B1(net635),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .Y(_1852_),
    .A2(net638));
 sg13g2_a22oi_1 _2432_ (.Y(_1853_),
    .B1(net633),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .A2(net677),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ));
 sg13g2_nand3_1 _2433_ (.B(_1852_),
    .C(_1853_),
    .A(_1850_),
    .Y(_1854_));
 sg13g2_a221oi_1 _2434_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .C1(_1854_),
    .B1(net623),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .Y(_1855_),
    .A2(net629));
 sg13g2_a21oi_1 _2435_ (.A1(_1851_),
    .A2(_1855_),
    .Y(_1856_),
    .B1(net565));
 sg13g2_or3_1 _2436_ (.A(_1811_),
    .B(_1849_),
    .C(_1856_),
    .X(net542));
 sg13g2_nor3_2 _2437_ (.A(net724),
    .B(_1576_),
    .C(_1675_),
    .Y(_1857_));
 sg13g2_inv_2 _2438_ (.Y(_1858_),
    .A(net675));
 sg13g2_mux2_1 _2439_ (.A0(\sap_3_inst.alu.flags[7] ),
    .A1(net542),
    .S(net675),
    .X(_0033_));
 sg13g2_a22oi_1 _2440_ (.Y(_1859_),
    .B1(net620),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .A2(net634),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ));
 sg13g2_a22oi_1 _2441_ (.Y(_1860_),
    .B1(_1801_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .A2(_1797_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ));
 sg13g2_and2_1 _2442_ (.A(_1859_),
    .B(_1860_),
    .X(_1861_));
 sg13g2_a221oi_1 _2443_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .C1(net639),
    .B1(net636),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ),
    .Y(_1862_),
    .A2(net677));
 sg13g2_a22oi_1 _2444_ (.Y(_1863_),
    .B1(net625),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .A2(net629),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ));
 sg13g2_a22oi_1 _2445_ (.Y(_1864_),
    .B1(net621),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .A2(net627),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ));
 sg13g2_and3_1 _2446_ (.X(_1865_),
    .A(_1862_),
    .B(_1863_),
    .C(_1864_));
 sg13g2_a22oi_1 _2447_ (.Y(_1866_),
    .B1(_1861_),
    .B2(_1865_),
    .A2(net639),
    .A1(_1479_));
 sg13g2_and2_1 _2448_ (.A(\sap_3_inst.alu.flags[6] ),
    .B(_1828_),
    .X(_1867_));
 sg13g2_a221oi_1 _2449_ (.B2(net7),
    .C1(_1867_),
    .B1(_1847_),
    .A1(net745),
    .Y(_1868_),
    .A2(_1827_));
 sg13g2_a22oi_1 _2450_ (.Y(_1869_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .A2(_1796_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ));
 sg13g2_a22oi_1 _2451_ (.Y(_1870_),
    .B1(net623),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .A2(_1795_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ));
 sg13g2_nand2_1 _2452_ (.Y(_1871_),
    .A(_1869_),
    .B(_1870_));
 sg13g2_a221oi_1 _2453_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .C1(net621),
    .B1(net627),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ),
    .Y(_1872_),
    .A2(net677));
 sg13g2_a22oi_1 _2454_ (.Y(_1873_),
    .B1(_1803_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ),
    .A2(net639),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ));
 sg13g2_a22oi_1 _2455_ (.Y(_1874_),
    .B1(net626),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .A2(net630),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ));
 sg13g2_nand3_1 _2456_ (.B(_1873_),
    .C(_1874_),
    .A(_1872_),
    .Y(_1875_));
 sg13g2_nor2_1 _2457_ (.A(_1871_),
    .B(_1875_),
    .Y(_1876_));
 sg13g2_o21ai_1 _2458_ (.B1(_1868_),
    .Y(_1877_),
    .A1(net565),
    .A2(_1876_));
 sg13g2_a21oi_2 _2459_ (.B1(_1877_),
    .Y(_1878_),
    .A2(_1866_),
    .A1(_1723_));
 sg13g2_inv_2 _2460_ (.Y(net23),
    .A(net547));
 sg13g2_nor2_1 _2461_ (.A(\sap_3_inst.alu.flags[6] ),
    .B(net675),
    .Y(_1879_));
 sg13g2_a21oi_1 _2462_ (.A1(net675),
    .A2(_1878_),
    .Y(_0032_),
    .B1(_1879_));
 sg13g2_and2_1 _2463_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .B(net629),
    .X(_1880_));
 sg13g2_a221oi_1 _2464_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .C1(_1880_),
    .B1(net625),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .Y(_1881_),
    .A2(net627));
 sg13g2_a21oi_1 _2465_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .A2(net635),
    .Y(_1882_),
    .B1(net638));
 sg13g2_a22oi_1 _2466_ (.Y(_1883_),
    .B1(net621),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .A2(net633),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ));
 sg13g2_a22oi_1 _2467_ (.Y(_1884_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .A2(net677),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ));
 sg13g2_nand3_1 _2468_ (.B(_1883_),
    .C(_1884_),
    .A(_1882_),
    .Y(_1885_));
 sg13g2_a221oi_1 _2469_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .C1(_1885_),
    .B1(net619),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .Y(_1886_),
    .A2(net623));
 sg13g2_a22oi_1 _2470_ (.Y(_1887_),
    .B1(_1881_),
    .B2(_1886_),
    .A2(net639),
    .A1(_1475_));
 sg13g2_a22oi_1 _2471_ (.Y(_1888_),
    .B1(_1828_),
    .B2(\sap_3_inst.alu.flags[5] ),
    .A2(_1827_),
    .A1(net747));
 sg13g2_nand2_1 _2472_ (.Y(_1889_),
    .A(net6),
    .B(_1847_));
 sg13g2_a22oi_1 _2473_ (.Y(_1890_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .A2(net635),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ));
 sg13g2_a22oi_1 _2474_ (.Y(_1891_),
    .B1(net623),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .A2(net638),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ));
 sg13g2_and2_1 _2475_ (.A(_1890_),
    .B(_1891_),
    .X(_1892_));
 sg13g2_a221oi_1 _2476_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .C1(net621),
    .B1(net629),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .Y(_1893_),
    .A2(net677));
 sg13g2_a22oi_1 _2477_ (.Y(_1894_),
    .B1(net625),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .A2(net633),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ));
 sg13g2_a22oi_1 _2478_ (.Y(_1895_),
    .B1(net619),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .A2(net627),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ));
 sg13g2_and3_1 _2479_ (.X(_1896_),
    .A(_1893_),
    .B(_1894_),
    .C(_1895_));
 sg13g2_a21oi_1 _2480_ (.A1(_1892_),
    .A2(_1896_),
    .Y(_1897_),
    .B1(net565));
 sg13g2_a21oi_1 _2481_ (.A1(_1723_),
    .A2(_1887_),
    .Y(_1898_),
    .B1(_1897_));
 sg13g2_and3_2 _2482_ (.X(_1899_),
    .A(_1888_),
    .B(_1889_),
    .C(_1898_));
 sg13g2_inv_4 _2483_ (.A(_1899_),
    .Y(net22));
 sg13g2_nor2_1 _2484_ (.A(\sap_3_inst.alu.flags[5] ),
    .B(net676),
    .Y(_1900_));
 sg13g2_a21oi_1 _2485_ (.A1(net676),
    .A2(_1899_),
    .Y(_0031_),
    .B1(_1900_));
 sg13g2_a22oi_1 _2486_ (.Y(_1901_),
    .B1(net619),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .A2(net633),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ));
 sg13g2_a22oi_1 _2487_ (.Y(_1902_),
    .B1(net629),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .A2(net631),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ));
 sg13g2_and2_1 _2488_ (.A(_1901_),
    .B(_1902_),
    .X(_1903_));
 sg13g2_a221oi_1 _2489_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .C1(net638),
    .B1(net621),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .Y(_1904_),
    .A2(net623));
 sg13g2_a22oi_1 _2490_ (.Y(_1905_),
    .B1(net627),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .A2(net635),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ));
 sg13g2_a22oi_1 _2491_ (.Y(_1906_),
    .B1(net625),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .A2(net677),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ));
 sg13g2_and3_1 _2492_ (.X(_1907_),
    .A(_1904_),
    .B(_1905_),
    .C(_1906_));
 sg13g2_a22oi_1 _2493_ (.Y(_1908_),
    .B1(_1903_),
    .B2(_1907_),
    .A2(net638),
    .A1(_1468_));
 sg13g2_a22oi_1 _2494_ (.Y(_1909_),
    .B1(_1828_),
    .B2(\sap_3_inst.alu.flags[4] ),
    .A2(_1827_),
    .A1(net751));
 sg13g2_nand2_1 _2495_ (.Y(_1910_),
    .A(net5),
    .B(_1847_));
 sg13g2_a22oi_1 _2496_ (.Y(_1911_),
    .B1(net623),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .A2(net635),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ));
 sg13g2_a22oi_1 _2497_ (.Y(_1912_),
    .B1(net625),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ),
    .A2(net633),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ));
 sg13g2_and2_1 _2498_ (.A(_1911_),
    .B(_1912_),
    .X(_1913_));
 sg13g2_a221oi_1 _2499_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .C1(net621),
    .B1(net638),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ),
    .Y(_1914_),
    .A2(net677));
 sg13g2_a22oi_1 _2500_ (.Y(_1915_),
    .B1(net619),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .A2(net627),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ));
 sg13g2_a22oi_1 _2501_ (.Y(_1916_),
    .B1(net629),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .A2(net631),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ));
 sg13g2_and3_1 _2502_ (.X(_1917_),
    .A(_1914_),
    .B(_1915_),
    .C(_1916_));
 sg13g2_a21oi_1 _2503_ (.A1(_1913_),
    .A2(_1917_),
    .Y(_1918_),
    .B1(net565));
 sg13g2_a21oi_1 _2504_ (.A1(_1723_),
    .A2(_1908_),
    .Y(_1919_),
    .B1(_1918_));
 sg13g2_and3_2 _2505_ (.X(_1920_),
    .A(_1909_),
    .B(_1910_),
    .C(_1919_));
 sg13g2_inv_2 _2506_ (.Y(net21),
    .A(_1920_));
 sg13g2_nor2_1 _2507_ (.A(\sap_3_inst.alu.flags[4] ),
    .B(net676),
    .Y(_1921_));
 sg13g2_a21oi_1 _2508_ (.A1(net676),
    .A2(_1920_),
    .Y(_0030_),
    .B1(_1921_));
 sg13g2_a21oi_1 _2509_ (.A1(_1540_),
    .A2(net688),
    .Y(_1922_),
    .B1(net682));
 sg13g2_nand2_1 _2510_ (.Y(_1923_),
    .A(_1546_),
    .B(net688));
 sg13g2_a21oi_1 _2511_ (.A1(net725),
    .A2(net685),
    .Y(_1924_),
    .B1(_1821_));
 sg13g2_nor2_1 _2512_ (.A(net728),
    .B(_1924_),
    .Y(_1925_));
 sg13g2_inv_1 _2513_ (.Y(_1926_),
    .A(_1925_));
 sg13g2_a21oi_1 _2514_ (.A1(net688),
    .A2(_1568_),
    .Y(_1927_),
    .B1(_1925_));
 sg13g2_o21ai_1 _2515_ (.B1(_1923_),
    .Y(_1928_),
    .A1(net690),
    .A2(_1927_));
 sg13g2_nor3_1 _2516_ (.A(net694),
    .B(_1550_),
    .C(_1716_),
    .Y(_1929_));
 sg13g2_nand2b_1 _2517_ (.Y(_1930_),
    .B(net682),
    .A_N(_1929_));
 sg13g2_a21o_1 _2518_ (.A2(net685),
    .A1(_1549_),
    .B1(_1930_),
    .X(_1931_));
 sg13g2_nand2_1 _2519_ (.Y(_1932_),
    .A(_1559_),
    .B(_1627_));
 sg13g2_a21oi_1 _2520_ (.A1(net706),
    .A2(_1932_),
    .Y(_1933_),
    .B1(_1715_));
 sg13g2_nor2_1 _2521_ (.A(net690),
    .B(_1933_),
    .Y(_1934_));
 sg13g2_nor3_1 _2522_ (.A(_1928_),
    .B(_1931_),
    .C(_1934_),
    .Y(_1935_));
 sg13g2_nor2b_2 _2523_ (.A(_1922_),
    .B_N(_1931_),
    .Y(_1936_));
 sg13g2_inv_1 _2524_ (.Y(_1937_),
    .A(_1936_));
 sg13g2_nor2_1 _2525_ (.A(_1922_),
    .B(_1935_),
    .Y(_1938_));
 sg13g2_o21ai_1 _2526_ (.B1(_1858_),
    .Y(_1939_),
    .A1(_1922_),
    .A2(_1935_));
 sg13g2_inv_2 _2527_ (.Y(_1940_),
    .A(_1939_));
 sg13g2_nand4_1 _2528_ (.B(net725),
    .C(_1508_),
    .A(net729),
    .Y(_1941_),
    .D(net688));
 sg13g2_nand3_1 _2529_ (.B(_1551_),
    .C(_1925_),
    .A(net730),
    .Y(_1942_));
 sg13g2_and2_1 _2530_ (.A(_1941_),
    .B(_1942_),
    .X(_1943_));
 sg13g2_nor3_2 _2531_ (.A(_1521_),
    .B(net695),
    .C(net709),
    .Y(_1944_));
 sg13g2_nand2b_2 _2532_ (.Y(_1945_),
    .B(_1943_),
    .A_N(_1944_));
 sg13g2_nor2_2 _2533_ (.A(_1943_),
    .B(_1944_),
    .Y(_1946_));
 sg13g2_nor2_2 _2534_ (.A(_1550_),
    .B(_1747_),
    .Y(_1947_));
 sg13g2_a21oi_1 _2535_ (.A1(net735),
    .A2(_1928_),
    .Y(_1948_),
    .B1(_1947_));
 sg13g2_o21ai_1 _2536_ (.B1(_1948_),
    .Y(_1949_),
    .A1(_1612_),
    .A2(_1627_));
 sg13g2_and2_1 _2537_ (.A(net732),
    .B(_1928_),
    .X(_1950_));
 sg13g2_nand2_2 _2538_ (.Y(_1951_),
    .A(net732),
    .B(_1928_));
 sg13g2_nand2_1 _2539_ (.Y(_1952_),
    .A(net618),
    .B(_1950_));
 sg13g2_nand2_1 _2540_ (.Y(_1953_),
    .A(_1946_),
    .B(_1952_));
 sg13g2_nand2_1 _2541_ (.Y(_1954_),
    .A(_1945_),
    .B(_1953_));
 sg13g2_a21oi_1 _2542_ (.A1(_1945_),
    .A2(_1953_),
    .Y(_1955_),
    .B1(_1940_));
 sg13g2_a22oi_1 _2543_ (.Y(_1956_),
    .B1(net622),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .A2(net636),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ));
 sg13g2_a22oi_1 _2544_ (.Y(_1957_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .A2(net634),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ));
 sg13g2_and2_1 _2545_ (.A(_1956_),
    .B(_1957_),
    .X(_1958_));
 sg13g2_a221oi_1 _2546_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .C1(net637),
    .B1(net624),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .Y(_1959_),
    .A2(net678));
 sg13g2_a22oi_1 _2547_ (.Y(_1960_),
    .B1(net620),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .A2(net630),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ));
 sg13g2_a22oi_1 _2548_ (.Y(_1961_),
    .B1(net626),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .A2(net628),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ));
 sg13g2_and3_1 _2549_ (.X(_1962_),
    .A(_1959_),
    .B(_1960_),
    .C(_1961_));
 sg13g2_a22oi_1 _2550_ (.Y(_1963_),
    .B1(_1958_),
    .B2(_1962_),
    .A2(net637),
    .A1(_1440_));
 sg13g2_a22oi_1 _2551_ (.Y(_1964_),
    .B1(_1828_),
    .B2(\sap_3_inst.alu.flags[3] ),
    .A2(_1827_),
    .A1(net754));
 sg13g2_nand2_1 _2552_ (.Y(_1965_),
    .A(net4),
    .B(_1847_));
 sg13g2_a22oi_1 _2553_ (.Y(_1966_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .A2(_1794_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ));
 sg13g2_a22oi_1 _2554_ (.Y(_1967_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .A2(net636),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ));
 sg13g2_and2_1 _2555_ (.A(_1966_),
    .B(_1967_),
    .X(_1968_));
 sg13g2_a221oi_1 _2556_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .C1(net622),
    .B1(net624),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .Y(_1969_),
    .A2(net678));
 sg13g2_a22oi_1 _2557_ (.Y(_1970_),
    .B1(net620),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .A2(net630),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ));
 sg13g2_a22oi_1 _2558_ (.Y(_1971_),
    .B1(net626),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .A2(net628),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ));
 sg13g2_and3_1 _2559_ (.X(_1972_),
    .A(_1969_),
    .B(_1970_),
    .C(_1971_));
 sg13g2_a21oi_1 _2560_ (.A1(_1968_),
    .A2(_1972_),
    .Y(_1973_),
    .B1(net566));
 sg13g2_a21oi_1 _2561_ (.A1(_1723_),
    .A2(_1963_),
    .Y(_1974_),
    .B1(_1973_));
 sg13g2_and3_2 _2562_ (.X(_1975_),
    .A(_1964_),
    .B(_1965_),
    .C(_1974_));
 sg13g2_inv_1 _2563_ (.Y(net20),
    .A(net546));
 sg13g2_nor2_1 _2564_ (.A(net743),
    .B(net675),
    .Y(_1976_));
 sg13g2_a21oi_1 _2565_ (.A1(net675),
    .A2(_1975_),
    .Y(_1977_),
    .B1(_1976_));
 sg13g2_mux2_1 _2566_ (.A0(\sap_3_inst.alu.flags[3] ),
    .A1(_1977_),
    .S(_1955_),
    .X(_0029_));
 sg13g2_nand2b_1 _2567_ (.Y(_1978_),
    .B(\sap_3_inst.alu.flags[2] ),
    .A_N(_1955_));
 sg13g2_a22oi_1 _2568_ (.Y(_1979_),
    .B1(net620),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .A2(net626),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ));
 sg13g2_a22oi_1 _2569_ (.Y(_1980_),
    .B1(net632),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .A2(net634),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ));
 sg13g2_a22oi_1 _2570_ (.Y(_1981_),
    .B1(net636),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .A2(net679),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ));
 sg13g2_and2_1 _2571_ (.A(_1979_),
    .B(_1981_),
    .X(_1982_));
 sg13g2_a221oi_1 _2572_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .C1(net637),
    .B1(net622),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .Y(_1983_),
    .A2(net624));
 sg13g2_nand2_1 _2573_ (.Y(_1984_),
    .A(_1980_),
    .B(_1983_));
 sg13g2_a221oi_1 _2574_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .C1(_1984_),
    .B1(net628),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .Y(_1985_),
    .A2(net630));
 sg13g2_a22oi_1 _2575_ (.Y(_1986_),
    .B1(_1982_),
    .B2(_1985_),
    .A2(net637),
    .A1(_1444_));
 sg13g2_and2_1 _2576_ (.A(\sap_3_inst.alu.flags[2] ),
    .B(_1828_),
    .X(_1987_));
 sg13g2_a221oi_1 _2577_ (.B2(net3),
    .C1(_1987_),
    .B1(_1847_),
    .A1(net756),
    .Y(_1988_),
    .A2(_1827_));
 sg13g2_a22oi_1 _2578_ (.Y(_1989_),
    .B1(net634),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .A2(net637),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ));
 sg13g2_a22oi_1 _2579_ (.Y(_1990_),
    .B1(net626),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .A2(net630),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ));
 sg13g2_nand2_1 _2580_ (.Y(_1991_),
    .A(_1989_),
    .B(_1990_));
 sg13g2_a221oi_1 _2581_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .C1(net622),
    .B1(net624),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .Y(_1992_),
    .A2(net679));
 sg13g2_a22oi_1 _2582_ (.Y(_1993_),
    .B1(net628),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ),
    .A2(net636),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ));
 sg13g2_a22oi_1 _2583_ (.Y(_1994_),
    .B1(net620),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ),
    .A2(net632),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ));
 sg13g2_nand3_1 _2584_ (.B(_1993_),
    .C(_1994_),
    .A(_1992_),
    .Y(_1995_));
 sg13g2_nor2_1 _2585_ (.A(_1991_),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_o21ai_1 _2586_ (.B1(_1988_),
    .Y(_1997_),
    .A1(net567),
    .A2(_1996_));
 sg13g2_a21o_2 _2587_ (.A2(_1986_),
    .A1(_1723_),
    .B1(_1997_),
    .X(net545));
 sg13g2_nor2_1 _2588_ (.A(_1858_),
    .B(net545),
    .Y(_1998_));
 sg13g2_xor2_1 _2589_ (.B(net760),
    .A(net757),
    .X(_1999_));
 sg13g2_xor2_1 _2590_ (.B(net756),
    .A(net754),
    .X(_2000_));
 sg13g2_xnor2_1 _2591_ (.Y(_2001_),
    .A(_1999_),
    .B(_2000_));
 sg13g2_xor2_1 _2592_ (.B(net745),
    .A(net743),
    .X(_2002_));
 sg13g2_xor2_1 _2593_ (.B(net751),
    .A(net747),
    .X(_2003_));
 sg13g2_xnor2_1 _2594_ (.Y(_2004_),
    .A(_2002_),
    .B(_2003_));
 sg13g2_xnor2_1 _2595_ (.Y(_2005_),
    .A(_2001_),
    .B(_2004_));
 sg13g2_o21ai_1 _2596_ (.B1(_1955_),
    .Y(_2006_),
    .A1(net675),
    .A2(_2005_));
 sg13g2_o21ai_1 _2597_ (.B1(_1978_),
    .Y(_0028_),
    .A1(_1998_),
    .A2(_2006_));
 sg13g2_or2_1 _2598_ (.X(_2007_),
    .B(_1952_),
    .A(_1945_));
 sg13g2_inv_1 _2599_ (.Y(_2008_),
    .A(net564));
 sg13g2_nand2_2 _2600_ (.Y(_0197_),
    .A(_1946_),
    .B(_1951_));
 sg13g2_nand2_2 _2601_ (.Y(_0198_),
    .A(_1943_),
    .B(_1944_));
 sg13g2_nand3_1 _2602_ (.B(_0197_),
    .C(_0198_),
    .A(net564),
    .Y(_0199_));
 sg13g2_nor2_2 _2603_ (.A(_1936_),
    .B(_1945_),
    .Y(_0200_));
 sg13g2_nor2_2 _2604_ (.A(net618),
    .B(_1951_),
    .Y(_0201_));
 sg13g2_nor2b_2 _2605_ (.A(_1943_),
    .B_N(_1944_),
    .Y(_0202_));
 sg13g2_nor2b_1 _2606_ (.A(_1952_),
    .B_N(_0202_),
    .Y(_0203_));
 sg13g2_nor4_1 _2607_ (.A(_0199_),
    .B(_0200_),
    .C(_0201_),
    .D(_0203_),
    .Y(_0204_));
 sg13g2_o21ai_1 _2608_ (.B1(net720),
    .Y(_0205_),
    .A1(_1940_),
    .A2(_0204_));
 sg13g2_and2_1 _2609_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .B(net624),
    .X(_0206_));
 sg13g2_a22oi_1 _2610_ (.Y(_0207_),
    .B1(net628),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .A2(net632),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ));
 sg13g2_a22oi_1 _2611_ (.Y(_0208_),
    .B1(net620),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .A2(net622),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ));
 sg13g2_a221oi_1 _2612_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .C1(_0206_),
    .B1(net626),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .Y(_0209_),
    .A2(net630));
 sg13g2_a21oi_1 _2613_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .A2(net636),
    .Y(_0210_),
    .B1(net637));
 sg13g2_nand3_1 _2614_ (.B(_0208_),
    .C(_0210_),
    .A(_0207_),
    .Y(_0211_));
 sg13g2_a221oi_1 _2615_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .C1(_0211_),
    .B1(net634),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .Y(_0212_),
    .A2(net679));
 sg13g2_a22oi_1 _2616_ (.Y(_0213_),
    .B1(_0209_),
    .B2(_0212_),
    .A2(net637),
    .A1(_1457_));
 sg13g2_a22oi_1 _2617_ (.Y(_0214_),
    .B1(_1828_),
    .B2(net720),
    .A2(_1827_),
    .A1(net757));
 sg13g2_nand2_1 _2618_ (.Y(_0215_),
    .A(net2),
    .B(_1847_));
 sg13g2_a22oi_1 _2619_ (.Y(_0216_),
    .B1(net620),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .A2(net637),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ));
 sg13g2_a22oi_1 _2620_ (.Y(_0217_),
    .B1(net624),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .A2(net632),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ));
 sg13g2_and2_1 _2621_ (.A(_0216_),
    .B(_0217_),
    .X(_0218_));
 sg13g2_a221oi_1 _2622_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .C1(net622),
    .B1(net634),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ),
    .Y(_0219_),
    .A2(net679));
 sg13g2_a22oi_1 _2623_ (.Y(_0220_),
    .B1(net630),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .A2(net636),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ));
 sg13g2_a22oi_1 _2624_ (.Y(_0221_),
    .B1(net626),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .A2(net628),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ));
 sg13g2_and3_1 _2625_ (.X(_0222_),
    .A(_0219_),
    .B(_0220_),
    .C(_0221_));
 sg13g2_a21oi_1 _2626_ (.A1(_0218_),
    .A2(_0222_),
    .Y(_0223_),
    .B1(net567));
 sg13g2_a21oi_1 _2627_ (.A1(_1723_),
    .A2(_0213_),
    .Y(_0224_),
    .B1(_0223_));
 sg13g2_nand3_1 _2628_ (.B(_0215_),
    .C(_0224_),
    .A(_0214_),
    .Y(net18));
 sg13g2_inv_1 _2629_ (.Y(_0225_),
    .A(net32));
 sg13g2_nor2_1 _2630_ (.A(\sap_3_inst.alu.carry ),
    .B(net675),
    .Y(_0226_));
 sg13g2_nor3_1 _2631_ (.A(_1940_),
    .B(_0204_),
    .C(_0226_),
    .Y(_0227_));
 sg13g2_o21ai_1 _2632_ (.B1(_0227_),
    .Y(_0228_),
    .A1(_1858_),
    .A2(net32));
 sg13g2_nand2_1 _2633_ (.Y(_0027_),
    .A(_0205_),
    .B(_0228_));
 sg13g2_a22oi_1 _2634_ (.Y(_0229_),
    .B1(net629),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .A2(net633),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ));
 sg13g2_a22oi_1 _2635_ (.Y(_0230_),
    .B1(net624),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .A2(net635),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ));
 sg13g2_and2_1 _2636_ (.A(_0229_),
    .B(_0230_),
    .X(_0231_));
 sg13g2_a221oi_1 _2637_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .C1(net639),
    .B1(net622),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .Y(_0232_),
    .A2(net678));
 sg13g2_a22oi_1 _2638_ (.Y(_0233_),
    .B1(net625),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .A2(_1799_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ));
 sg13g2_a22oi_1 _2639_ (.Y(_0234_),
    .B1(net619),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .A2(net632),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ));
 sg13g2_and3_1 _2640_ (.X(_0235_),
    .A(_0232_),
    .B(_0233_),
    .C(_0234_));
 sg13g2_a22oi_1 _2641_ (.Y(_0236_),
    .B1(_0231_),
    .B2(_0235_),
    .A2(net639),
    .A1(_1460_));
 sg13g2_and2_1 _2642_ (.A(_1723_),
    .B(_0236_),
    .X(_0237_));
 sg13g2_a22oi_1 _2643_ (.Y(_0238_),
    .B1(_1828_),
    .B2(\sap_3_inst.alu.flags[0] ),
    .A2(_1827_),
    .A1(net760));
 sg13g2_nand2_1 _2644_ (.Y(_0239_),
    .A(net1),
    .B(_1847_));
 sg13g2_nand2_1 _2645_ (.Y(_0240_),
    .A(_0238_),
    .B(_0239_));
 sg13g2_a22oi_1 _2646_ (.Y(_0241_),
    .B1(_1800_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .A2(_1798_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ));
 sg13g2_a22oi_1 _2647_ (.Y(_0242_),
    .B1(net628),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .A2(net678),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ));
 sg13g2_a22oi_1 _2648_ (.Y(_0243_),
    .B1(net631),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .A2(net639),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ));
 sg13g2_a221oi_1 _2649_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .C1(_1802_),
    .B1(net633),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .Y(_0244_),
    .A2(net635));
 sg13g2_nand3_1 _2650_ (.B(_0242_),
    .C(_0244_),
    .A(_0241_),
    .Y(_0245_));
 sg13g2_a221oi_1 _2651_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .C1(_0245_),
    .B1(net619),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .Y(_0246_),
    .A2(net623));
 sg13g2_a21oi_1 _2652_ (.A1(_0243_),
    .A2(_0246_),
    .Y(_0247_),
    .B1(net566));
 sg13g2_or3_1 _2653_ (.A(_0237_),
    .B(_0240_),
    .C(_0247_),
    .X(net17));
 sg13g2_nor2_1 _2654_ (.A(_1566_),
    .B(_1940_),
    .Y(_0248_));
 sg13g2_nor4_1 _2655_ (.A(net754),
    .B(net744),
    .C(net756),
    .D(net746),
    .Y(_0249_));
 sg13g2_nor4_1 _2656_ (.A(net757),
    .B(net759),
    .C(net749),
    .D(net752),
    .Y(_0250_));
 sg13g2_nand3_1 _2657_ (.B(_0249_),
    .C(_0250_),
    .A(_1954_),
    .Y(_0251_));
 sg13g2_nor4_1 _2658_ (.A(\sap_3_inst.alu.act[1] ),
    .B(\sap_3_inst.alu.act[0] ),
    .C(\sap_3_inst.alu.act[3] ),
    .D(\sap_3_inst.alu.act[2] ),
    .Y(_0252_));
 sg13g2_nor4_1 _2659_ (.A(\sap_3_inst.alu.act[5] ),
    .B(\sap_3_inst.alu.act[4] ),
    .C(\sap_3_inst.alu.act[7] ),
    .D(\sap_3_inst.alu.act[6] ),
    .Y(_0253_));
 sg13g2_nand2_1 _2660_ (.Y(_0254_),
    .A(_0252_),
    .B(_0253_));
 sg13g2_o21ai_1 _2661_ (.B1(_0251_),
    .Y(_0255_),
    .A1(_1954_),
    .A2(_0254_));
 sg13g2_mux2_1 _2662_ (.A0(net31),
    .A1(_0255_),
    .S(_1858_),
    .X(_0256_));
 sg13g2_mux2_1 _2663_ (.A0(\sap_3_inst.alu.flags[0] ),
    .A1(_0256_),
    .S(_0248_),
    .X(_0026_));
 sg13g2_a21oi_1 _2664_ (.A1(_1604_),
    .A2(_1698_),
    .Y(_0257_),
    .B1(_1768_));
 sg13g2_nand4_1 _2665_ (.B(_1699_),
    .C(net682),
    .A(_1686_),
    .Y(_0258_),
    .D(_0257_));
 sg13g2_o21ai_1 _2666_ (.B1(_1823_),
    .Y(_0259_),
    .A1(_1816_),
    .A2(_0258_));
 sg13g2_a21oi_1 _2667_ (.A1(_1812_),
    .A2(_0259_),
    .Y(mem_ram_we),
    .B1(_1526_));
 sg13g2_nand4_1 _2668_ (.B(_1561_),
    .C(_1591_),
    .A(net700),
    .Y(_0260_),
    .D(_1620_));
 sg13g2_o21ai_1 _2669_ (.B1(_1646_),
    .Y(_0261_),
    .A1(_1575_),
    .A2(_1583_));
 sg13g2_a21oi_1 _2670_ (.A1(net673),
    .A2(_0261_),
    .Y(_0262_),
    .B1(net708));
 sg13g2_nand2b_1 _2671_ (.Y(_0263_),
    .B(_1569_),
    .A_N(_1786_));
 sg13g2_nor2_1 _2672_ (.A(_0262_),
    .B(_0263_),
    .Y(_0264_));
 sg13g2_a22oi_1 _2673_ (.Y(_0265_),
    .B1(_1646_),
    .B2(_1592_),
    .A2(_1637_),
    .A1(net707));
 sg13g2_o21ai_1 _2674_ (.B1(_1626_),
    .Y(_0266_),
    .A1(_1589_),
    .A2(_1596_));
 sg13g2_nand4_1 _2675_ (.B(_1750_),
    .C(_0265_),
    .A(_1659_),
    .Y(_0267_),
    .D(_0266_));
 sg13g2_o21ai_1 _2676_ (.B1(_1587_),
    .Y(_0268_),
    .A1(net696),
    .A2(_1646_));
 sg13g2_o21ai_1 _2677_ (.B1(_1599_),
    .Y(_0269_),
    .A1(net696),
    .A2(_1626_));
 sg13g2_o21ai_1 _2678_ (.B1(_1605_),
    .Y(_0270_),
    .A1(net696),
    .A2(_1637_));
 sg13g2_nand3_1 _2679_ (.B(_0269_),
    .C(_0270_),
    .A(_0268_),
    .Y(_0271_));
 sg13g2_a21oi_1 _2680_ (.A1(_1623_),
    .A2(_0271_),
    .Y(_0272_),
    .B1(_0267_));
 sg13g2_a21oi_2 _2681_ (.B1(_1606_),
    .Y(_0273_),
    .A2(_1622_),
    .A1(net700));
 sg13g2_nand3_1 _2682_ (.B(_0264_),
    .C(_0272_),
    .A(_1815_),
    .Y(_0274_));
 sg13g2_a221oi_1 _2683_ (.B2(_1555_),
    .C1(_1569_),
    .B1(_1690_),
    .A1(net688),
    .Y(_0275_),
    .A2(_1568_));
 sg13g2_a21oi_1 _2684_ (.A1(_1926_),
    .A2(_0275_),
    .Y(_0276_),
    .B1(net690));
 sg13g2_a221oi_1 _2685_ (.B2(_0276_),
    .C1(_1930_),
    .B1(_0274_),
    .A1(net690),
    .Y(_0277_),
    .A2(net688));
 sg13g2_a21oi_1 _2686_ (.A1(net698),
    .A2(_1713_),
    .Y(_0278_),
    .B1(_1823_));
 sg13g2_nor4_1 _2687_ (.A(net713),
    .B(net712),
    .C(_0277_),
    .D(_0278_),
    .Y(_0279_));
 sg13g2_a21oi_1 _2688_ (.A1(net703),
    .A2(_1515_),
    .Y(_0280_),
    .B1(_1675_));
 sg13g2_nor3_1 _2689_ (.A(_1526_),
    .B(_0279_),
    .C(_0280_),
    .Y(_0281_));
 sg13g2_a221oi_1 _2690_ (.B2(_1499_),
    .C1(_0281_),
    .B1(_1528_),
    .A1(_1508_),
    .Y(_0282_),
    .A2(net712));
 sg13g2_nor2_1 _2691_ (.A(net719),
    .B(_0282_),
    .Y(_0002_));
 sg13g2_nor2_1 _2692_ (.A(_1535_),
    .B(_0282_),
    .Y(_0003_));
 sg13g2_nor3_1 _2693_ (.A(_1635_),
    .B(_1744_),
    .C(_0282_),
    .Y(_0004_));
 sg13g2_nor2_1 _2694_ (.A(net716),
    .B(_1635_),
    .Y(_0283_));
 sg13g2_nor3_1 _2695_ (.A(_1637_),
    .B(_0282_),
    .C(_0283_),
    .Y(_0005_));
 sg13g2_nor2b_2 _2696_ (.A(net566),
    .B_N(_0236_),
    .Y(net9));
 sg13g2_nor2b_2 _2697_ (.A(net567),
    .B_N(_0213_),
    .Y(net10));
 sg13g2_nor2b_2 _2698_ (.A(net567),
    .B_N(_1986_),
    .Y(net11));
 sg13g2_nor2b_2 _2699_ (.A(net566),
    .B_N(_1963_),
    .Y(net12));
 sg13g2_nor2b_2 _2700_ (.A(net565),
    .B_N(_1908_),
    .Y(net13));
 sg13g2_nor2b_2 _2701_ (.A(net565),
    .B_N(_1887_),
    .Y(net14));
 sg13g2_nor2b_2 _2702_ (.A(net565),
    .B_N(_1866_),
    .Y(net15));
 sg13g2_nor2b_2 _2703_ (.A(net565),
    .B_N(_1810_),
    .Y(net16));
 sg13g2_nand3_1 _2704_ (.B(_1514_),
    .C(net699),
    .A(_1508_),
    .Y(_0001_));
 sg13g2_nor2_1 _2705_ (.A(net707),
    .B(_1628_),
    .Y(_0284_));
 sg13g2_a21oi_1 _2706_ (.A1(_1616_),
    .A2(_0284_),
    .Y(_0285_),
    .B1(net696));
 sg13g2_nand2_1 _2707_ (.Y(_0286_),
    .A(_1653_),
    .B(_0285_));
 sg13g2_a221oi_1 _2708_ (.B2(_1655_),
    .C1(net681),
    .B1(net687),
    .A1(net700),
    .Y(_0287_),
    .A2(_1553_));
 sg13g2_nand3_1 _2709_ (.B(_1578_),
    .C(_1642_),
    .A(net694),
    .Y(_0288_));
 sg13g2_nand4_1 _2710_ (.B(_1593_),
    .C(_1597_),
    .A(_1590_),
    .Y(_0289_),
    .D(_1708_));
 sg13g2_a22oi_1 _2711_ (.Y(_0290_),
    .B1(_0288_),
    .B2(_1709_),
    .A2(_0286_),
    .A1(_1677_));
 sg13g2_nand3_1 _2712_ (.B(_1602_),
    .C(_0289_),
    .A(_1580_),
    .Y(_0291_));
 sg13g2_nand3_1 _2713_ (.B(_0290_),
    .C(_0291_),
    .A(_0287_),
    .Y(_0292_));
 sg13g2_nand2_1 _2714_ (.Y(_0293_),
    .A(_1619_),
    .B(_0292_));
 sg13g2_a21oi_1 _2715_ (.A1(_1569_),
    .A2(_0293_),
    .Y(_0294_),
    .B1(_1572_));
 sg13g2_o21ai_1 _2716_ (.B1(_1538_),
    .Y(_0295_),
    .A1(_1548_),
    .A2(_0294_));
 sg13g2_nand2_1 _2717_ (.Y(_0296_),
    .A(net703),
    .B(_0295_));
 sg13g2_nand2_1 _2718_ (.Y(_0297_),
    .A(_1537_),
    .B(_0296_));
 sg13g2_nand2_1 _2719_ (.Y(mem_mar_we),
    .A(_1503_),
    .B(_0297_));
 sg13g2_nor2_2 _2720_ (.A(\u_ser.state[0] ),
    .B(\u_ser.state[1] ),
    .Y(_0186_));
 sg13g2_mux2_1 _2721_ (.A0(net70),
    .A1(\sap_3_inst.out[0] ),
    .S(net766),
    .X(_0018_));
 sg13g2_mux2_1 _2722_ (.A0(net61),
    .A1(\sap_3_inst.out[1] ),
    .S(net766),
    .X(_0019_));
 sg13g2_mux2_1 _2723_ (.A0(net62),
    .A1(\sap_3_inst.out[2] ),
    .S(net766),
    .X(_0020_));
 sg13g2_mux2_1 _2724_ (.A0(net57),
    .A1(\sap_3_inst.out[3] ),
    .S(net766),
    .X(_0021_));
 sg13g2_mux2_1 _2725_ (.A0(net74),
    .A1(\sap_3_inst.out[4] ),
    .S(net766),
    .X(_0022_));
 sg13g2_mux2_1 _2726_ (.A0(net65),
    .A1(\sap_3_inst.out[5] ),
    .S(net766),
    .X(_0023_));
 sg13g2_mux2_1 _2727_ (.A0(net56),
    .A1(\sap_3_inst.out[6] ),
    .S(_0186_),
    .X(_0024_));
 sg13g2_mux2_1 _2728_ (.A0(net60),
    .A1(\sap_3_inst.out[7] ),
    .S(_0186_),
    .X(_0025_));
 sg13g2_nand3_1 _2729_ (.B(_1504_),
    .C(net713),
    .A(net733),
    .Y(_0298_));
 sg13g2_nor2_1 _2730_ (.A(_1546_),
    .B(_1718_),
    .Y(_0299_));
 sg13g2_nand2b_1 _2731_ (.Y(_0300_),
    .B(_1839_),
    .A_N(_1716_));
 sg13g2_nand2_1 _2732_ (.Y(_0301_),
    .A(_1551_),
    .B(_1757_));
 sg13g2_o21ai_1 _2733_ (.B1(_1612_),
    .Y(_0302_),
    .A1(net723),
    .A2(_1576_));
 sg13g2_a21oi_1 _2734_ (.A1(_1690_),
    .A2(_0302_),
    .Y(_0303_),
    .B1(_1837_));
 sg13g2_nor2b_1 _2735_ (.A(_0301_),
    .B_N(_1832_),
    .Y(_0304_));
 sg13g2_nand3_1 _2736_ (.B(_0303_),
    .C(_0304_),
    .A(_0300_),
    .Y(_0305_));
 sg13g2_a21oi_1 _2737_ (.A1(_0299_),
    .A2(_0305_),
    .Y(_0306_),
    .B1(_1715_));
 sg13g2_nor3_1 _2738_ (.A(_1511_),
    .B(net695),
    .C(_1716_),
    .Y(_0307_));
 sg13g2_nor3_1 _2739_ (.A(net683),
    .B(_1845_),
    .C(_0307_),
    .Y(_0308_));
 sg13g2_or3_1 _2740_ (.A(net713),
    .B(_0306_),
    .C(_0308_),
    .X(_0309_));
 sg13g2_o21ai_1 _2741_ (.B1(_0309_),
    .Y(_0310_),
    .A1(_1675_),
    .A2(_0298_));
 sg13g2_or2_1 _2742_ (.X(_0311_),
    .B(net617),
    .A(_1938_));
 sg13g2_a21oi_1 _2743_ (.A1(_1611_),
    .A2(_1639_),
    .Y(_0312_),
    .B1(net689));
 sg13g2_o21ai_1 _2744_ (.B1(net683),
    .Y(_0313_),
    .A1(_1551_),
    .A2(_1814_));
 sg13g2_o21ai_1 _2745_ (.B1(_1822_),
    .Y(_0314_),
    .A1(_0312_),
    .A2(_0313_));
 sg13g2_nand3_1 _2746_ (.B(net618),
    .C(_1950_),
    .A(_1946_),
    .Y(_0315_));
 sg13g2_and2_1 _2747_ (.A(net618),
    .B(_1951_),
    .X(_0316_));
 sg13g2_nand2b_1 _2748_ (.Y(_0317_),
    .B(_0202_),
    .A_N(_0316_));
 sg13g2_o21ai_1 _2749_ (.B1(_0315_),
    .Y(_0318_),
    .A1(_0311_),
    .A2(net670));
 sg13g2_nand2b_1 _2750_ (.Y(_0319_),
    .B(_0317_),
    .A_N(_0318_));
 sg13g2_nand2_1 _2751_ (.Y(_0320_),
    .A(net759),
    .B(\sap_3_inst.alu.tmp[0] ));
 sg13g2_xor2_1 _2752_ (.B(\sap_3_inst.alu.tmp[0] ),
    .A(net759),
    .X(_0321_));
 sg13g2_and2_1 _2753_ (.A(_0200_),
    .B(_0201_),
    .X(_0322_));
 sg13g2_nand2_2 _2754_ (.Y(_0323_),
    .A(_0200_),
    .B(_0201_));
 sg13g2_and2_1 _2755_ (.A(_0200_),
    .B(_0316_),
    .X(_0324_));
 sg13g2_nand2_1 _2756_ (.Y(_0325_),
    .A(_0200_),
    .B(_0316_));
 sg13g2_nor2_1 _2757_ (.A(_0322_),
    .B(_0324_),
    .Y(_0326_));
 sg13g2_nand2_2 _2758_ (.Y(_0327_),
    .A(_0202_),
    .B(_0316_));
 sg13g2_a21oi_1 _2759_ (.A1(_0202_),
    .A2(_0316_),
    .Y(_0328_),
    .B1(_1936_));
 sg13g2_nand2_1 _2760_ (.Y(_0329_),
    .A(_0326_),
    .B(_0328_));
 sg13g2_and2_1 _2761_ (.A(_1946_),
    .B(_0201_),
    .X(_0330_));
 sg13g2_nor3_1 _2762_ (.A(_0199_),
    .B(_0329_),
    .C(net563),
    .Y(_0331_));
 sg13g2_inv_1 _2763_ (.Y(_0332_),
    .A(net543));
 sg13g2_nor2b_2 _2764_ (.A(_0197_),
    .B_N(net618),
    .Y(_0333_));
 sg13g2_or2_1 _2765_ (.X(_0334_),
    .B(_0333_),
    .A(_0322_));
 sg13g2_o21ai_1 _2766_ (.B1(_0321_),
    .Y(_0335_),
    .A1(net544),
    .A2(_0334_));
 sg13g2_o21ai_1 _2767_ (.B1(net563),
    .Y(_0336_),
    .A1(net759),
    .A2(\sap_3_inst.alu.tmp[0] ));
 sg13g2_and2_1 _2768_ (.A(net720),
    .B(_1950_),
    .X(_0337_));
 sg13g2_nor2_1 _2769_ (.A(_1949_),
    .B(_0198_),
    .Y(_0338_));
 sg13g2_nor2b_2 _2770_ (.A(_0198_),
    .B_N(_1949_),
    .Y(_0339_));
 sg13g2_nor2_2 _2771_ (.A(_1949_),
    .B(_0197_),
    .Y(_0340_));
 sg13g2_nand2b_1 _2772_ (.Y(_0341_),
    .B(_0340_),
    .A_N(_0320_));
 sg13g2_nor2_1 _2773_ (.A(net760),
    .B(_0328_),
    .Y(_0342_));
 sg13g2_nand2b_1 _2774_ (.Y(_0343_),
    .B(net720),
    .A_N(_0321_));
 sg13g2_nand2b_1 _2775_ (.Y(_0344_),
    .B(_0321_),
    .A_N(net720));
 sg13g2_nand2_1 _2776_ (.Y(_0345_),
    .A(net720),
    .B(_0321_));
 sg13g2_a22oi_1 _2777_ (.Y(_0346_),
    .B1(_0343_),
    .B2(_0344_),
    .A2(_0325_),
    .A1(net564));
 sg13g2_a221oi_1 _2778_ (.B2(net757),
    .C1(net670),
    .B1(net572),
    .A1(_0337_),
    .Y(_0347_),
    .A2(net573));
 sg13g2_nand2_1 _2779_ (.Y(_0348_),
    .A(_0336_),
    .B(_0341_));
 sg13g2_nor3_1 _2780_ (.A(_0342_),
    .B(_0346_),
    .C(_0348_),
    .Y(_0349_));
 sg13g2_nand3_1 _2781_ (.B(_0347_),
    .C(_0349_),
    .A(_0335_),
    .Y(_0350_));
 sg13g2_a21oi_1 _2782_ (.A1(_1462_),
    .A2(net670),
    .Y(_0351_),
    .B1(net617));
 sg13g2_a221oi_1 _2783_ (.B2(_0351_),
    .C1(net555),
    .B1(_0350_),
    .A1(net31),
    .Y(_0352_),
    .A2(net617));
 sg13g2_a21oi_1 _2784_ (.A1(_1456_),
    .A2(net555),
    .Y(_0034_),
    .B1(_0352_));
 sg13g2_nand2_1 _2785_ (.Y(_0353_),
    .A(net757),
    .B(\sap_3_inst.alu.tmp[1] ));
 sg13g2_nand2_1 _2786_ (.Y(_0354_),
    .A(_1455_),
    .B(_1463_));
 sg13g2_xor2_1 _2787_ (.B(\sap_3_inst.alu.tmp[1] ),
    .A(net758),
    .X(_0355_));
 sg13g2_nand2b_1 _2788_ (.Y(_0356_),
    .B(\sap_3_inst.alu.tmp[0] ),
    .A_N(net759));
 sg13g2_nor2b_1 _2789_ (.A(_0355_),
    .B_N(_0356_),
    .Y(_0357_));
 sg13g2_xnor2_1 _2790_ (.Y(_0358_),
    .A(_0355_),
    .B(_0356_));
 sg13g2_nor2_1 _2791_ (.A(_0343_),
    .B(_0358_),
    .Y(_0359_));
 sg13g2_and2_1 _2792_ (.A(_0343_),
    .B(_0358_),
    .X(_0360_));
 sg13g2_o21ai_1 _2793_ (.B1(_2008_),
    .Y(_0361_),
    .A1(_0359_),
    .A2(_0360_));
 sg13g2_o21ai_1 _2794_ (.B1(_0361_),
    .Y(_0362_),
    .A1(net757),
    .A2(_0327_));
 sg13g2_a221oi_1 _2795_ (.B2(_0322_),
    .C1(_0362_),
    .B1(_0358_),
    .A1(net563),
    .Y(_0363_),
    .A2(_0354_));
 sg13g2_nor3_1 _2796_ (.A(net618),
    .B(_0197_),
    .C(_0353_),
    .Y(_0364_));
 sg13g2_a221oi_1 _2797_ (.B2(_0333_),
    .C1(_0364_),
    .B1(_0355_),
    .A1(net759),
    .Y(_0365_),
    .A2(net573));
 sg13g2_nand3_1 _2798_ (.B(_0321_),
    .C(_0355_),
    .A(net720),
    .Y(_0366_));
 sg13g2_nand2b_1 _2799_ (.Y(_0367_),
    .B(_0355_),
    .A_N(_0320_));
 sg13g2_xor2_1 _2800_ (.B(_0355_),
    .A(_0320_),
    .X(_0368_));
 sg13g2_a21oi_1 _2801_ (.A1(_0345_),
    .A2(_0368_),
    .Y(_0369_),
    .B1(_0325_));
 sg13g2_nor3_1 _2802_ (.A(_1455_),
    .B(_1550_),
    .C(_1747_),
    .Y(_0370_));
 sg13g2_o21ai_1 _2803_ (.B1(_1455_),
    .Y(_0371_),
    .A1(_1550_),
    .A2(_1747_));
 sg13g2_nor2b_1 _2804_ (.A(_0370_),
    .B_N(_0371_),
    .Y(_0372_));
 sg13g2_o21ai_1 _2805_ (.B1(_1936_),
    .Y(_0373_),
    .A1(net760),
    .A2(_0372_));
 sg13g2_a21oi_1 _2806_ (.A1(net759),
    .A2(_0372_),
    .Y(_0374_),
    .B1(_0373_));
 sg13g2_a221oi_1 _2807_ (.B2(_0369_),
    .C1(_0374_),
    .B1(_0366_),
    .A1(net756),
    .Y(_0375_),
    .A2(net572));
 sg13g2_nand3_1 _2808_ (.B(_0365_),
    .C(_0375_),
    .A(_0363_),
    .Y(_0376_));
 sg13g2_a21oi_1 _2809_ (.A1(net544),
    .A2(_0368_),
    .Y(_0377_),
    .B1(net670));
 sg13g2_o21ai_1 _2810_ (.B1(_0377_),
    .Y(_0378_),
    .A1(net544),
    .A2(_0376_));
 sg13g2_a21oi_1 _2811_ (.A1(\sap_3_inst.alu.act[1] ),
    .A2(net670),
    .Y(_0379_),
    .B1(net617));
 sg13g2_a221oi_1 _2812_ (.B2(_0379_),
    .C1(net555),
    .B1(_0378_),
    .A1(_0225_),
    .Y(_0380_),
    .A2(net617));
 sg13g2_a21o_1 _2813_ (.A2(net555),
    .A1(net757),
    .B1(_0380_),
    .X(_0035_));
 sg13g2_nor2b_1 _2814_ (.A(net545),
    .B_N(net616),
    .Y(_0381_));
 sg13g2_xnor2_1 _2815_ (.Y(_0382_),
    .A(net755),
    .B(\sap_3_inst.alu.tmp[2] ));
 sg13g2_inv_1 _2816_ (.Y(_0383_),
    .A(_0382_));
 sg13g2_a21oi_1 _2817_ (.A1(_0353_),
    .A2(_0367_),
    .Y(_0384_),
    .B1(_0382_));
 sg13g2_nand3_1 _2818_ (.B(_0367_),
    .C(_0382_),
    .A(_0353_),
    .Y(_0385_));
 sg13g2_nor2b_1 _2819_ (.A(_0384_),
    .B_N(_0385_),
    .Y(_0386_));
 sg13g2_inv_1 _2820_ (.Y(_0387_),
    .A(_0386_));
 sg13g2_xnor2_1 _2821_ (.Y(_0388_),
    .A(_0366_),
    .B(_0386_));
 sg13g2_a21oi_1 _2822_ (.A1(net758),
    .A2(_1463_),
    .Y(_0389_),
    .B1(_0357_));
 sg13g2_nor2_1 _2823_ (.A(_0383_),
    .B(_0389_),
    .Y(_0390_));
 sg13g2_xnor2_1 _2824_ (.Y(_0391_),
    .A(_0382_),
    .B(_0389_));
 sg13g2_nand2b_1 _2825_ (.Y(_0392_),
    .B(_0359_),
    .A_N(_0391_));
 sg13g2_xor2_1 _2826_ (.B(_0391_),
    .A(_0359_),
    .X(_0393_));
 sg13g2_o21ai_1 _2827_ (.B1(net563),
    .Y(_0394_),
    .A1(net755),
    .A2(\sap_3_inst.alu.tmp[2] ));
 sg13g2_o21ai_1 _2828_ (.B1(_0394_),
    .Y(_0395_),
    .A1(net755),
    .A2(_0327_));
 sg13g2_a221oi_1 _2829_ (.B2(_2008_),
    .C1(_0395_),
    .B1(_0393_),
    .A1(_0324_),
    .Y(_0396_),
    .A2(_0388_));
 sg13g2_and3_1 _2830_ (.X(_0397_),
    .A(net755),
    .B(\sap_3_inst.alu.tmp[2] ),
    .C(_0340_));
 sg13g2_a221oi_1 _2831_ (.B2(_0333_),
    .C1(_0397_),
    .B1(_0383_),
    .A1(net753),
    .Y(_0398_),
    .A2(net572));
 sg13g2_nand2_1 _2832_ (.Y(_0399_),
    .A(net756),
    .B(net672));
 sg13g2_xnor2_1 _2833_ (.Y(_0400_),
    .A(net756),
    .B(_1947_));
 sg13g2_a21oi_1 _2834_ (.A1(net760),
    .A2(_0371_),
    .Y(_0401_),
    .B1(_0370_));
 sg13g2_nand2_1 _2835_ (.Y(_0402_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_or2_1 _2836_ (.X(_0403_),
    .B(_0401_),
    .A(_0400_));
 sg13g2_and3_1 _2837_ (.X(_0404_),
    .A(_1936_),
    .B(_0402_),
    .C(_0403_));
 sg13g2_a221oi_1 _2838_ (.B2(_0322_),
    .C1(_0404_),
    .B1(_0391_),
    .A1(net758),
    .Y(_0405_),
    .A2(net573));
 sg13g2_nand4_1 _2839_ (.B(_0396_),
    .C(_0398_),
    .A(_0332_),
    .Y(_0406_),
    .D(_0405_));
 sg13g2_a21oi_1 _2840_ (.A1(net543),
    .A2(_0387_),
    .Y(_0407_),
    .B1(net669));
 sg13g2_a221oi_1 _2841_ (.B2(_0407_),
    .C1(net616),
    .B1(_0406_),
    .A1(\sap_3_inst.alu.act[2] ),
    .Y(_0408_),
    .A2(net669));
 sg13g2_nor3_1 _2842_ (.A(net554),
    .B(_0381_),
    .C(_0408_),
    .Y(_0409_));
 sg13g2_a21o_1 _2843_ (.A2(net554),
    .A1(\sap_3_inst.alu.acc[2] ),
    .B1(_0409_),
    .X(_0036_));
 sg13g2_nand2_1 _2844_ (.Y(_0410_),
    .A(_0399_),
    .B(_0403_));
 sg13g2_nor2_1 _2845_ (.A(net754),
    .B(net672),
    .Y(_0411_));
 sg13g2_xnor2_1 _2846_ (.Y(_0412_),
    .A(net753),
    .B(net672));
 sg13g2_a21oi_1 _2847_ (.A1(_0399_),
    .A2(_0403_),
    .Y(_0413_),
    .B1(_0411_));
 sg13g2_xnor2_1 _2848_ (.Y(_0414_),
    .A(_0410_),
    .B(_0412_));
 sg13g2_and2_1 _2849_ (.A(net753),
    .B(\sap_3_inst.alu.tmp[3] ),
    .X(_0415_));
 sg13g2_nand2_1 _2850_ (.Y(_0416_),
    .A(net753),
    .B(\sap_3_inst.alu.tmp[3] ));
 sg13g2_nor2_1 _2851_ (.A(net753),
    .B(\sap_3_inst.alu.tmp[3] ),
    .Y(_0417_));
 sg13g2_a21oi_1 _2852_ (.A1(_0333_),
    .A2(_0416_),
    .Y(_0418_),
    .B1(net563));
 sg13g2_a22oi_1 _2853_ (.Y(_0419_),
    .B1(_0340_),
    .B2(_0415_),
    .A2(net573),
    .A1(net755));
 sg13g2_o21ai_1 _2854_ (.B1(_0419_),
    .Y(_0420_),
    .A1(_0417_),
    .A2(_0418_));
 sg13g2_a221oi_1 _2855_ (.B2(_1936_),
    .C1(_0420_),
    .B1(_0414_),
    .A1(net752),
    .Y(_0421_),
    .A2(net572));
 sg13g2_or2_1 _2856_ (.X(_0422_),
    .B(_0417_),
    .A(_0415_));
 sg13g2_inv_1 _2857_ (.Y(_0423_),
    .A(_0422_));
 sg13g2_a21oi_1 _2858_ (.A1(net755),
    .A2(\sap_3_inst.alu.tmp[2] ),
    .Y(_0424_),
    .B1(_0384_));
 sg13g2_xnor2_1 _2859_ (.Y(_0425_),
    .A(_0422_),
    .B(_0424_));
 sg13g2_or3_1 _2860_ (.A(_0366_),
    .B(_0387_),
    .C(_0425_),
    .X(_0426_));
 sg13g2_o21ai_1 _2861_ (.B1(_0425_),
    .Y(_0427_),
    .A1(_0366_),
    .A2(_0387_));
 sg13g2_nand3_1 _2862_ (.B(_0426_),
    .C(_0427_),
    .A(_0324_),
    .Y(_0428_));
 sg13g2_a21oi_1 _2863_ (.A1(net755),
    .A2(_1464_),
    .Y(_0429_),
    .B1(_0390_));
 sg13g2_nor2_1 _2864_ (.A(_0423_),
    .B(_0429_),
    .Y(_0430_));
 sg13g2_xnor2_1 _2865_ (.Y(_0431_),
    .A(_0423_),
    .B(_0429_));
 sg13g2_nand2b_2 _2866_ (.Y(_0432_),
    .B(_0431_),
    .A_N(_0392_));
 sg13g2_xnor2_1 _2867_ (.Y(_0433_),
    .A(_0392_),
    .B(_0431_));
 sg13g2_o21ai_1 _2868_ (.B1(_0428_),
    .Y(_0434_),
    .A1(net564),
    .A2(_0433_));
 sg13g2_nor2_1 _2869_ (.A(_0323_),
    .B(_0431_),
    .Y(_0435_));
 sg13g2_nor2_1 _2870_ (.A(net753),
    .B(_0327_),
    .Y(_0436_));
 sg13g2_nor4_1 _2871_ (.A(net543),
    .B(_0434_),
    .C(_0435_),
    .D(_0436_),
    .Y(_0437_));
 sg13g2_a221oi_1 _2872_ (.B2(_0421_),
    .C1(net669),
    .B1(_0437_),
    .A1(net543),
    .Y(_0438_),
    .A2(_0425_));
 sg13g2_inv_1 _2873_ (.Y(_0439_),
    .A(_0438_));
 sg13g2_a21oi_1 _2874_ (.A1(\sap_3_inst.alu.act[3] ),
    .A2(net669),
    .Y(_0440_),
    .B1(net616));
 sg13g2_a221oi_1 _2875_ (.B2(_0440_),
    .C1(net554),
    .B1(_0439_),
    .A1(net546),
    .Y(_0441_),
    .A2(net616));
 sg13g2_a21o_1 _2876_ (.A2(net554),
    .A1(net753),
    .B1(_0441_),
    .X(_0037_));
 sg13g2_xnor2_1 _2877_ (.Y(_0442_),
    .A(net751),
    .B(net671));
 sg13g2_a21oi_1 _2878_ (.A1(net754),
    .A2(net671),
    .Y(_0443_),
    .B1(_0413_));
 sg13g2_nor2_1 _2879_ (.A(_0442_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_a21o_1 _2880_ (.A2(_0443_),
    .A1(_0442_),
    .B1(_1937_),
    .X(_0445_));
 sg13g2_and3_1 _2881_ (.X(_0446_),
    .A(net750),
    .B(\sap_3_inst.alu.tmp[4] ),
    .C(_0340_));
 sg13g2_xor2_1 _2882_ (.B(\sap_3_inst.alu.tmp[4] ),
    .A(net750),
    .X(_0447_));
 sg13g2_a21oi_1 _2883_ (.A1(_0416_),
    .A2(_0424_),
    .Y(_0448_),
    .B1(_0417_));
 sg13g2_and2_1 _2884_ (.A(_0447_),
    .B(_0448_),
    .X(_0449_));
 sg13g2_xnor2_1 _2885_ (.Y(_0450_),
    .A(_0447_),
    .B(_0448_));
 sg13g2_nand2_1 _2886_ (.Y(_0451_),
    .A(_0426_),
    .B(_0450_));
 sg13g2_nor2_1 _2887_ (.A(_0426_),
    .B(_0450_),
    .Y(_0452_));
 sg13g2_nand3b_1 _2888_ (.B(_0324_),
    .C(_0451_),
    .Y(_0453_),
    .A_N(_0452_));
 sg13g2_o21ai_1 _2889_ (.B1(_0453_),
    .Y(_0454_),
    .A1(net750),
    .A2(_0327_));
 sg13g2_o21ai_1 _2890_ (.B1(net563),
    .Y(_0455_),
    .A1(net750),
    .A2(\sap_3_inst.alu.tmp[4] ));
 sg13g2_a21oi_1 _2891_ (.A1(net754),
    .A2(_1465_),
    .Y(_0456_),
    .B1(_0430_));
 sg13g2_or2_1 _2892_ (.X(_0457_),
    .B(_0456_),
    .A(_0447_));
 sg13g2_xor2_1 _2893_ (.B(_0456_),
    .A(_0447_),
    .X(_0458_));
 sg13g2_nor2_1 _2894_ (.A(_0432_),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_a22oi_1 _2895_ (.Y(_0460_),
    .B1(_0458_),
    .B2(_0322_),
    .A2(net572),
    .A1(net749));
 sg13g2_a221oi_1 _2896_ (.B2(_0333_),
    .C1(_0446_),
    .B1(_0447_),
    .A1(\sap_3_inst.alu.acc[3] ),
    .Y(_0461_),
    .A2(net573));
 sg13g2_nand2_1 _2897_ (.Y(_0462_),
    .A(_0460_),
    .B(_0461_));
 sg13g2_xor2_1 _2898_ (.B(_0458_),
    .A(_0432_),
    .X(_0463_));
 sg13g2_o21ai_1 _2899_ (.B1(_0455_),
    .Y(_0464_),
    .A1(net564),
    .A2(_0463_));
 sg13g2_nor4_1 _2900_ (.A(net543),
    .B(_0454_),
    .C(_0462_),
    .D(_0464_),
    .Y(_0465_));
 sg13g2_o21ai_1 _2901_ (.B1(_0465_),
    .Y(_0466_),
    .A1(_0444_),
    .A2(_0445_));
 sg13g2_a21oi_1 _2902_ (.A1(net544),
    .A2(_0450_),
    .Y(_0467_),
    .B1(_0314_));
 sg13g2_nand2_1 _2903_ (.Y(_0468_),
    .A(_0466_),
    .B(_0467_));
 sg13g2_a21oi_1 _2904_ (.A1(\sap_3_inst.alu.act[4] ),
    .A2(net669),
    .Y(_0469_),
    .B1(net616));
 sg13g2_a221oi_1 _2905_ (.B2(_0469_),
    .C1(net554),
    .B1(_0468_),
    .A1(_1920_),
    .Y(_0470_),
    .A2(net616));
 sg13g2_a21o_1 _2906_ (.A2(net554),
    .A1(net751),
    .B1(_0470_),
    .X(_0038_));
 sg13g2_a21o_1 _2907_ (.A2(net671),
    .A1(net751),
    .B1(_0444_),
    .X(_0471_));
 sg13g2_nand2_1 _2908_ (.Y(_0472_),
    .A(net747),
    .B(net671));
 sg13g2_xor2_1 _2909_ (.B(net671),
    .A(net747),
    .X(_0473_));
 sg13g2_a21oi_1 _2910_ (.A1(_0471_),
    .A2(_0473_),
    .Y(_0474_),
    .B1(_1937_));
 sg13g2_o21ai_1 _2911_ (.B1(_0474_),
    .Y(_0475_),
    .A1(_0471_),
    .A2(_0473_));
 sg13g2_a22oi_1 _2912_ (.Y(_0476_),
    .B1(_0339_),
    .B2(net746),
    .A2(_0338_),
    .A1(net752));
 sg13g2_and2_1 _2913_ (.A(net747),
    .B(\sap_3_inst.alu.tmp[5] ),
    .X(_0477_));
 sg13g2_or2_1 _2914_ (.X(_0478_),
    .B(\sap_3_inst.alu.tmp[5] ),
    .A(net747));
 sg13g2_nor2b_2 _2915_ (.A(_0477_),
    .B_N(_0478_),
    .Y(_0479_));
 sg13g2_a22oi_1 _2916_ (.Y(_0480_),
    .B1(_0479_),
    .B2(_0333_),
    .A2(_0477_),
    .A1(_0340_));
 sg13g2_nand2_1 _2917_ (.Y(_0481_),
    .A(_0476_),
    .B(_0480_));
 sg13g2_nor3_1 _2918_ (.A(_0432_),
    .B(_0447_),
    .C(_0479_),
    .Y(_0482_));
 sg13g2_a22oi_1 _2919_ (.Y(_0483_),
    .B1(_0482_),
    .B2(_2008_),
    .A2(_0478_),
    .A1(net563));
 sg13g2_o21ai_1 _2920_ (.B1(_0483_),
    .Y(_0484_),
    .A1(net748),
    .A2(_0327_));
 sg13g2_nand2b_1 _2921_ (.Y(_0485_),
    .B(net750),
    .A_N(\sap_3_inst.alu.tmp[4] ));
 sg13g2_and3_1 _2922_ (.X(_0486_),
    .A(_0457_),
    .B(_0479_),
    .C(_0485_));
 sg13g2_a21oi_1 _2923_ (.A1(_0457_),
    .A2(_0485_),
    .Y(_0487_),
    .B1(_0479_));
 sg13g2_nor2_1 _2924_ (.A(_0486_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_o21ai_1 _2925_ (.B1(_0323_),
    .Y(_0489_),
    .A1(net564),
    .A2(_0459_));
 sg13g2_a21oi_1 _2926_ (.A1(net750),
    .A2(\sap_3_inst.alu.tmp[4] ),
    .Y(_0490_),
    .B1(_0449_));
 sg13g2_xor2_1 _2927_ (.B(_0490_),
    .A(_0479_),
    .X(_0491_));
 sg13g2_nand2b_1 _2928_ (.Y(_0492_),
    .B(_0452_),
    .A_N(_0491_));
 sg13g2_xnor2_1 _2929_ (.Y(_0493_),
    .A(_0452_),
    .B(_0491_));
 sg13g2_nor3_1 _2930_ (.A(net544),
    .B(_0481_),
    .C(_0484_),
    .Y(_0494_));
 sg13g2_a22oi_1 _2931_ (.Y(_0495_),
    .B1(_0493_),
    .B2(_0324_),
    .A2(_0489_),
    .A1(_0488_));
 sg13g2_nand3_1 _2932_ (.B(_0494_),
    .C(_0495_),
    .A(_0475_),
    .Y(_0496_));
 sg13g2_a21oi_1 _2933_ (.A1(net543),
    .A2(_0491_),
    .Y(_0497_),
    .B1(_0314_));
 sg13g2_a221oi_1 _2934_ (.B2(_0497_),
    .C1(_0310_),
    .B1(_0496_),
    .A1(\sap_3_inst.alu.act[5] ),
    .Y(_0498_),
    .A2(net669));
 sg13g2_a21oi_1 _2935_ (.A1(_1899_),
    .A2(net616),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_mux2_1 _2936_ (.A0(_0499_),
    .A1(net747),
    .S(net555),
    .X(_0039_));
 sg13g2_xnor2_1 _2937_ (.Y(_0500_),
    .A(net745),
    .B(net671));
 sg13g2_o21ai_1 _2938_ (.B1(_0471_),
    .Y(_0501_),
    .A1(net747),
    .A2(net671));
 sg13g2_a21oi_1 _2939_ (.A1(_0472_),
    .A2(_0501_),
    .Y(_0502_),
    .B1(_0500_));
 sg13g2_nand3_1 _2940_ (.B(_0500_),
    .C(_0501_),
    .A(_0472_),
    .Y(_0503_));
 sg13g2_nand3b_1 _2941_ (.B(_0503_),
    .C(_1936_),
    .Y(_0504_),
    .A_N(_0502_));
 sg13g2_nor2_2 _2942_ (.A(net745),
    .B(\sap_3_inst.alu.tmp[6] ),
    .Y(_0505_));
 sg13g2_nand2_2 _2943_ (.Y(_0506_),
    .A(net745),
    .B(\sap_3_inst.alu.tmp[6] ));
 sg13g2_nor2b_2 _2944_ (.A(_0505_),
    .B_N(_0506_),
    .Y(_0507_));
 sg13g2_a21oi_1 _2945_ (.A1(net748),
    .A2(_1466_),
    .Y(_0508_),
    .B1(_0487_));
 sg13g2_nor2_1 _2946_ (.A(_0507_),
    .B(_0508_),
    .Y(_0509_));
 sg13g2_xnor2_1 _2947_ (.Y(_0510_),
    .A(_0507_),
    .B(_0508_));
 sg13g2_nand2_1 _2948_ (.Y(_0511_),
    .A(_0482_),
    .B(_0510_));
 sg13g2_or2_1 _2949_ (.X(_0512_),
    .B(_0510_),
    .A(_0482_));
 sg13g2_a21oi_1 _2950_ (.A1(_0511_),
    .A2(_0512_),
    .Y(_0513_),
    .B1(_2007_));
 sg13g2_a21o_1 _2951_ (.A2(\sap_3_inst.alu.tmp[4] ),
    .A1(net750),
    .B1(_0477_),
    .X(_0514_));
 sg13g2_o21ai_1 _2952_ (.B1(_0478_),
    .Y(_0515_),
    .A1(_0449_),
    .A2(_0514_));
 sg13g2_xor2_1 _2953_ (.B(_0515_),
    .A(_0507_),
    .X(_0516_));
 sg13g2_and2_1 _2954_ (.A(_0492_),
    .B(_0516_),
    .X(_0517_));
 sg13g2_nor2_1 _2955_ (.A(_0492_),
    .B(_0516_),
    .Y(_0518_));
 sg13g2_nor3_1 _2956_ (.A(_0325_),
    .B(_0517_),
    .C(_0518_),
    .Y(_0519_));
 sg13g2_a21oi_1 _2957_ (.A1(_0333_),
    .A2(_0506_),
    .Y(_0520_),
    .B1(net563));
 sg13g2_nor3_1 _2958_ (.A(net618),
    .B(_0197_),
    .C(_0506_),
    .Y(_0521_));
 sg13g2_a221oi_1 _2959_ (.B2(net744),
    .C1(_0521_),
    .B1(net572),
    .A1(net748),
    .Y(_0522_),
    .A2(net573));
 sg13g2_or2_1 _2960_ (.X(_0523_),
    .B(_0510_),
    .A(_0323_));
 sg13g2_o21ai_1 _2961_ (.B1(_0522_),
    .Y(_0524_),
    .A1(_0505_),
    .A2(_0520_));
 sg13g2_o21ai_1 _2962_ (.B1(_0523_),
    .Y(_0525_),
    .A1(net745),
    .A2(_0327_));
 sg13g2_nor4_1 _2963_ (.A(_0513_),
    .B(_0519_),
    .C(_0524_),
    .D(_0525_),
    .Y(_0526_));
 sg13g2_nor2b_1 _2964_ (.A(net544),
    .B_N(_0526_),
    .Y(_0527_));
 sg13g2_nand2_1 _2965_ (.Y(_0528_),
    .A(net543),
    .B(_0516_));
 sg13g2_a21oi_1 _2966_ (.A1(_0504_),
    .A2(_0527_),
    .Y(_0529_),
    .B1(net670));
 sg13g2_nand2_1 _2967_ (.Y(_0530_),
    .A(_0528_),
    .B(_0529_));
 sg13g2_a21oi_1 _2968_ (.A1(\sap_3_inst.alu.act[6] ),
    .A2(net669),
    .Y(_0531_),
    .B1(net616));
 sg13g2_a221oi_1 _2969_ (.B2(_0531_),
    .C1(net554),
    .B1(_0530_),
    .A1(net547),
    .Y(_0532_),
    .A2(_0310_));
 sg13g2_a21o_1 _2970_ (.A2(net554),
    .A1(net745),
    .B1(_0532_),
    .X(_0040_));
 sg13g2_nor2b_1 _2971_ (.A(net542),
    .B_N(net617),
    .Y(_0533_));
 sg13g2_a21oi_1 _2972_ (.A1(net745),
    .A2(net672),
    .Y(_0534_),
    .B1(_0502_));
 sg13g2_xnor2_1 _2973_ (.Y(_0535_),
    .A(net743),
    .B(net671));
 sg13g2_o21ai_1 _2974_ (.B1(_1936_),
    .Y(_0536_),
    .A1(_0534_),
    .A2(_0535_));
 sg13g2_a21oi_1 _2975_ (.A1(_0534_),
    .A2(_0535_),
    .Y(_0537_),
    .B1(_0536_));
 sg13g2_or2_1 _2976_ (.X(_0538_),
    .B(\sap_3_inst.alu.tmp[7] ),
    .A(net743));
 sg13g2_and2_1 _2977_ (.A(net743),
    .B(\sap_3_inst.alu.tmp[7] ),
    .X(_0539_));
 sg13g2_xor2_1 _2978_ (.B(\sap_3_inst.alu.tmp[7] ),
    .A(net743),
    .X(_0540_));
 sg13g2_a21oi_1 _2979_ (.A1(net746),
    .A2(_1467_),
    .Y(_0541_),
    .B1(_0509_));
 sg13g2_xnor2_1 _2980_ (.Y(_0542_),
    .A(_0540_),
    .B(_0541_));
 sg13g2_nand2b_1 _2981_ (.Y(_0543_),
    .B(_0542_),
    .A_N(_0511_));
 sg13g2_xnor2_1 _2982_ (.Y(_0544_),
    .A(_0511_),
    .B(_0542_));
 sg13g2_a22oi_1 _2983_ (.Y(_0545_),
    .B1(_0340_),
    .B2(_0539_),
    .A2(net572),
    .A1(_0337_));
 sg13g2_a22oi_1 _2984_ (.Y(_0546_),
    .B1(_0540_),
    .B2(_0333_),
    .A2(net573),
    .A1(net746));
 sg13g2_nand2_1 _2985_ (.Y(_0547_),
    .A(_0330_),
    .B(_0538_));
 sg13g2_or2_1 _2986_ (.X(_0548_),
    .B(_0327_),
    .A(net744));
 sg13g2_and4_1 _2987_ (.A(_0545_),
    .B(_0546_),
    .C(_0547_),
    .D(_0548_),
    .X(_0549_));
 sg13g2_o21ai_1 _2988_ (.B1(_0549_),
    .Y(_0550_),
    .A1(_0323_),
    .A2(_0542_));
 sg13g2_o21ai_1 _2989_ (.B1(_0506_),
    .Y(_0551_),
    .A1(_0505_),
    .A2(_0515_));
 sg13g2_xnor2_1 _2990_ (.Y(_0552_),
    .A(_0540_),
    .B(_0551_));
 sg13g2_xnor2_1 _2991_ (.Y(_0553_),
    .A(_0518_),
    .B(_0552_));
 sg13g2_nand2_1 _2992_ (.Y(_0554_),
    .A(_0324_),
    .B(_0553_));
 sg13g2_o21ai_1 _2993_ (.B1(_0554_),
    .Y(_0555_),
    .A1(_2007_),
    .A2(_0544_));
 sg13g2_or4_1 _2994_ (.A(net544),
    .B(_0537_),
    .C(_0550_),
    .D(_0555_),
    .X(_0556_));
 sg13g2_a21oi_1 _2995_ (.A1(net543),
    .A2(_0552_),
    .Y(_0557_),
    .B1(net670));
 sg13g2_a221oi_1 _2996_ (.B2(_0557_),
    .C1(_0310_),
    .B1(_0556_),
    .A1(\sap_3_inst.alu.act[7] ),
    .Y(_0558_),
    .A2(net669));
 sg13g2_nor3_1 _2997_ (.A(net555),
    .B(_0533_),
    .C(_0558_),
    .Y(_0559_));
 sg13g2_a21o_1 _2998_ (.A2(net555),
    .A1(net743),
    .B1(_0559_),
    .X(_0041_));
 sg13g2_nand2_1 _2999_ (.Y(_0560_),
    .A(\sap_3_inst.out[0] ),
    .B(net673));
 sg13g2_o21ai_1 _3000_ (.B1(_0560_),
    .Y(_0042_),
    .A1(_1456_),
    .A2(net673));
 sg13g2_nand2_1 _3001_ (.Y(_0561_),
    .A(\sap_3_inst.out[1] ),
    .B(net673));
 sg13g2_o21ai_1 _3002_ (.B1(_0561_),
    .Y(_0043_),
    .A1(_1455_),
    .A2(net673));
 sg13g2_mux2_1 _3003_ (.A0(net756),
    .A1(\sap_3_inst.out[2] ),
    .S(net673),
    .X(_0044_));
 sg13g2_mux2_1 _3004_ (.A0(net754),
    .A1(\sap_3_inst.out[3] ),
    .S(net674),
    .X(_0045_));
 sg13g2_mux2_1 _3005_ (.A0(net752),
    .A1(\sap_3_inst.out[4] ),
    .S(net674),
    .X(_0046_));
 sg13g2_mux2_1 _3006_ (.A0(net749),
    .A1(\sap_3_inst.out[5] ),
    .S(net674),
    .X(_0047_));
 sg13g2_mux2_1 _3007_ (.A0(net746),
    .A1(\sap_3_inst.out[6] ),
    .S(net674),
    .X(_0048_));
 sg13g2_mux2_1 _3008_ (.A0(net744),
    .A1(\sap_3_inst.out[7] ),
    .S(net673),
    .X(_0049_));
 sg13g2_nand2b_1 _3009_ (.Y(_0562_),
    .B(_1938_),
    .A_N(_0204_));
 sg13g2_nor2b_1 _3010_ (.A(\sap_3_inst.alu.acc[7] ),
    .B_N(\sap_3_inst.alu.tmp[7] ),
    .Y(_0563_));
 sg13g2_nand2b_1 _3011_ (.Y(_0564_),
    .B(net744),
    .A_N(\sap_3_inst.alu.tmp[7] ));
 sg13g2_o21ai_1 _3012_ (.B1(_0564_),
    .Y(_0565_),
    .A1(_0541_),
    .A2(_0563_));
 sg13g2_a21oi_1 _3013_ (.A1(_0543_),
    .A2(_0565_),
    .Y(_0566_),
    .B1(net564));
 sg13g2_o21ai_1 _3014_ (.B1(_1944_),
    .Y(_0567_),
    .A1(net732),
    .A2(_1943_));
 sg13g2_nand4_1 _3015_ (.B(net564),
    .C(_0326_),
    .A(_1953_),
    .Y(_0568_),
    .D(_0567_));
 sg13g2_and3_1 _3016_ (.X(_0569_),
    .A(_0479_),
    .B(_0507_),
    .C(_0540_));
 sg13g2_nand2_1 _3017_ (.Y(_0570_),
    .A(_0447_),
    .B(_0569_));
 sg13g2_and4_1 _3018_ (.A(_0478_),
    .B(_0507_),
    .C(_0514_),
    .D(_0540_),
    .X(_0571_));
 sg13g2_a21o_1 _3019_ (.A2(\sap_3_inst.alu.tmp[6] ),
    .A1(net746),
    .B1(_0539_),
    .X(_0572_));
 sg13g2_a221oi_1 _3020_ (.B2(_0538_),
    .C1(_0571_),
    .B1(_0572_),
    .A1(_0449_),
    .Y(_0573_),
    .A2(_0569_));
 sg13g2_o21ai_1 _3021_ (.B1(_0573_),
    .Y(_0574_),
    .A1(_0426_),
    .A2(_0570_));
 sg13g2_nand2_1 _3022_ (.Y(_0575_),
    .A(_0324_),
    .B(_0574_));
 sg13g2_nand2_1 _3023_ (.Y(_0576_),
    .A(\sap_3_inst.alu.flags[1] ),
    .B(net618));
 sg13g2_nand3_1 _3024_ (.B(_0202_),
    .C(_0576_),
    .A(_1950_),
    .Y(_0577_));
 sg13g2_a22oi_1 _3025_ (.Y(_0578_),
    .B1(net572),
    .B2(net760),
    .A2(net573),
    .A1(net744));
 sg13g2_nand3_1 _3026_ (.B(_0577_),
    .C(_0578_),
    .A(_0575_),
    .Y(_0579_));
 sg13g2_o21ai_1 _3027_ (.B1(_0568_),
    .Y(_0580_),
    .A1(_0323_),
    .A2(_0565_));
 sg13g2_nor3_1 _3028_ (.A(_0566_),
    .B(_0579_),
    .C(_0580_),
    .Y(_0581_));
 sg13g2_nor2b_1 _3029_ (.A(_0568_),
    .B_N(_0573_),
    .Y(_0582_));
 sg13g2_nor3_1 _3030_ (.A(_0562_),
    .B(_0581_),
    .C(_0582_),
    .Y(_0583_));
 sg13g2_a21o_1 _3031_ (.A2(_0562_),
    .A1(\sap_3_inst.alu.carry ),
    .B1(_0583_),
    .X(_0050_));
 sg13g2_nand2_1 _3032_ (.Y(_0584_),
    .A(_1545_),
    .B(_1729_));
 sg13g2_o21ai_1 _3033_ (.B1(_1843_),
    .Y(_0585_),
    .A1(_1836_),
    .A2(_0584_));
 sg13g2_mux2_1 _3034_ (.A0(net17),
    .A1(\sap_3_inst.alu.tmp[0] ),
    .S(net668),
    .X(_0051_));
 sg13g2_nor2_1 _3035_ (.A(net18),
    .B(net668),
    .Y(_0586_));
 sg13g2_a21oi_1 _3036_ (.A1(_1463_),
    .A2(net668),
    .Y(_0052_),
    .B1(_0586_));
 sg13g2_mux2_1 _3037_ (.A0(net19),
    .A1(\sap_3_inst.alu.tmp[2] ),
    .S(net667),
    .X(_0053_));
 sg13g2_nand2_1 _3038_ (.Y(_0587_),
    .A(\sap_3_inst.alu.tmp[3] ),
    .B(net667));
 sg13g2_o21ai_1 _3039_ (.B1(_0587_),
    .Y(_0054_),
    .A1(net546),
    .A2(net667));
 sg13g2_nand2_1 _3040_ (.Y(_0588_),
    .A(\sap_3_inst.alu.tmp[4] ),
    .B(net667));
 sg13g2_o21ai_1 _3041_ (.B1(_0588_),
    .Y(_0055_),
    .A1(_1920_),
    .A2(net667));
 sg13g2_nand2_1 _3042_ (.Y(_0589_),
    .A(\sap_3_inst.alu.tmp[5] ),
    .B(net667));
 sg13g2_o21ai_1 _3043_ (.B1(_0589_),
    .Y(_0056_),
    .A1(_1899_),
    .A2(net667));
 sg13g2_nand2_1 _3044_ (.Y(_0590_),
    .A(\sap_3_inst.alu.tmp[6] ),
    .B(net668));
 sg13g2_o21ai_1 _3045_ (.B1(_0590_),
    .Y(_0057_),
    .A1(net547),
    .A2(net667));
 sg13g2_mux2_1 _3046_ (.A0(net24),
    .A1(\sap_3_inst.alu.tmp[7] ),
    .S(net668),
    .X(_0058_));
 sg13g2_mux2_1 _3047_ (.A0(net31),
    .A1(\sap_3_inst.controller.opcode[0] ),
    .S(net692),
    .X(_0059_));
 sg13g2_nand2_1 _3048_ (.Y(_0591_),
    .A(\sap_3_inst.controller.opcode[1] ),
    .B(net693));
 sg13g2_o21ai_1 _3049_ (.B1(_0591_),
    .Y(_0060_),
    .A1(net693),
    .A2(_0225_));
 sg13g2_nor2_1 _3050_ (.A(net692),
    .B(net19),
    .Y(_0592_));
 sg13g2_a21oi_1 _3051_ (.A1(_1436_),
    .A2(net692),
    .Y(_0061_),
    .B1(_0592_));
 sg13g2_nand2_1 _3052_ (.Y(_0593_),
    .A(net734),
    .B(net691));
 sg13g2_o21ai_1 _3053_ (.B1(_0593_),
    .Y(_0062_),
    .A1(net691),
    .A2(net546));
 sg13g2_nand2_1 _3054_ (.Y(_0594_),
    .A(net731),
    .B(net691));
 sg13g2_o21ai_1 _3055_ (.B1(_0594_),
    .Y(_0063_),
    .A1(net691),
    .A2(_1920_));
 sg13g2_nand2_1 _3056_ (.Y(_0595_),
    .A(net729),
    .B(net691));
 sg13g2_o21ai_1 _3057_ (.B1(_0595_),
    .Y(_0064_),
    .A1(net691),
    .A2(_1899_));
 sg13g2_nand2_1 _3058_ (.Y(_0596_),
    .A(net727),
    .B(net691));
 sg13g2_o21ai_1 _3059_ (.B1(_0596_),
    .Y(_0065_),
    .A1(net691),
    .A2(net547));
 sg13g2_nor2_1 _3060_ (.A(net692),
    .B(net24),
    .Y(_0597_));
 sg13g2_a21oi_1 _3061_ (.A1(_1439_),
    .A2(net692),
    .Y(_0066_),
    .B1(_0597_));
 sg13g2_nand3_1 _3062_ (.B(net696),
    .C(_1716_),
    .A(_1510_),
    .Y(_0598_));
 sg13g2_o21ai_1 _3063_ (.B1(net706),
    .Y(_0599_),
    .A1(_1577_),
    .A2(_1638_));
 sg13g2_nor2_1 _3064_ (.A(_1635_),
    .B(net684),
    .Y(_0600_));
 sg13g2_o21ai_1 _3065_ (.B1(_1594_),
    .Y(_0601_),
    .A1(_1581_),
    .A2(_1646_));
 sg13g2_a221oi_1 _3066_ (.B2(_1716_),
    .C1(net689),
    .B1(_1839_),
    .A1(net723),
    .Y(_0602_),
    .A2(_1838_));
 sg13g2_nor2_1 _3067_ (.A(_1582_),
    .B(_1662_),
    .Y(_0603_));
 sg13g2_o21ai_1 _3068_ (.B1(_1601_),
    .Y(_0604_),
    .A1(_1581_),
    .A2(_1626_));
 sg13g2_o21ai_1 _3069_ (.B1(_0604_),
    .Y(_0605_),
    .A1(_1607_),
    .A2(_0600_));
 sg13g2_nand4_1 _3070_ (.B(_0599_),
    .C(_0601_),
    .A(_1730_),
    .Y(_0606_),
    .D(_0602_));
 sg13g2_nor4_1 _3071_ (.A(_1835_),
    .B(_0603_),
    .C(_0605_),
    .D(_0606_),
    .Y(_0607_));
 sg13g2_o21ai_1 _3072_ (.B1(_0598_),
    .Y(_0608_),
    .A1(_0313_),
    .A2(_0607_));
 sg13g2_a21oi_1 _3073_ (.A1(_1515_),
    .A2(_0608_),
    .Y(_0609_),
    .B1(net713));
 sg13g2_nand3b_1 _3074_ (.B(_1830_),
    .C(_0298_),
    .Y(_0610_),
    .A_N(_0609_));
 sg13g2_o21ai_1 _3075_ (.B1(_0273_),
    .Y(_0611_),
    .A1(net700),
    .A2(_1704_));
 sg13g2_o21ai_1 _3076_ (.B1(_1615_),
    .Y(_0612_),
    .A1(net687),
    .A2(_1691_));
 sg13g2_nand2b_1 _3077_ (.Y(_0613_),
    .B(_1575_),
    .A_N(_1703_));
 sg13g2_and2_1 _3078_ (.A(net673),
    .B(_0613_),
    .X(_0614_));
 sg13g2_nand2_1 _3079_ (.Y(_0615_),
    .A(_1589_),
    .B(_1932_));
 sg13g2_o21ai_1 _3080_ (.B1(net687),
    .Y(_0616_),
    .A1(_1587_),
    .A2(_1592_));
 sg13g2_nor3_1 _3081_ (.A(net695),
    .B(_1588_),
    .C(_1622_),
    .Y(_0617_));
 sg13g2_nor4_1 _3082_ (.A(_1596_),
    .B(_1599_),
    .C(net707),
    .D(_1661_),
    .Y(_0618_));
 sg13g2_nand3_1 _3083_ (.B(_0614_),
    .C(_0615_),
    .A(_0612_),
    .Y(_0619_));
 sg13g2_a21oi_1 _3084_ (.A1(_0616_),
    .A2(_0618_),
    .Y(_0620_),
    .B1(_1703_));
 sg13g2_nor4_1 _3085_ (.A(_0263_),
    .B(_0617_),
    .C(_0619_),
    .D(_0620_),
    .Y(_0621_));
 sg13g2_a21oi_1 _3086_ (.A1(_0611_),
    .A2(_0621_),
    .Y(_0622_),
    .B1(_0275_));
 sg13g2_nand2_1 _3087_ (.Y(_0623_),
    .A(net698),
    .B(_1712_));
 sg13g2_o21ai_1 _3088_ (.B1(_1534_),
    .Y(_0624_),
    .A1(net733),
    .A2(_0623_));
 sg13g2_or2_1 _3089_ (.X(_0625_),
    .B(_0624_),
    .A(_0622_));
 sg13g2_nor2_1 _3090_ (.A(net707),
    .B(_0273_),
    .Y(_0626_));
 sg13g2_nand3_1 _3091_ (.B(net700),
    .C(_1712_),
    .A(net735),
    .Y(_0627_));
 sg13g2_nand2b_1 _3092_ (.Y(_0628_),
    .B(_1583_),
    .A_N(_1579_));
 sg13g2_o21ai_1 _3093_ (.B1(_0627_),
    .Y(_0629_),
    .A1(net708),
    .A2(_0628_));
 sg13g2_nor3_1 _3094_ (.A(net695),
    .B(_1606_),
    .C(_1622_),
    .Y(_0630_));
 sg13g2_nor3_1 _3095_ (.A(_0617_),
    .B(_0629_),
    .C(_0630_),
    .Y(_0631_));
 sg13g2_o21ai_1 _3096_ (.B1(_0631_),
    .Y(_0632_),
    .A1(_1651_),
    .A2(_0626_));
 sg13g2_inv_4 _3097_ (.A(net666),
    .Y(_0633_));
 sg13g2_nor2_1 _3098_ (.A(net660),
    .B(net666),
    .Y(_0634_));
 sg13g2_and2_1 _3099_ (.A(_0610_),
    .B(_0634_),
    .X(_0635_));
 sg13g2_nand4_1 _3100_ (.B(_1553_),
    .C(net684),
    .A(net731),
    .Y(_0636_),
    .D(_1716_));
 sg13g2_nand3_1 _3101_ (.B(_1549_),
    .C(net687),
    .A(net731),
    .Y(_0637_));
 sg13g2_nand3_1 _3102_ (.B(net714),
    .C(net704),
    .A(net731),
    .Y(_0638_));
 sg13g2_nand3_1 _3103_ (.B(_1581_),
    .C(_1620_),
    .A(_1575_),
    .Y(_0639_));
 sg13g2_and3_1 _3104_ (.X(_0640_),
    .A(_0613_),
    .B(_0628_),
    .C(_0639_));
 sg13g2_nand2b_1 _3105_ (.Y(_0641_),
    .B(net680),
    .A_N(_0640_));
 sg13g2_a21o_1 _3106_ (.A2(_1651_),
    .A1(net686),
    .B1(_1607_),
    .X(_0642_));
 sg13g2_a21o_1 _3107_ (.A2(_1658_),
    .A1(net686),
    .B1(_1616_),
    .X(_0643_));
 sg13g2_nand2_1 _3108_ (.Y(_0644_),
    .A(net686),
    .B(_1703_));
 sg13g2_o21ai_1 _3109_ (.B1(net686),
    .Y(_0645_),
    .A1(_1590_),
    .A2(_0638_));
 sg13g2_a22oi_1 _3110_ (.Y(_0646_),
    .B1(_0645_),
    .B2(_1594_),
    .A2(_0644_),
    .A1(_1601_));
 sg13g2_nor3_1 _3111_ (.A(_1715_),
    .B(_1818_),
    .C(_0603_),
    .Y(_0647_));
 sg13g2_and4_1 _3112_ (.A(_1730_),
    .B(_0636_),
    .C(_0637_),
    .D(_0643_),
    .X(_0648_));
 sg13g2_and4_1 _3113_ (.A(_0642_),
    .B(_0646_),
    .C(_0647_),
    .D(_0648_),
    .X(_0649_));
 sg13g2_a21oi_1 _3114_ (.A1(_0598_),
    .A2(_0623_),
    .Y(_0650_),
    .B1(_1437_));
 sg13g2_o21ai_1 _3115_ (.B1(_1515_),
    .Y(_0651_),
    .A1(net682),
    .A2(_0650_));
 sg13g2_a21o_2 _3116_ (.A2(_0649_),
    .A1(_0641_),
    .B1(_0651_),
    .X(_0652_));
 sg13g2_nand2_1 _3117_ (.Y(_0653_),
    .A(net702),
    .B(_0652_));
 sg13g2_a21oi_1 _3118_ (.A1(net731),
    .A2(_1716_),
    .Y(_0654_),
    .B1(net702));
 sg13g2_or3_1 _3119_ (.A(_1502_),
    .B(_1831_),
    .C(_0654_),
    .X(_0655_));
 sg13g2_inv_1 _3120_ (.Y(_0656_),
    .A(_0655_));
 sg13g2_a21oi_2 _3121_ (.B1(_0655_),
    .Y(_0657_),
    .A2(_0652_),
    .A1(net702));
 sg13g2_a21o_2 _3122_ (.A2(_0652_),
    .A1(net702),
    .B1(_0655_),
    .X(_0658_));
 sg13g2_nor2_1 _3123_ (.A(_1504_),
    .B(_1675_),
    .Y(_0659_));
 sg13g2_nand4_1 _3124_ (.B(_1439_),
    .C(_1508_),
    .A(net733),
    .Y(_0660_),
    .D(_0659_));
 sg13g2_o21ai_1 _3125_ (.B1(net733),
    .Y(_0661_),
    .A1(_1749_),
    .A2(_1814_));
 sg13g2_nand2_1 _3126_ (.Y(_0662_),
    .A(_1601_),
    .B(_1690_));
 sg13g2_nand4_1 _3127_ (.B(net724),
    .C(_1510_),
    .A(net734),
    .Y(_0663_),
    .D(net697));
 sg13g2_a22oi_1 _3128_ (.Y(_0664_),
    .B1(_0659_),
    .B2(_1575_),
    .A2(net706),
    .A1(_1577_));
 sg13g2_nand3_1 _3129_ (.B(_0663_),
    .C(_0664_),
    .A(_0662_),
    .Y(_0665_));
 sg13g2_nor3_1 _3130_ (.A(_1587_),
    .B(_1592_),
    .C(_1605_),
    .Y(_0666_));
 sg13g2_nor3_1 _3131_ (.A(_1594_),
    .B(_1608_),
    .C(_1609_),
    .Y(_0667_));
 sg13g2_o21ai_1 _3132_ (.B1(_0661_),
    .Y(_0668_),
    .A1(_1675_),
    .A2(_0667_));
 sg13g2_o21ai_1 _3133_ (.B1(net702),
    .Y(_0669_),
    .A1(_0665_),
    .A2(_0668_));
 sg13g2_and2_1 _3134_ (.A(_0660_),
    .B(_0669_),
    .X(_0670_));
 sg13g2_nand2_1 _3135_ (.Y(_0671_),
    .A(_0660_),
    .B(_0669_));
 sg13g2_nor2_2 _3136_ (.A(_0657_),
    .B(net665),
    .Y(_0672_));
 sg13g2_nand2_1 _3137_ (.Y(_0673_),
    .A(_0658_),
    .B(_0670_));
 sg13g2_nand3_1 _3138_ (.B(_0614_),
    .C(_0628_),
    .A(net680),
    .Y(_0674_));
 sg13g2_nand2_1 _3139_ (.Y(_0675_),
    .A(_1535_),
    .B(_1633_));
 sg13g2_nand2_1 _3140_ (.Y(_0676_),
    .A(_1627_),
    .B(_1703_));
 sg13g2_nor2_1 _3141_ (.A(_1604_),
    .B(_0675_),
    .Y(_0677_));
 sg13g2_nand4_1 _3142_ (.B(_1627_),
    .C(_1703_),
    .A(net694),
    .Y(_0678_),
    .D(_0675_));
 sg13g2_a21oi_1 _3143_ (.A1(_0273_),
    .A2(_0678_),
    .Y(_0679_),
    .B1(_0677_));
 sg13g2_a21oi_1 _3144_ (.A1(net695),
    .A2(_1703_),
    .Y(_0680_),
    .B1(_1588_));
 sg13g2_nand2_1 _3145_ (.Y(_0681_),
    .A(_1623_),
    .B(_0680_));
 sg13g2_o21ai_1 _3146_ (.B1(_0676_),
    .Y(_0682_),
    .A1(_1601_),
    .A2(net708));
 sg13g2_nand3_1 _3147_ (.B(_0681_),
    .C(_0682_),
    .A(_0679_),
    .Y(_0683_));
 sg13g2_a21oi_1 _3148_ (.A1(_1593_),
    .A2(_1662_),
    .Y(_0684_),
    .B1(_1703_));
 sg13g2_nor2_1 _3149_ (.A(_1786_),
    .B(_0684_),
    .Y(_0685_));
 sg13g2_nor2b_1 _3150_ (.A(net680),
    .B_N(_0685_),
    .Y(_0686_));
 sg13g2_nor3_2 _3151_ (.A(_1438_),
    .B(_1590_),
    .C(_0638_),
    .Y(_0687_));
 sg13g2_a221oi_1 _3152_ (.B2(_1589_),
    .C1(_0687_),
    .B1(_1932_),
    .A1(_1615_),
    .Y(_0688_),
    .A2(_1704_));
 sg13g2_nand3b_1 _3153_ (.B(_0685_),
    .C(_0688_),
    .Y(_0689_),
    .A_N(net680));
 sg13g2_o21ai_1 _3154_ (.B1(_0674_),
    .Y(_0690_),
    .A1(_0683_),
    .A2(_0689_));
 sg13g2_a21o_2 _3155_ (.A2(_0690_),
    .A1(_1569_),
    .B1(_0275_),
    .X(_0691_));
 sg13g2_nand2_1 _3156_ (.Y(_0692_),
    .A(_1534_),
    .B(_0623_));
 sg13g2_nand2_1 _3157_ (.Y(_0693_),
    .A(net724),
    .B(_1534_));
 sg13g2_nand2_2 _3158_ (.Y(_0694_),
    .A(_0692_),
    .B(_0693_));
 sg13g2_nand2_2 _3159_ (.Y(_0695_),
    .A(_0691_),
    .B(_0694_));
 sg13g2_a21oi_1 _3160_ (.A1(_0618_),
    .A2(_0666_),
    .Y(_0696_),
    .B1(net686));
 sg13g2_nand3_1 _3161_ (.B(_1614_),
    .C(net704),
    .A(net714),
    .Y(_0697_));
 sg13g2_a21o_1 _3162_ (.A2(_0697_),
    .A1(net686),
    .B1(_1590_),
    .X(_0698_));
 sg13g2_nand3_1 _3163_ (.B(_1581_),
    .C(_1614_),
    .A(_1575_),
    .Y(_0699_));
 sg13g2_nand3_1 _3164_ (.B(net684),
    .C(_1782_),
    .A(_1553_),
    .Y(_0700_));
 sg13g2_nand3_1 _3165_ (.B(_0699_),
    .C(_0700_),
    .A(_0698_),
    .Y(_0701_));
 sg13g2_o21ai_1 _3166_ (.B1(net734),
    .Y(_0702_),
    .A1(_1638_),
    .A2(_1641_));
 sg13g2_o21ai_1 _3167_ (.B1(_0643_),
    .Y(_0703_),
    .A1(_1616_),
    .A2(_0702_));
 sg13g2_nand3_1 _3168_ (.B(_1549_),
    .C(net687),
    .A(net729),
    .Y(_0704_));
 sg13g2_nand4_1 _3169_ (.B(_1730_),
    .C(_0599_),
    .A(net682),
    .Y(_0705_),
    .D(_0704_));
 sg13g2_nor4_1 _3170_ (.A(_0696_),
    .B(_0701_),
    .C(_0703_),
    .D(_0705_),
    .Y(_0706_));
 sg13g2_a21oi_1 _3171_ (.A1(net697),
    .A2(_1614_),
    .Y(_0707_),
    .B1(net682));
 sg13g2_nand2b_1 _3172_ (.Y(_0708_),
    .B(net713),
    .A_N(_1782_));
 sg13g2_o21ai_1 _3173_ (.B1(net702),
    .Y(_0709_),
    .A1(_0706_),
    .A2(_0707_));
 sg13g2_and3_2 _3174_ (.X(_0710_),
    .A(_1830_),
    .B(_0708_),
    .C(_0709_));
 sg13g2_nand3_1 _3175_ (.B(_0708_),
    .C(_0709_),
    .A(_1830_),
    .Y(_0711_));
 sg13g2_and3_2 _3176_ (.X(_0712_),
    .A(_0691_),
    .B(_0694_),
    .C(_0711_));
 sg13g2_nand3_1 _3177_ (.B(_0694_),
    .C(_0711_),
    .A(_0691_),
    .Y(_0713_));
 sg13g2_nor2_1 _3178_ (.A(_0673_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_nand2_2 _3179_ (.Y(_0715_),
    .A(_0672_),
    .B(net659));
 sg13g2_nand2b_2 _3180_ (.Y(_0716_),
    .B(net614),
    .A_N(_0635_));
 sg13g2_inv_4 _3181_ (.A(_0716_),
    .Y(_0717_));
 sg13g2_nand2_1 _3182_ (.Y(_0718_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][0] ),
    .B(_0716_));
 sg13g2_nor2_2 _3183_ (.A(_0658_),
    .B(net665),
    .Y(_0719_));
 sg13g2_nand2_1 _3184_ (.Y(_0720_),
    .A(_0657_),
    .B(_0670_));
 sg13g2_and2_1 _3185_ (.A(_0695_),
    .B(_0719_),
    .X(_0721_));
 sg13g2_nand2_2 _3186_ (.Y(_0722_),
    .A(_0695_),
    .B(_0719_));
 sg13g2_a221oi_1 _3187_ (.B2(_0694_),
    .C1(net665),
    .B1(_0691_),
    .A1(_0653_),
    .Y(_0723_),
    .A2(_0656_));
 sg13g2_nand2_2 _3188_ (.Y(_0724_),
    .A(_0672_),
    .B(_0695_));
 sg13g2_a22oi_1 _3189_ (.Y(_0725_),
    .B1(net657),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .A2(net609),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ));
 sg13g2_nor3_1 _3190_ (.A(_0657_),
    .B(net665),
    .C(_0711_),
    .Y(_0726_));
 sg13g2_nand2_2 _3191_ (.Y(_0727_),
    .A(_0672_),
    .B(_0710_));
 sg13g2_a221oi_1 _3192_ (.B2(_0669_),
    .C1(_0655_),
    .B1(_0660_),
    .A1(net702),
    .Y(_0728_),
    .A2(_0652_));
 sg13g2_and2_1 _3193_ (.A(_0710_),
    .B(_0728_),
    .X(_0729_));
 sg13g2_a22oi_1 _3194_ (.Y(_0730_),
    .B1(net649),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .A2(net653),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ));
 sg13g2_nand2_1 _3195_ (.Y(_0731_),
    .A(_0658_),
    .B(net665));
 sg13g2_nor3_1 _3196_ (.A(_0657_),
    .B(_0670_),
    .C(_0711_),
    .Y(_0732_));
 sg13g2_nor3_1 _3197_ (.A(_0658_),
    .B(net665),
    .C(_0711_),
    .Y(_0733_));
 sg13g2_nand2_2 _3198_ (.Y(_0734_),
    .A(_0710_),
    .B(_0719_));
 sg13g2_a22oi_1 _3199_ (.Y(_0735_),
    .B1(net644),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .A2(net646),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ));
 sg13g2_nand4_1 _3200_ (.B(_0725_),
    .C(_0730_),
    .A(net610),
    .Y(_0736_),
    .D(_0735_));
 sg13g2_and4_1 _3201_ (.A(_0691_),
    .B(_0694_),
    .C(_0711_),
    .D(_0728_),
    .X(_0737_));
 sg13g2_nor2_1 _3202_ (.A(_0713_),
    .B(_0720_),
    .Y(_0738_));
 sg13g2_nand2_1 _3203_ (.Y(_0739_),
    .A(net659),
    .B(_0719_));
 sg13g2_nor2_2 _3204_ (.A(_0713_),
    .B(_0731_),
    .Y(_0740_));
 sg13g2_a22oi_1 _3205_ (.Y(_0741_),
    .B1(net588),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ));
 sg13g2_o21ai_1 _3206_ (.B1(_0741_),
    .Y(_0742_),
    .A1(_1461_),
    .A2(net590));
 sg13g2_nand2_1 _3207_ (.Y(_0743_),
    .A(_1460_),
    .B(net615));
 sg13g2_o21ai_1 _3208_ (.B1(_0743_),
    .Y(_0744_),
    .A1(_0736_),
    .A2(_0742_));
 sg13g2_a22oi_1 _3209_ (.Y(_0745_),
    .B1(net646),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .A2(net649),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ));
 sg13g2_a22oi_1 _3210_ (.Y(_0746_),
    .B1(net643),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .A2(net652),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ));
 sg13g2_nand2_1 _3211_ (.Y(_0747_),
    .A(_0745_),
    .B(_0746_));
 sg13g2_a221oi_1 _3212_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ),
    .C1(_0747_),
    .B1(net658),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .Y(_0748_),
    .A2(net606));
 sg13g2_a22oi_1 _3213_ (.Y(_0749_),
    .B1(net587),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .A2(net592),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ));
 sg13g2_a22oi_1 _3214_ (.Y(_0750_),
    .B1(net640),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .A2(net612),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ));
 sg13g2_and3_2 _3215_ (.X(_0751_),
    .A(_0748_),
    .B(_0749_),
    .C(_0750_));
 sg13g2_a22oi_1 _3216_ (.Y(_0752_),
    .B1(net644),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .A2(net653),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ));
 sg13g2_a22oi_1 _3217_ (.Y(_0753_),
    .B1(net646),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .A2(_0729_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ));
 sg13g2_a22oi_1 _3218_ (.Y(_0754_),
    .B1(net593),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ));
 sg13g2_a22oi_1 _3219_ (.Y(_0755_),
    .B1(net588),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .A2(net657),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ));
 sg13g2_nand4_1 _3220_ (.B(_0753_),
    .C(_0754_),
    .A(_0752_),
    .Y(_0756_),
    .D(_0755_));
 sg13g2_a221oi_1 _3221_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .C1(_0756_),
    .B1(net609),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .Y(_0757_),
    .A2(net615));
 sg13g2_nand2_1 _3222_ (.Y(_0758_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .B(net606));
 sg13g2_nand2_1 _3223_ (.Y(_0759_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .B(net655));
 sg13g2_a22oi_1 _3224_ (.Y(_0760_),
    .B1(net649),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .A2(net651),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ));
 sg13g2_a22oi_1 _3225_ (.Y(_0761_),
    .B1(net643),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ),
    .A2(net646),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ));
 sg13g2_nand2_1 _3226_ (.Y(_0762_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .B(net640));
 sg13g2_nand3_1 _3227_ (.B(net659),
    .C(_0719_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .Y(_0763_));
 sg13g2_a22oi_1 _3228_ (.Y(_0764_),
    .B1(net587),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .A2(net613),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ));
 sg13g2_and4_1 _3229_ (.A(_0760_),
    .B(_0761_),
    .C(_0762_),
    .D(_0763_),
    .X(_0765_));
 sg13g2_and4_1 _3230_ (.A(_0758_),
    .B(_0759_),
    .C(_0764_),
    .D(_0765_),
    .X(_0766_));
 sg13g2_nand4_1 _3231_ (.B(_0759_),
    .C(_0764_),
    .A(_0758_),
    .Y(_0767_),
    .D(_0765_));
 sg13g2_a22oi_1 _3232_ (.Y(_0768_),
    .B1(net643),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .A2(net646),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ));
 sg13g2_a22oi_1 _3233_ (.Y(_0769_),
    .B1(net649),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .A2(net651),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ));
 sg13g2_nand2_1 _3234_ (.Y(_0770_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .B(net613));
 sg13g2_nand2_1 _3235_ (.Y(_0771_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ),
    .B(net640));
 sg13g2_a22oi_1 _3236_ (.Y(_0772_),
    .B1(net587),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .A2(net592),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ));
 sg13g2_a22oi_1 _3237_ (.Y(_0773_),
    .B1(net658),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .A2(net606),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ));
 sg13g2_and3_1 _3238_ (.X(_0774_),
    .A(_0768_),
    .B(_0769_),
    .C(_0771_));
 sg13g2_and4_1 _3239_ (.A(_0770_),
    .B(_0772_),
    .C(_0773_),
    .D(_0774_),
    .X(_0775_));
 sg13g2_nand4_1 _3240_ (.B(_0772_),
    .C(_0773_),
    .A(_0770_),
    .Y(_0776_),
    .D(_0774_));
 sg13g2_and2_1 _3241_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .B(net608),
    .X(_0777_));
 sg13g2_and2_1 _3242_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .B(net656),
    .X(_0778_));
 sg13g2_a22oi_1 _3243_ (.Y(_0779_),
    .B1(net648),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .A2(net650),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ));
 sg13g2_a22oi_1 _3244_ (.Y(_0780_),
    .B1(net645),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ),
    .A2(net653),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ));
 sg13g2_nand2_1 _3245_ (.Y(_0781_),
    .A(_0779_),
    .B(_0780_));
 sg13g2_nand2_1 _3246_ (.Y(_0782_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .B(net641));
 sg13g2_nand3_1 _3247_ (.B(net659),
    .C(_0719_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .Y(_0783_));
 sg13g2_nand3_1 _3248_ (.B(_0672_),
    .C(net659),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .Y(_0784_));
 sg13g2_nand4_1 _3249_ (.B(_0658_),
    .C(net665),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ),
    .Y(_0785_),
    .D(net659));
 sg13g2_nand4_1 _3250_ (.B(_0783_),
    .C(_0784_),
    .A(_0782_),
    .Y(_0786_),
    .D(_0785_));
 sg13g2_nor4_2 _3251_ (.A(_0777_),
    .B(_0778_),
    .C(_0781_),
    .Y(_0787_),
    .D(_0786_));
 sg13g2_or4_1 _3252_ (.A(_0777_),
    .B(_0778_),
    .C(_0781_),
    .D(_0786_),
    .X(_0788_));
 sg13g2_a22oi_1 _3253_ (.Y(_0789_),
    .B1(net644),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .A2(net654),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ));
 sg13g2_a22oi_1 _3254_ (.Y(_0790_),
    .B1(net647),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .A2(net650),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ));
 sg13g2_nand2_1 _3255_ (.Y(_0791_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .B(net642));
 sg13g2_nand2_1 _3256_ (.Y(_0792_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .B(net593));
 sg13g2_a22oi_1 _3257_ (.Y(_0793_),
    .B1(net588),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .A2(net615),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ));
 sg13g2_a22oi_1 _3258_ (.Y(_0794_),
    .B1(net657),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .A2(net609),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ));
 sg13g2_and3_1 _3259_ (.X(_0795_),
    .A(_0789_),
    .B(_0790_),
    .C(_0791_));
 sg13g2_and4_1 _3260_ (.A(_0792_),
    .B(_0793_),
    .C(_0794_),
    .D(_0795_),
    .X(_0796_));
 sg13g2_inv_2 _3261_ (.Y(_0797_),
    .A(net560));
 sg13g2_nand2_1 _3262_ (.Y(_0798_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ),
    .B(net656));
 sg13g2_a22oi_1 _3263_ (.Y(_0799_),
    .B1(net645),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ),
    .A2(net648),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ));
 sg13g2_a22oi_1 _3264_ (.Y(_0800_),
    .B1(net650),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .A2(net653),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ));
 sg13g2_nand3_1 _3265_ (.B(_0695_),
    .C(_0719_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .Y(_0801_));
 sg13g2_and4_1 _3266_ (.A(_0798_),
    .B(_0799_),
    .C(_0800_),
    .D(_0801_),
    .X(_0802_));
 sg13g2_nor3_1 _3267_ (.A(_1454_),
    .B(_0673_),
    .C(_0713_),
    .Y(_0803_));
 sg13g2_and2_1 _3268_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .B(net640),
    .X(_0804_));
 sg13g2_nor3_1 _3269_ (.A(_1453_),
    .B(_0713_),
    .C(_0731_),
    .Y(_0805_));
 sg13g2_nor3_1 _3270_ (.A(_1452_),
    .B(_0713_),
    .C(_0720_),
    .Y(_0806_));
 sg13g2_nor4_1 _3271_ (.A(_0803_),
    .B(_0804_),
    .C(_0805_),
    .D(_0806_),
    .Y(_0807_));
 sg13g2_and2_1 _3272_ (.A(_0802_),
    .B(_0807_),
    .X(_0808_));
 sg13g2_nand4_1 _3273_ (.B(_0658_),
    .C(_0670_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .Y(_0809_),
    .D(_0710_));
 sg13g2_nand3_1 _3274_ (.B(_0710_),
    .C(_0728_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .Y(_0810_));
 sg13g2_nand4_1 _3275_ (.B(_0658_),
    .C(net665),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .Y(_0811_),
    .D(_0710_));
 sg13g2_nand4_1 _3276_ (.B(_0657_),
    .C(_0670_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .Y(_0812_),
    .D(_0710_));
 sg13g2_nand4_1 _3277_ (.B(_0810_),
    .C(_0811_),
    .A(_0809_),
    .Y(_0813_),
    .D(_0812_));
 sg13g2_a221oi_1 _3278_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .C1(_0813_),
    .B1(net656),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .Y(_0814_),
    .A2(net608));
 sg13g2_nand4_1 _3279_ (.B(_0658_),
    .C(_0671_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .Y(_0815_),
    .D(net659));
 sg13g2_nand2_1 _3280_ (.Y(_0816_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .B(net641));
 sg13g2_nand3_1 _3281_ (.B(net659),
    .C(_0719_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .Y(_0817_));
 sg13g2_nand3_1 _3282_ (.B(_0672_),
    .C(_0712_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .Y(_0818_));
 sg13g2_and4_1 _3283_ (.A(_0815_),
    .B(_0816_),
    .C(_0817_),
    .D(_0818_),
    .X(_0819_));
 sg13g2_and2_1 _3284_ (.A(_0814_),
    .B(_0819_),
    .X(_0820_));
 sg13g2_nand2_1 _3285_ (.Y(_0821_),
    .A(net561),
    .B(_0820_));
 sg13g2_nand3_1 _3286_ (.B(_0808_),
    .C(_0820_),
    .A(net561),
    .Y(_0822_));
 sg13g2_and4_1 _3287_ (.A(_0787_),
    .B(net560),
    .C(_0808_),
    .D(_0820_),
    .X(_0823_));
 sg13g2_nand3_1 _3288_ (.B(_0775_),
    .C(_0823_),
    .A(_0766_),
    .Y(_0824_));
 sg13g2_and4_1 _3289_ (.A(_0757_),
    .B(_0766_),
    .C(_0775_),
    .D(_0823_),
    .X(_0825_));
 sg13g2_nand2_1 _3290_ (.Y(_0826_),
    .A(net553),
    .B(_0825_));
 sg13g2_nand3_1 _3291_ (.B(net553),
    .C(_0825_),
    .A(_0744_),
    .Y(_0827_));
 sg13g2_xnor2_1 _3292_ (.Y(_0828_),
    .A(_0744_),
    .B(_0826_));
 sg13g2_nor2_1 _3293_ (.A(net660),
    .B(_0633_),
    .Y(_0829_));
 sg13g2_nand2b_2 _3294_ (.Y(_0830_),
    .B(net666),
    .A_N(net660));
 sg13g2_mux2_1 _3295_ (.A0(_0797_),
    .A1(_0828_),
    .S(net614),
    .X(_0831_));
 sg13g2_a21oi_1 _3296_ (.A1(_1589_),
    .A2(_0676_),
    .Y(_0832_),
    .B1(_1657_));
 sg13g2_nand3_1 _3297_ (.B(_0686_),
    .C(_0832_),
    .A(_0612_),
    .Y(_0833_));
 sg13g2_o21ai_1 _3298_ (.B1(_0674_),
    .Y(_0834_),
    .A1(_0683_),
    .A2(_0833_));
 sg13g2_a21oi_1 _3299_ (.A1(_1569_),
    .A2(_0834_),
    .Y(_0835_),
    .B1(_0275_));
 sg13g2_nor2_2 _3300_ (.A(_0692_),
    .B(_0835_),
    .Y(_0836_));
 sg13g2_nand2b_1 _3301_ (.Y(_0837_),
    .B(net614),
    .A_N(_0836_));
 sg13g2_inv_4 _3302_ (.A(net571),
    .Y(_0838_));
 sg13g2_nand2_1 _3303_ (.Y(_0839_),
    .A(net31),
    .B(net571));
 sg13g2_a21oi_1 _3304_ (.A1(net9),
    .A2(_0838_),
    .Y(_0840_),
    .B1(net584));
 sg13g2_a22oi_1 _3305_ (.Y(_0841_),
    .B1(_0839_),
    .B2(_0840_),
    .A2(_0831_),
    .A1(net586));
 sg13g2_and2_1 _3306_ (.A(net660),
    .B(_0633_),
    .X(_0842_));
 sg13g2_nand2_2 _3307_ (.Y(_0843_),
    .A(net660),
    .B(_0633_));
 sg13g2_and2_1 _3308_ (.A(net660),
    .B(net666),
    .X(_0844_));
 sg13g2_nand2_1 _3309_ (.Y(_0845_),
    .A(net661),
    .B(net666));
 sg13g2_o21ai_1 _3310_ (.B1(net575),
    .Y(_0846_),
    .A1(net561),
    .A2(net574));
 sg13g2_inv_1 _3311_ (.Y(_0847_),
    .A(_0846_));
 sg13g2_nor2_1 _3312_ (.A(_0841_),
    .B(_0846_),
    .Y(_0848_));
 sg13g2_a22oi_1 _3313_ (.Y(_0849_),
    .B1(_0814_),
    .B2(_0819_),
    .A2(_0807_),
    .A1(_0802_));
 sg13g2_or2_1 _3314_ (.X(_0850_),
    .B(_0820_),
    .A(_0808_));
 sg13g2_nand2_1 _3315_ (.Y(_0851_),
    .A(_0788_),
    .B(_0849_));
 sg13g2_nor2_1 _3316_ (.A(_0775_),
    .B(_0851_),
    .Y(_0852_));
 sg13g2_nand3_1 _3317_ (.B(_0788_),
    .C(_0849_),
    .A(_0776_),
    .Y(_0853_));
 sg13g2_nand4_1 _3318_ (.B(_0776_),
    .C(_0788_),
    .A(_0767_),
    .Y(_0854_),
    .D(_0849_));
 sg13g2_or2_1 _3319_ (.X(_0855_),
    .B(_0854_),
    .A(_0757_));
 sg13g2_or2_1 _3320_ (.X(_0856_),
    .B(_0855_),
    .A(net553));
 sg13g2_nor4_2 _3321_ (.A(_0744_),
    .B(net553),
    .C(_0757_),
    .Y(_0857_),
    .D(_0854_));
 sg13g2_nor2_1 _3322_ (.A(net559),
    .B(_0856_),
    .Y(_0858_));
 sg13g2_nand2_1 _3323_ (.Y(_0859_),
    .A(_0797_),
    .B(_0857_));
 sg13g2_xnor2_1 _3324_ (.Y(_0860_),
    .A(_0744_),
    .B(_0858_));
 sg13g2_nor2_1 _3325_ (.A(net575),
    .B(_0860_),
    .Y(_0861_));
 sg13g2_o21ai_1 _3326_ (.B1(_0717_),
    .Y(_0862_),
    .A1(_0843_),
    .A2(_0860_));
 sg13g2_o21ai_1 _3327_ (.B1(_0718_),
    .Y(_0067_),
    .A1(_0848_),
    .A2(_0862_));
 sg13g2_nor2_1 _3328_ (.A(_1457_),
    .B(_0717_),
    .Y(_0863_));
 sg13g2_a22oi_1 _3329_ (.Y(_0864_),
    .B1(net656),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .A2(net608),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ));
 sg13g2_a22oi_1 _3330_ (.Y(_0865_),
    .B1(net645),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .A2(net648),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ));
 sg13g2_a22oi_1 _3331_ (.Y(_0866_),
    .B1(net650),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .A2(net653),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ));
 sg13g2_and3_1 _3332_ (.X(_0867_),
    .A(net611),
    .B(_0865_),
    .C(_0866_));
 sg13g2_nand2_1 _3333_ (.Y(_0868_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .B(net641));
 sg13g2_a22oi_1 _3334_ (.Y(_0869_),
    .B1(net588),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .A2(net592),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ));
 sg13g2_nand4_1 _3335_ (.B(_0867_),
    .C(_0868_),
    .A(_0864_),
    .Y(_0870_),
    .D(_0869_));
 sg13g2_o21ai_1 _3336_ (.B1(_0870_),
    .Y(_0871_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[0][1] ),
    .A2(net610));
 sg13g2_inv_2 _3337_ (.Y(_0872_),
    .A(_0871_));
 sg13g2_nand2_2 _3338_ (.Y(_0873_),
    .A(_0857_),
    .B(_0872_));
 sg13g2_xnor2_1 _3339_ (.Y(_0874_),
    .A(_0859_),
    .B(_0871_));
 sg13g2_or2_1 _3340_ (.X(_0875_),
    .B(_0820_),
    .A(net561));
 sg13g2_and2_1 _3341_ (.A(_0821_),
    .B(_0875_),
    .X(_0876_));
 sg13g2_a21oi_1 _3342_ (.A1(net582),
    .A2(_0874_),
    .Y(_0877_),
    .B1(net562));
 sg13g2_nand2b_1 _3343_ (.Y(_0878_),
    .B(_0838_),
    .A_N(net10));
 sg13g2_o21ai_1 _3344_ (.B1(_0878_),
    .Y(_0879_),
    .A1(net32),
    .A2(_0838_));
 sg13g2_nand2_1 _3345_ (.Y(_0880_),
    .A(_0820_),
    .B(_0844_));
 sg13g2_and2_1 _3346_ (.A(_0744_),
    .B(_0871_),
    .X(_0881_));
 sg13g2_and3_2 _3347_ (.X(_0882_),
    .A(net553),
    .B(_0825_),
    .C(_0881_));
 sg13g2_xnor2_1 _3348_ (.Y(_0883_),
    .A(_0827_),
    .B(_0872_));
 sg13g2_nand2_2 _3349_ (.Y(_0884_),
    .A(net584),
    .B(_0883_));
 sg13g2_inv_1 _3350_ (.Y(_0885_),
    .A(_0884_));
 sg13g2_nand4_1 _3351_ (.B(_0879_),
    .C(_0880_),
    .A(net576),
    .Y(_0886_),
    .D(_0884_));
 sg13g2_a21o_1 _3352_ (.A2(_0886_),
    .A1(_0877_),
    .B1(_0863_),
    .X(_0068_));
 sg13g2_a22oi_1 _3353_ (.Y(_0887_),
    .B1(net648),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .A2(net650),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ));
 sg13g2_a22oi_1 _3354_ (.Y(_0888_),
    .B1(net645),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .A2(net653),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ));
 sg13g2_and3_1 _3355_ (.X(_0889_),
    .A(net611),
    .B(_0887_),
    .C(_0888_));
 sg13g2_a22oi_1 _3356_ (.Y(_0890_),
    .B1(net656),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .A2(net608),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ));
 sg13g2_nand2_1 _3357_ (.Y(_0891_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .B(net592));
 sg13g2_a22oi_1 _3358_ (.Y(_0892_),
    .B1(net588),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ));
 sg13g2_nand4_1 _3359_ (.B(_0890_),
    .C(_0891_),
    .A(_0889_),
    .Y(_0893_),
    .D(_0892_));
 sg13g2_o21ai_1 _3360_ (.B1(_0893_),
    .Y(_0894_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[0][2] ),
    .A2(net610));
 sg13g2_inv_1 _3361_ (.Y(_0895_),
    .A(_0894_));
 sg13g2_o21ai_1 _3362_ (.B1(_0894_),
    .Y(_0896_),
    .A1(net560),
    .A2(_0873_));
 sg13g2_nand4_1 _3363_ (.B(_0857_),
    .C(_0872_),
    .A(_0797_),
    .Y(_0897_),
    .D(_0895_));
 sg13g2_and2_1 _3364_ (.A(_0896_),
    .B(_0897_),
    .X(_0898_));
 sg13g2_nand2_1 _3365_ (.Y(_0899_),
    .A(net577),
    .B(_0898_));
 sg13g2_xnor2_1 _3366_ (.Y(_0900_),
    .A(_0882_),
    .B(_0894_));
 sg13g2_a22oi_1 _3367_ (.Y(_0901_),
    .B1(_0900_),
    .B2(net584),
    .A2(_0898_),
    .A1(net577));
 sg13g2_nor2_1 _3368_ (.A(net19),
    .B(_0838_),
    .Y(_0902_));
 sg13g2_nor2_1 _3369_ (.A(net11),
    .B(net571),
    .Y(_0903_));
 sg13g2_nor3_1 _3370_ (.A(_0610_),
    .B(_0902_),
    .C(_0903_),
    .Y(_0904_));
 sg13g2_a22oi_1 _3371_ (.Y(_0905_),
    .B1(_0904_),
    .B2(net614),
    .A2(net562),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[0][2] ));
 sg13g2_xnor2_1 _3372_ (.Y(_0906_),
    .A(_0808_),
    .B(_0875_));
 sg13g2_nand2b_1 _3373_ (.Y(_0907_),
    .B(_0821_),
    .A_N(_0808_));
 sg13g2_o21ai_1 _3374_ (.B1(_0905_),
    .Y(_0069_),
    .A1(net562),
    .A2(_0901_));
 sg13g2_nand2_1 _3375_ (.Y(_0908_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][3] ),
    .B(_0716_));
 sg13g2_a22oi_1 _3376_ (.Y(_0909_),
    .B1(net588),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .A2(net641),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ));
 sg13g2_o21ai_1 _3377_ (.B1(_0909_),
    .Y(_0910_),
    .A1(_1443_),
    .A2(net590));
 sg13g2_a22oi_1 _3378_ (.Y(_0911_),
    .B1(net656),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .A2(net608),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ));
 sg13g2_a22oi_1 _3379_ (.Y(_0912_),
    .B1(net648),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .A2(net653),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ));
 sg13g2_a22oi_1 _3380_ (.Y(_0913_),
    .B1(net645),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .A2(net650),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ));
 sg13g2_nand4_1 _3381_ (.B(_0911_),
    .C(_0912_),
    .A(net611),
    .Y(_0914_),
    .D(_0913_));
 sg13g2_nand2_1 _3382_ (.Y(_0915_),
    .A(_1440_),
    .B(net615));
 sg13g2_o21ai_1 _3383_ (.B1(_0915_),
    .Y(_0916_),
    .A1(_0910_),
    .A2(_0914_));
 sg13g2_inv_1 _3384_ (.Y(_0917_),
    .A(_0916_));
 sg13g2_nand4_1 _3385_ (.B(_0872_),
    .C(_0895_),
    .A(_0857_),
    .Y(_0918_),
    .D(_0917_));
 sg13g2_nor2_1 _3386_ (.A(net560),
    .B(_0918_),
    .Y(_0919_));
 sg13g2_a21o_1 _3387_ (.A2(_0916_),
    .A1(_0897_),
    .B1(_0919_),
    .X(_0920_));
 sg13g2_nand2_2 _3388_ (.Y(_0921_),
    .A(net577),
    .B(_0920_));
 sg13g2_nand2b_1 _3389_ (.Y(_0922_),
    .B(_0797_),
    .A_N(_0851_));
 sg13g2_o21ai_1 _3390_ (.B1(_0787_),
    .Y(_0923_),
    .A1(net560),
    .A2(_0850_));
 sg13g2_and2_1 _3391_ (.A(_0922_),
    .B(_0923_),
    .X(_0924_));
 sg13g2_nand2_1 _3392_ (.Y(_0925_),
    .A(_0717_),
    .B(_0921_));
 sg13g2_nor2_1 _3393_ (.A(net12),
    .B(net571),
    .Y(_0926_));
 sg13g2_a21oi_1 _3394_ (.A1(net546),
    .A2(_0837_),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_a21oi_1 _3395_ (.A1(_0787_),
    .A2(_0850_),
    .Y(_0928_),
    .B1(net574));
 sg13g2_a21o_2 _3396_ (.A2(_0928_),
    .A1(_0851_),
    .B1(net580),
    .X(_0929_));
 sg13g2_and2_1 _3397_ (.A(_0894_),
    .B(_0916_),
    .X(_0930_));
 sg13g2_nand4_1 _3398_ (.B(_0825_),
    .C(_0881_),
    .A(net553),
    .Y(_0931_),
    .D(_0930_));
 sg13g2_a21o_1 _3399_ (.A2(_0894_),
    .A1(_0882_),
    .B1(_0916_),
    .X(_0932_));
 sg13g2_a21oi_2 _3400_ (.B1(net583),
    .Y(_0933_),
    .A2(_0932_),
    .A1(_0931_));
 sg13g2_nor3_1 _3401_ (.A(_0927_),
    .B(_0929_),
    .C(_0933_),
    .Y(_0934_));
 sg13g2_xnor2_1 _3402_ (.Y(_0935_),
    .A(_0787_),
    .B(_0822_));
 sg13g2_o21ai_1 _3403_ (.B1(_0908_),
    .Y(_0070_),
    .A1(_0925_),
    .A2(_0934_));
 sg13g2_nand2_1 _3404_ (.Y(_0936_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[0][4] ),
    .B(net562));
 sg13g2_a22oi_1 _3405_ (.Y(_0937_),
    .B1(net655),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .A2(net606),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ));
 sg13g2_a22oi_1 _3406_ (.Y(_0938_),
    .B1(net643),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .A2(net646),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ));
 sg13g2_a22oi_1 _3407_ (.Y(_0939_),
    .B1(net649),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .A2(net651),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ));
 sg13g2_nand4_1 _3408_ (.B(_0937_),
    .C(_0938_),
    .A(net610),
    .Y(_0940_),
    .D(_0939_));
 sg13g2_a22oi_1 _3409_ (.Y(_0941_),
    .B1(net587),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .A2(net640),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ));
 sg13g2_o21ai_1 _3410_ (.B1(_0941_),
    .Y(_0942_),
    .A1(_1474_),
    .A2(net589));
 sg13g2_nand2_1 _3411_ (.Y(_0943_),
    .A(_1468_),
    .B(net612));
 sg13g2_o21ai_1 _3412_ (.B1(_0943_),
    .Y(_0944_),
    .A1(_0940_),
    .A2(_0942_));
 sg13g2_inv_1 _3413_ (.Y(_0945_),
    .A(net552));
 sg13g2_xnor2_1 _3414_ (.Y(_0946_),
    .A(_0931_),
    .B(_0945_));
 sg13g2_xnor2_1 _3415_ (.Y(_0947_),
    .A(_0775_),
    .B(_0823_));
 sg13g2_mux2_1 _3416_ (.A0(_0946_),
    .A1(_0947_),
    .S(net610),
    .X(_0948_));
 sg13g2_nand2_1 _3417_ (.Y(_0949_),
    .A(_1920_),
    .B(net571));
 sg13g2_nand2b_1 _3418_ (.Y(_0950_),
    .B(_0838_),
    .A_N(net13));
 sg13g2_a21oi_1 _3419_ (.A1(_0788_),
    .A2(_0849_),
    .Y(_0951_),
    .B1(_0776_));
 sg13g2_nor3_1 _3420_ (.A(net574),
    .B(_0852_),
    .C(_0951_),
    .Y(_0952_));
 sg13g2_or2_1 _3421_ (.X(_0953_),
    .B(_0952_),
    .A(net579));
 sg13g2_a221oi_1 _3422_ (.B2(_0950_),
    .C1(_0953_),
    .B1(_0949_),
    .A1(net584),
    .Y(_0954_),
    .A2(_0948_));
 sg13g2_nor2_1 _3423_ (.A(_0918_),
    .B(net552),
    .Y(_0955_));
 sg13g2_nor3_1 _3424_ (.A(net559),
    .B(_0918_),
    .C(net552),
    .Y(_0956_));
 sg13g2_xnor2_1 _3425_ (.Y(_0957_),
    .A(_0919_),
    .B(net552));
 sg13g2_a22oi_1 _3426_ (.Y(_0958_),
    .B1(_0922_),
    .B2(_0775_),
    .A2(_0852_),
    .A1(_0797_));
 sg13g2_inv_1 _3427_ (.Y(_0959_),
    .A(_0958_));
 sg13g2_o21ai_1 _3428_ (.B1(_0717_),
    .Y(_0960_),
    .A1(net576),
    .A2(_0957_));
 sg13g2_o21ai_1 _3429_ (.B1(_0936_),
    .Y(_0071_),
    .A1(_0954_),
    .A2(_0960_));
 sg13g2_a22oi_1 _3430_ (.Y(_0961_),
    .B1(net655),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .A2(net606),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ));
 sg13g2_a22oi_1 _3431_ (.Y(_0962_),
    .B1(net643),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .A2(net651),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ));
 sg13g2_a22oi_1 _3432_ (.Y(_0963_),
    .B1(net646),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .A2(net649),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ));
 sg13g2_nand4_1 _3433_ (.B(_0961_),
    .C(_0962_),
    .A(net610),
    .Y(_0964_),
    .D(_0963_));
 sg13g2_nand2_1 _3434_ (.Y(_0965_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .B(net587));
 sg13g2_a22oi_1 _3435_ (.Y(_0966_),
    .B1(net592),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .A2(net640),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ));
 sg13g2_nand3b_1 _3436_ (.B(_0965_),
    .C(_0966_),
    .Y(_0967_),
    .A_N(_0964_));
 sg13g2_nand2_1 _3437_ (.Y(_0968_),
    .A(_1475_),
    .B(net612));
 sg13g2_and2_1 _3438_ (.A(_0967_),
    .B(_0968_),
    .X(_0969_));
 sg13g2_nand2_2 _3439_ (.Y(_0970_),
    .A(_0967_),
    .B(_0968_));
 sg13g2_nand4_1 _3440_ (.B(_0930_),
    .C(net552),
    .A(_0882_),
    .Y(_0971_),
    .D(_0970_));
 sg13g2_o21ai_1 _3441_ (.B1(_0969_),
    .Y(_0972_),
    .A1(_0931_),
    .A2(_0945_));
 sg13g2_nand2_1 _3442_ (.Y(_0973_),
    .A(_0971_),
    .B(_0972_));
 sg13g2_a21o_1 _3443_ (.A2(_0823_),
    .A1(_0775_),
    .B1(_0766_),
    .X(_0974_));
 sg13g2_and2_1 _3444_ (.A(_0824_),
    .B(_0974_),
    .X(_0975_));
 sg13g2_o21ai_1 _3445_ (.B1(net585),
    .Y(_0976_),
    .A1(net612),
    .A2(_0975_));
 sg13g2_a21oi_1 _3446_ (.A1(net612),
    .A2(_0973_),
    .Y(_0977_),
    .B1(_0976_));
 sg13g2_a21oi_1 _3447_ (.A1(net14),
    .A2(_0838_),
    .Y(_0978_),
    .B1(_0632_));
 sg13g2_o21ai_1 _3448_ (.B1(_0978_),
    .Y(_0979_),
    .A1(_1899_),
    .A2(_0838_));
 sg13g2_nor2b_1 _3449_ (.A(net661),
    .B_N(_0979_),
    .Y(_0980_));
 sg13g2_nand2b_1 _3450_ (.Y(_0981_),
    .B(_0980_),
    .A_N(_0977_));
 sg13g2_or4_1 _3451_ (.A(net559),
    .B(_0918_),
    .C(net552),
    .D(_0970_),
    .X(_0982_));
 sg13g2_xnor2_1 _3452_ (.Y(_0983_),
    .A(_0956_),
    .B(_0970_));
 sg13g2_nand2_1 _3453_ (.Y(_0984_),
    .A(net578),
    .B(_0983_));
 sg13g2_a21oi_1 _3454_ (.A1(net578),
    .A2(_0983_),
    .Y(_0985_),
    .B1(net562));
 sg13g2_o21ai_1 _3455_ (.B1(_0766_),
    .Y(_0986_),
    .A1(net559),
    .A2(_0853_));
 sg13g2_o21ai_1 _3456_ (.B1(_0986_),
    .Y(_0987_),
    .A1(net559),
    .A2(_0854_));
 sg13g2_a22oi_1 _3457_ (.Y(_0072_),
    .B1(_0981_),
    .B2(_0985_),
    .A2(net562),
    .A1(_1475_));
 sg13g2_and2_1 _3458_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .B(net641),
    .X(_0988_));
 sg13g2_a221oi_1 _3459_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .C1(_0988_),
    .B1(net588),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .Y(_0989_),
    .A2(net593));
 sg13g2_a22oi_1 _3460_ (.Y(_0990_),
    .B1(net649),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .A2(net654),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ));
 sg13g2_a22oi_1 _3461_ (.Y(_0991_),
    .B1(net644),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .A2(net647),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ));
 sg13g2_nand3_1 _3462_ (.B(_0990_),
    .C(_0991_),
    .A(net611),
    .Y(_0992_));
 sg13g2_a221oi_1 _3463_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .C1(_0992_),
    .B1(net657),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ),
    .Y(_0993_),
    .A2(net609));
 sg13g2_a22oi_1 _3464_ (.Y(_0994_),
    .B1(_0989_),
    .B2(_0993_),
    .A2(net615),
    .A1(_1479_));
 sg13g2_inv_1 _3465_ (.Y(_0995_),
    .A(_0994_));
 sg13g2_nand2_1 _3466_ (.Y(_0996_),
    .A(_0969_),
    .B(_0994_));
 sg13g2_nor3_1 _3467_ (.A(_0918_),
    .B(net552),
    .C(_0996_),
    .Y(_0997_));
 sg13g2_nor4_1 _3468_ (.A(net559),
    .B(_0918_),
    .C(_0944_),
    .D(_0996_),
    .Y(_0998_));
 sg13g2_a21oi_2 _3469_ (.B1(_0998_),
    .Y(_0999_),
    .A2(_0995_),
    .A1(_0982_));
 sg13g2_o21ai_1 _3470_ (.B1(_0757_),
    .Y(_1000_),
    .A1(net559),
    .A2(_0854_));
 sg13g2_o21ai_1 _3471_ (.B1(_1000_),
    .Y(_1001_),
    .A1(net560),
    .A2(_0855_));
 sg13g2_nor2_2 _3472_ (.A(net575),
    .B(_1001_),
    .Y(_1002_));
 sg13g2_a21oi_1 _3473_ (.A1(net611),
    .A2(_1001_),
    .Y(_1003_),
    .B1(net575));
 sg13g2_o21ai_1 _3474_ (.B1(_1003_),
    .Y(_1004_),
    .A1(net611),
    .A2(_0999_));
 sg13g2_nor4_1 _3475_ (.A(_0931_),
    .B(_0945_),
    .C(_0969_),
    .D(_0994_),
    .Y(_1005_));
 sg13g2_xnor2_1 _3476_ (.Y(_1006_),
    .A(_0971_),
    .B(_0994_));
 sg13g2_xor2_1 _3477_ (.B(_0824_),
    .A(_0757_),
    .X(_1007_));
 sg13g2_o21ai_1 _3478_ (.B1(net586),
    .Y(_1008_),
    .A1(net615),
    .A2(_1007_));
 sg13g2_inv_1 _3479_ (.Y(_1009_),
    .A(_1008_));
 sg13g2_o21ai_1 _3480_ (.B1(_1009_),
    .Y(_1010_),
    .A1(net611),
    .A2(_1006_));
 sg13g2_nand2_1 _3481_ (.Y(_1011_),
    .A(net547),
    .B(net571));
 sg13g2_o21ai_1 _3482_ (.B1(_1011_),
    .Y(_1012_),
    .A1(net15),
    .A2(net571));
 sg13g2_nand3_1 _3483_ (.B(_1010_),
    .C(_1012_),
    .A(_1004_),
    .Y(_1013_));
 sg13g2_mux2_1 _3484_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[0][6] ),
    .A1(_1013_),
    .S(_0717_),
    .X(_0073_));
 sg13g2_a22oi_1 _3485_ (.Y(_1014_),
    .B1(net646),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .A2(net649),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ));
 sg13g2_a22oi_1 _3486_ (.Y(_1015_),
    .B1(net643),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .A2(net651),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ));
 sg13g2_a22oi_1 _3487_ (.Y(_1016_),
    .B1(net658),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .A2(net606),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ));
 sg13g2_nand4_1 _3488_ (.B(_1014_),
    .C(_1015_),
    .A(net610),
    .Y(_1017_),
    .D(_1016_));
 sg13g2_nand2_1 _3489_ (.Y(_1018_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .B(net640));
 sg13g2_a221oi_1 _3490_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .C1(_1017_),
    .B1(net587),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .Y(_1019_),
    .A2(net592));
 sg13g2_a22oi_1 _3491_ (.Y(_1020_),
    .B1(_1018_),
    .B2(_1019_),
    .A2(net612),
    .A1(_1490_));
 sg13g2_xnor2_1 _3492_ (.Y(_1021_),
    .A(_0998_),
    .B(_1020_));
 sg13g2_nand2b_1 _3493_ (.Y(_1022_),
    .B(net612),
    .A_N(_1021_));
 sg13g2_o21ai_1 _3494_ (.B1(net553),
    .Y(_1023_),
    .A1(net559),
    .A2(_0855_));
 sg13g2_nor2b_2 _3495_ (.A(_0858_),
    .B_N(_1023_),
    .Y(_1024_));
 sg13g2_nor2_1 _3496_ (.A(net576),
    .B(_1024_),
    .Y(_1025_));
 sg13g2_a21oi_1 _3497_ (.A1(net610),
    .A2(_1024_),
    .Y(_1026_),
    .B1(net576));
 sg13g2_xnor2_1 _3498_ (.Y(_1027_),
    .A(_1005_),
    .B(_1020_));
 sg13g2_xnor2_1 _3499_ (.Y(_1028_),
    .A(net553),
    .B(_0825_));
 sg13g2_o21ai_1 _3500_ (.B1(net585),
    .Y(_1029_),
    .A1(net612),
    .A2(_1028_));
 sg13g2_a21o_1 _3501_ (.A2(_1027_),
    .A1(net613),
    .B1(_1029_),
    .X(_1030_));
 sg13g2_mux2_1 _3502_ (.A0(net24),
    .A1(net16),
    .S(_0838_),
    .X(_1031_));
 sg13g2_xnor2_1 _3503_ (.Y(_1032_),
    .A(_0751_),
    .B(_0855_));
 sg13g2_nor2_1 _3504_ (.A(net574),
    .B(_1032_),
    .Y(_1033_));
 sg13g2_nor3_1 _3505_ (.A(net578),
    .B(_1031_),
    .C(_1033_),
    .Y(_1034_));
 sg13g2_a221oi_1 _3506_ (.B2(_1034_),
    .C1(net562),
    .B1(_1030_),
    .A1(_1022_),
    .Y(_1035_),
    .A2(_1026_));
 sg13g2_a21o_1 _3507_ (.A2(net562),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[0][7] ),
    .B1(_1035_),
    .X(_0074_));
 sg13g2_a21oi_1 _3508_ (.A1(_0610_),
    .A2(net614),
    .Y(_1036_),
    .B1(net587));
 sg13g2_a21o_1 _3509_ (.A2(_1036_),
    .A1(net571),
    .B1(_0635_),
    .X(_1037_));
 sg13g2_nand2_1 _3510_ (.Y(_1038_),
    .A(net561),
    .B(net586));
 sg13g2_inv_1 _3511_ (.Y(_1039_),
    .A(_1038_));
 sg13g2_nor3_2 _3512_ (.A(net31),
    .B(_0846_),
    .C(_1039_),
    .Y(_1040_));
 sg13g2_nor2_2 _3513_ (.A(net561),
    .B(net575),
    .Y(_1041_));
 sg13g2_nor3_1 _3514_ (.A(net557),
    .B(_1040_),
    .C(_1041_),
    .Y(_1042_));
 sg13g2_a21o_1 _3515_ (.A2(net557),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .B1(_1042_),
    .X(_0075_));
 sg13g2_nor2_1 _3516_ (.A(net583),
    .B(_0876_),
    .Y(_1043_));
 sg13g2_o21ai_1 _3517_ (.B1(net586),
    .Y(_1044_),
    .A1(net655),
    .A2(_0876_));
 sg13g2_nor2b_1 _3518_ (.A(net660),
    .B_N(_1044_),
    .Y(_1045_));
 sg13g2_or2_1 _3519_ (.X(_1046_),
    .B(_1043_),
    .A(net32));
 sg13g2_a21o_2 _3520_ (.A2(_0876_),
    .A1(net580),
    .B1(_1046_),
    .X(_1047_));
 sg13g2_mux2_1 _3521_ (.A0(_1047_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .S(net557),
    .X(_0076_));
 sg13g2_a21oi_1 _3522_ (.A1(_0822_),
    .A2(_0907_),
    .Y(_1048_),
    .B1(net583));
 sg13g2_nor2_2 _3523_ (.A(net19),
    .B(_1048_),
    .Y(_1049_));
 sg13g2_nor2_2 _3524_ (.A(net575),
    .B(_0906_),
    .Y(_1050_));
 sg13g2_nor2_1 _3525_ (.A(net557),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_a22oi_1 _3526_ (.Y(_0077_),
    .B1(_1049_),
    .B2(_1051_),
    .A2(net557),
    .A1(_1454_));
 sg13g2_nor2_1 _3527_ (.A(net583),
    .B(_0935_),
    .Y(_1052_));
 sg13g2_nor2_1 _3528_ (.A(_0929_),
    .B(_1052_),
    .Y(_1053_));
 sg13g2_nand2_1 _3529_ (.Y(_1054_),
    .A(_1975_),
    .B(_1053_));
 sg13g2_nand2b_2 _3530_ (.Y(_1055_),
    .B(net580),
    .A_N(_0924_));
 sg13g2_nor2b_1 _3531_ (.A(net557),
    .B_N(_1055_),
    .Y(_1056_));
 sg13g2_a22oi_1 _3532_ (.Y(_1057_),
    .B1(_1054_),
    .B2(_1056_),
    .A2(net557),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ));
 sg13g2_inv_1 _3533_ (.Y(_0078_),
    .A(_1057_));
 sg13g2_nand2_1 _3534_ (.Y(_1058_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .B(net558));
 sg13g2_a21o_2 _3535_ (.A2(_0947_),
    .A1(net584),
    .B1(net21),
    .X(_1059_));
 sg13g2_nor2_1 _3536_ (.A(_0953_),
    .B(_1059_),
    .Y(_1060_));
 sg13g2_o21ai_1 _3537_ (.B1(net579),
    .Y(_1061_),
    .A1(net587),
    .A2(_0959_));
 sg13g2_nand2b_1 _3538_ (.Y(_1062_),
    .B(_1061_),
    .A_N(net558));
 sg13g2_o21ai_1 _3539_ (.B1(_1058_),
    .Y(_0079_),
    .A1(_1060_),
    .A2(_1062_));
 sg13g2_nor2_2 _3540_ (.A(net583),
    .B(_0975_),
    .Y(_1063_));
 sg13g2_nor2_1 _3541_ (.A(net22),
    .B(_1063_),
    .Y(_1064_));
 sg13g2_nor2_1 _3542_ (.A(net576),
    .B(_0987_),
    .Y(_1065_));
 sg13g2_nor2_1 _3543_ (.A(net558),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_a22oi_1 _3544_ (.Y(_0080_),
    .B1(_1064_),
    .B2(_1066_),
    .A2(net558),
    .A1(_1478_));
 sg13g2_nand2_1 _3545_ (.Y(_1067_),
    .A(net586),
    .B(_1007_));
 sg13g2_nand2_2 _3546_ (.Y(_1068_),
    .A(net547),
    .B(_1067_));
 sg13g2_nand2_1 _3547_ (.Y(_1069_),
    .A(_0844_),
    .B(_0855_));
 sg13g2_a21oi_1 _3548_ (.A1(_0757_),
    .A2(_0854_),
    .Y(_1070_),
    .B1(_1069_));
 sg13g2_or2_1 _3549_ (.X(_1071_),
    .B(_1070_),
    .A(_1068_));
 sg13g2_nor3_1 _3550_ (.A(_1002_),
    .B(net557),
    .C(_1068_),
    .Y(_1072_));
 sg13g2_a21oi_1 _3551_ (.A1(_1489_),
    .A2(net558),
    .Y(_0081_),
    .B1(_1072_));
 sg13g2_nand2_1 _3552_ (.Y(_1073_),
    .A(net585),
    .B(_1028_));
 sg13g2_inv_1 _3553_ (.Y(_1074_),
    .A(_1073_));
 sg13g2_nor4_1 _3554_ (.A(net24),
    .B(net578),
    .C(_1033_),
    .D(_1074_),
    .Y(_1075_));
 sg13g2_nor3_1 _3555_ (.A(_1025_),
    .B(net558),
    .C(_1075_),
    .Y(_1076_));
 sg13g2_a21o_1 _3556_ (.A2(net558),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .B1(_1076_),
    .X(_0082_));
 sg13g2_nand2b_2 _3557_ (.Y(_1077_),
    .B(net592),
    .A_N(_0836_));
 sg13g2_inv_4 _3558_ (.A(net570),
    .Y(_1078_));
 sg13g2_nand2_1 _3559_ (.Y(_1079_),
    .A(net31),
    .B(_1077_));
 sg13g2_a21oi_1 _3560_ (.A1(net9),
    .A2(_1078_),
    .Y(_1080_),
    .B1(_0829_));
 sg13g2_a21oi_1 _3561_ (.A1(net590),
    .A2(net561),
    .Y(_1081_),
    .B1(_0830_));
 sg13g2_a22oi_1 _3562_ (.Y(_1082_),
    .B1(_1081_),
    .B2(_0828_),
    .A2(_1080_),
    .A1(_1079_));
 sg13g2_nor2_1 _3563_ (.A(_0846_),
    .B(_1082_),
    .Y(_1083_));
 sg13g2_nor3_1 _3564_ (.A(net590),
    .B(_0861_),
    .C(_1083_),
    .Y(_1084_));
 sg13g2_a21o_1 _3565_ (.A2(net590),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .B1(_1084_),
    .X(_0083_));
 sg13g2_mux2_1 _3566_ (.A0(net32),
    .A1(net10),
    .S(_1078_),
    .X(_1085_));
 sg13g2_nand2_2 _3567_ (.Y(_1086_),
    .A(net576),
    .B(_0880_));
 sg13g2_nor2_1 _3568_ (.A(_1085_),
    .B(_1086_),
    .Y(_1087_));
 sg13g2_a221oi_1 _3569_ (.B2(_1087_),
    .C1(net589),
    .B1(_0884_),
    .A1(net577),
    .Y(_1088_),
    .A2(_0874_));
 sg13g2_a21o_1 _3570_ (.A2(net589),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .B1(_1088_),
    .X(_0084_));
 sg13g2_a21o_1 _3571_ (.A2(net570),
    .A1(net19),
    .B1(net666),
    .X(_1089_));
 sg13g2_a21oi_1 _3572_ (.A1(net11),
    .A2(_1078_),
    .Y(_1090_),
    .B1(_1089_));
 sg13g2_nor2_1 _3573_ (.A(_0633_),
    .B(_0900_),
    .Y(_1091_));
 sg13g2_or3_1 _3574_ (.A(net660),
    .B(_1090_),
    .C(_1091_),
    .X(_1092_));
 sg13g2_a21oi_1 _3575_ (.A1(net577),
    .A2(_0898_),
    .Y(_1093_),
    .B1(net589));
 sg13g2_a22oi_1 _3576_ (.Y(_0085_),
    .B1(_1092_),
    .B2(_1093_),
    .A2(net589),
    .A1(_1453_));
 sg13g2_nand2_1 _3577_ (.Y(_1094_),
    .A(net590),
    .B(_0935_));
 sg13g2_nand2_1 _3578_ (.Y(_1095_),
    .A(net546),
    .B(net570));
 sg13g2_nand2b_1 _3579_ (.Y(_1096_),
    .B(_1078_),
    .A_N(net12));
 sg13g2_a221oi_1 _3580_ (.B2(_1096_),
    .C1(_0929_),
    .B1(_1095_),
    .A1(_0933_),
    .Y(_1097_),
    .A2(_1094_));
 sg13g2_nand3b_1 _3581_ (.B(net593),
    .C(_0921_),
    .Y(_1098_),
    .A_N(_1097_));
 sg13g2_o21ai_1 _3582_ (.B1(_1098_),
    .Y(_0086_),
    .A1(_1443_),
    .A2(net593));
 sg13g2_nor2_1 _3583_ (.A(net13),
    .B(net570),
    .Y(_1099_));
 sg13g2_a21oi_1 _3584_ (.A1(_1920_),
    .A2(net570),
    .Y(_1100_),
    .B1(_1099_));
 sg13g2_nor2_1 _3585_ (.A(net589),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_nand2_1 _3586_ (.Y(_1102_),
    .A(net577),
    .B(_0957_));
 sg13g2_a22oi_1 _3587_ (.Y(_1103_),
    .B1(_0957_),
    .B2(net577),
    .A2(_0946_),
    .A1(net584));
 sg13g2_a22oi_1 _3588_ (.Y(_0087_),
    .B1(_1101_),
    .B2(_1103_),
    .A2(net589),
    .A1(_1474_));
 sg13g2_nand2_1 _3589_ (.Y(_1104_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .B(net591));
 sg13g2_a221oi_1 _3590_ (.B2(net589),
    .C1(net583),
    .B1(_0975_),
    .A1(_0971_),
    .Y(_1105_),
    .A2(_0972_));
 sg13g2_nor2_1 _3591_ (.A(net14),
    .B(net570),
    .Y(_1106_));
 sg13g2_a21oi_1 _3592_ (.A1(_1899_),
    .A2(net570),
    .Y(_1107_),
    .B1(_1106_));
 sg13g2_nand2_1 _3593_ (.Y(_1108_),
    .A(_0844_),
    .B(_0854_));
 sg13g2_a21oi_1 _3594_ (.A1(_0766_),
    .A2(_0853_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_or2_1 _3595_ (.X(_1110_),
    .B(_1109_),
    .A(net578));
 sg13g2_nor3_1 _3596_ (.A(_1105_),
    .B(_1107_),
    .C(_1110_),
    .Y(_1111_));
 sg13g2_nand2b_2 _3597_ (.Y(_1112_),
    .B(net579),
    .A_N(_0983_));
 sg13g2_nand2_1 _3598_ (.Y(_1113_),
    .A(net592),
    .B(_1112_));
 sg13g2_o21ai_1 _3599_ (.B1(_1104_),
    .Y(_0088_),
    .A1(_1111_),
    .A2(_1113_));
 sg13g2_nand2_1 _3600_ (.Y(_1114_),
    .A(net581),
    .B(_0999_));
 sg13g2_a21oi_1 _3601_ (.A1(net581),
    .A2(_0999_),
    .Y(_1115_),
    .B1(net590));
 sg13g2_nand2b_1 _3602_ (.Y(_1116_),
    .B(net591),
    .A_N(_1007_));
 sg13g2_and2_1 _3603_ (.A(net586),
    .B(_1006_),
    .X(_1117_));
 sg13g2_nand2_1 _3604_ (.Y(_1118_),
    .A(net547),
    .B(_1077_));
 sg13g2_nand2b_1 _3605_ (.Y(_1119_),
    .B(_1078_),
    .A_N(net15));
 sg13g2_a221oi_1 _3606_ (.B2(_1119_),
    .C1(_1070_),
    .B1(_1118_),
    .A1(_1116_),
    .Y(_1120_),
    .A2(_1117_));
 sg13g2_a22oi_1 _3607_ (.Y(_0089_),
    .B1(_1115_),
    .B2(_1120_),
    .A2(net590),
    .A1(_1488_));
 sg13g2_nand2_1 _3608_ (.Y(_1121_),
    .A(net24),
    .B(net570));
 sg13g2_a21oi_1 _3609_ (.A1(net16),
    .A2(_1078_),
    .Y(_1122_),
    .B1(_0632_));
 sg13g2_a221oi_1 _3610_ (.B2(_1122_),
    .C1(net661),
    .B1(_1121_),
    .A1(net666),
    .Y(_1123_),
    .A2(_1027_));
 sg13g2_nor2_1 _3611_ (.A(net591),
    .B(_1123_),
    .Y(_1124_));
 sg13g2_nand2b_2 _3612_ (.Y(_1125_),
    .B(net579),
    .A_N(_1021_));
 sg13g2_a22oi_1 _3613_ (.Y(_0090_),
    .B1(_1124_),
    .B2(_1125_),
    .A2(net591),
    .A1(_1496_));
 sg13g2_nor2_2 _3614_ (.A(net640),
    .B(_1078_),
    .Y(_1126_));
 sg13g2_nor3_1 _3615_ (.A(_1040_),
    .B(_1041_),
    .C(net550),
    .Y(_1127_));
 sg13g2_a21o_1 _3616_ (.A2(net551),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .B1(_1127_),
    .X(_0091_));
 sg13g2_mux2_1 _3617_ (.A0(_1047_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .S(net550),
    .X(_0092_));
 sg13g2_nor2_1 _3618_ (.A(_1050_),
    .B(net551),
    .Y(_1128_));
 sg13g2_a22oi_1 _3619_ (.Y(_0093_),
    .B1(_1128_),
    .B2(_1049_),
    .A2(net551),
    .A1(_1452_));
 sg13g2_nand2_1 _3620_ (.Y(_1129_),
    .A(net580),
    .B(_0924_));
 sg13g2_nand3b_1 _3621_ (.B(_1129_),
    .C(net546),
    .Y(_1130_),
    .A_N(_1052_));
 sg13g2_mux2_1 _3622_ (.A0(_1130_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .S(net551),
    .X(_0094_));
 sg13g2_nand2_1 _3623_ (.Y(_1131_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .B(net550));
 sg13g2_o21ai_1 _3624_ (.B1(_1061_),
    .Y(_1132_),
    .A1(net642),
    .A2(_1078_));
 sg13g2_o21ai_1 _3625_ (.B1(_1131_),
    .Y(_0095_),
    .A1(_1060_),
    .A2(_1132_));
 sg13g2_nor3_2 _3626_ (.A(net22),
    .B(_1063_),
    .C(_1110_),
    .Y(_1133_));
 sg13g2_and2_1 _3627_ (.A(net579),
    .B(_0987_),
    .X(_1134_));
 sg13g2_nor3_1 _3628_ (.A(net550),
    .B(_1133_),
    .C(_1134_),
    .Y(_1135_));
 sg13g2_a21o_1 _3629_ (.A2(net550),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .B1(_1135_),
    .X(_0096_));
 sg13g2_nor3_1 _3630_ (.A(_1002_),
    .B(_1068_),
    .C(net550),
    .Y(_1136_));
 sg13g2_a21oi_1 _3631_ (.A1(_1487_),
    .A2(net551),
    .Y(_0097_),
    .B1(_1136_));
 sg13g2_nor3_1 _3632_ (.A(_1025_),
    .B(_1075_),
    .C(net550),
    .Y(_1137_));
 sg13g2_a21o_1 _3633_ (.A2(net550),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .B1(_1137_),
    .X(_0098_));
 sg13g2_o21ai_1 _3634_ (.B1(_0847_),
    .Y(_1138_),
    .A1(_0828_),
    .A2(_0830_));
 sg13g2_nand2b_1 _3635_ (.Y(_1139_),
    .B(net652),
    .A_N(_0836_));
 sg13g2_nand2b_1 _3636_ (.Y(_1140_),
    .B(net568),
    .A_N(net31));
 sg13g2_or2_1 _3637_ (.X(_1141_),
    .B(net569),
    .A(net9));
 sg13g2_a221oi_1 _3638_ (.B2(_1141_),
    .C1(_1138_),
    .B1(_1140_),
    .A1(_0727_),
    .Y(_1142_),
    .A2(_1039_));
 sg13g2_nor3_1 _3639_ (.A(net597),
    .B(_0861_),
    .C(_1142_),
    .Y(_1143_));
 sg13g2_a21o_1 _3640_ (.A2(net597),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .B1(_1143_),
    .X(_0099_));
 sg13g2_nor2_1 _3641_ (.A(net576),
    .B(_0874_),
    .Y(_1144_));
 sg13g2_mux2_1 _3642_ (.A0(net10),
    .A1(net32),
    .S(net568),
    .X(_1145_));
 sg13g2_nor4_1 _3643_ (.A(net596),
    .B(_0885_),
    .C(_1144_),
    .D(_1145_),
    .Y(_1146_));
 sg13g2_a21oi_1 _3644_ (.A1(_1459_),
    .A2(net596),
    .Y(_0100_),
    .B1(_1146_));
 sg13g2_mux2_1 _3645_ (.A0(net11),
    .A1(net19),
    .S(_0836_),
    .X(_1147_));
 sg13g2_nor2_1 _3646_ (.A(net596),
    .B(_1147_),
    .Y(_1148_));
 sg13g2_a22oi_1 _3647_ (.Y(_0101_),
    .B1(_0901_),
    .B2(_1148_),
    .A2(net596),
    .A1(_1451_));
 sg13g2_nand2_1 _3648_ (.Y(_1149_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .B(net597));
 sg13g2_nand2_1 _3649_ (.Y(_1150_),
    .A(net546),
    .B(net568));
 sg13g2_or2_1 _3650_ (.X(_1151_),
    .B(net569),
    .A(net12));
 sg13g2_nand2_1 _3651_ (.Y(_1152_),
    .A(_0727_),
    .B(_0935_));
 sg13g2_a221oi_1 _3652_ (.B2(_0933_),
    .C1(_0929_),
    .B1(_1152_),
    .A1(_1150_),
    .Y(_1153_),
    .A2(_1151_));
 sg13g2_nand2_1 _3653_ (.Y(_1154_),
    .A(net653),
    .B(_0921_));
 sg13g2_o21ai_1 _3654_ (.B1(_1149_),
    .Y(_0102_),
    .A1(_1153_),
    .A2(_1154_));
 sg13g2_o21ai_1 _3655_ (.B1(_0946_),
    .Y(_1155_),
    .A1(net652),
    .A2(_0947_));
 sg13g2_nor2_1 _3656_ (.A(net13),
    .B(net568),
    .Y(_1156_));
 sg13g2_a21oi_1 _3657_ (.A1(_1920_),
    .A2(net568),
    .Y(_1157_),
    .B1(_1156_));
 sg13g2_nor2_1 _3658_ (.A(net584),
    .B(_1157_),
    .Y(_1158_));
 sg13g2_a21oi_1 _3659_ (.A1(net584),
    .A2(_1155_),
    .Y(_1159_),
    .B1(_1158_));
 sg13g2_nor2_1 _3660_ (.A(net596),
    .B(_1159_),
    .Y(_1160_));
 sg13g2_a22oi_1 _3661_ (.Y(_0103_),
    .B1(_1102_),
    .B2(_1160_),
    .A2(net596),
    .A1(_1473_));
 sg13g2_nand2_1 _3662_ (.Y(_1161_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .B(net596));
 sg13g2_a221oi_1 _3663_ (.B2(net596),
    .C1(net583),
    .B1(_0975_),
    .A1(_0971_),
    .Y(_1162_),
    .A2(_0972_));
 sg13g2_nor2_1 _3664_ (.A(net14),
    .B(net568),
    .Y(_1163_));
 sg13g2_a21oi_1 _3665_ (.A1(_1899_),
    .A2(net568),
    .Y(_1164_),
    .B1(_1163_));
 sg13g2_nor3_1 _3666_ (.A(_1110_),
    .B(_1162_),
    .C(_1164_),
    .Y(_1165_));
 sg13g2_nand2_1 _3667_ (.Y(_1166_),
    .A(net651),
    .B(_1112_));
 sg13g2_o21ai_1 _3668_ (.B1(_1161_),
    .Y(_0104_),
    .A1(_1165_),
    .A2(_1166_));
 sg13g2_a21oi_1 _3669_ (.A1(net581),
    .A2(_0999_),
    .Y(_1167_),
    .B1(net597));
 sg13g2_nand2b_1 _3670_ (.Y(_1168_),
    .B(net597),
    .A_N(_1007_));
 sg13g2_nand2_1 _3671_ (.Y(_1169_),
    .A(net547),
    .B(net569));
 sg13g2_or2_1 _3672_ (.X(_1170_),
    .B(net569),
    .A(net15));
 sg13g2_a221oi_1 _3673_ (.B2(_1170_),
    .C1(_1070_),
    .B1(_1169_),
    .A1(_1117_),
    .Y(_1171_),
    .A2(_1168_));
 sg13g2_a22oi_1 _3674_ (.Y(_0105_),
    .B1(_1167_),
    .B2(_1171_),
    .A2(net597),
    .A1(_1486_));
 sg13g2_nor2_1 _3675_ (.A(net606),
    .B(_1032_),
    .Y(_1172_));
 sg13g2_nor2_1 _3676_ (.A(net574),
    .B(_1172_),
    .Y(_1173_));
 sg13g2_nor2_1 _3677_ (.A(net578),
    .B(_1173_),
    .Y(_1174_));
 sg13g2_mux2_1 _3678_ (.A0(net16),
    .A1(net24),
    .S(net568),
    .X(_1175_));
 sg13g2_or2_1 _3679_ (.X(_1176_),
    .B(_1175_),
    .A(net661));
 sg13g2_o21ai_1 _3680_ (.B1(net585),
    .Y(_1177_),
    .A1(net651),
    .A2(_1028_));
 sg13g2_nor2_1 _3681_ (.A(_1027_),
    .B(_1177_),
    .Y(_1178_));
 sg13g2_o21ai_1 _3682_ (.B1(_1174_),
    .Y(_1179_),
    .A1(_1176_),
    .A2(_1178_));
 sg13g2_and2_1 _3683_ (.A(net651),
    .B(_1125_),
    .X(_1180_));
 sg13g2_a22oi_1 _3684_ (.Y(_0106_),
    .B1(_1179_),
    .B2(_1180_),
    .A2(net597),
    .A1(_1495_));
 sg13g2_nor2b_2 _3685_ (.A(net647),
    .B_N(net569),
    .Y(_1181_));
 sg13g2_nand2b_2 _3686_ (.Y(_1182_),
    .B(net569),
    .A_N(net647));
 sg13g2_nor3_1 _3687_ (.A(_1040_),
    .B(_1041_),
    .C(_1181_),
    .Y(_1183_));
 sg13g2_a21o_1 _3688_ (.A2(_1181_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .B1(_1183_),
    .X(_0107_));
 sg13g2_nor2_2 _3689_ (.A(_1046_),
    .B(_1086_),
    .Y(_1184_));
 sg13g2_nor2_2 _3690_ (.A(net575),
    .B(_0876_),
    .Y(_1185_));
 sg13g2_nor3_1 _3691_ (.A(_1181_),
    .B(_1184_),
    .C(_1185_),
    .Y(_1186_));
 sg13g2_a21o_1 _3692_ (.A2(_1181_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .B1(_1186_),
    .X(_0108_));
 sg13g2_nor2_1 _3693_ (.A(_1050_),
    .B(_1181_),
    .Y(_1187_));
 sg13g2_a22oi_1 _3694_ (.Y(_0109_),
    .B1(_1187_),
    .B2(_1049_),
    .A2(_1181_),
    .A1(_1450_));
 sg13g2_mux2_1 _3695_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .A1(_1130_),
    .S(_1182_),
    .X(_0110_));
 sg13g2_a21o_2 _3696_ (.A2(_0958_),
    .A1(net579),
    .B1(_1059_),
    .X(_1188_));
 sg13g2_mux2_1 _3697_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .A1(_1188_),
    .S(_1182_),
    .X(_0111_));
 sg13g2_nor2_1 _3698_ (.A(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .B(_1182_),
    .Y(_1189_));
 sg13g2_nor3_1 _3699_ (.A(net22),
    .B(_1063_),
    .C(_1065_),
    .Y(_1190_));
 sg13g2_a21oi_1 _3700_ (.A1(_1182_),
    .A2(_1190_),
    .Y(_0112_),
    .B1(_1189_));
 sg13g2_nand2_1 _3701_ (.Y(_1191_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .B(_1181_));
 sg13g2_o21ai_1 _3702_ (.B1(net580),
    .Y(_1192_),
    .A1(net647),
    .A2(_1001_));
 sg13g2_o21ai_1 _3703_ (.B1(_1192_),
    .Y(_1193_),
    .A1(net581),
    .A2(_1071_));
 sg13g2_o21ai_1 _3704_ (.B1(_1191_),
    .Y(_0113_),
    .A1(_1181_),
    .A2(_1193_));
 sg13g2_nand2b_1 _3705_ (.Y(_1194_),
    .B(_1073_),
    .A_N(net24));
 sg13g2_a21o_2 _3706_ (.A2(_1024_),
    .A1(net578),
    .B1(_1194_),
    .X(_1195_));
 sg13g2_mux2_1 _3707_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .A1(_1195_),
    .S(_1182_),
    .X(_0114_));
 sg13g2_nor3_1 _3708_ (.A(net594),
    .B(_0861_),
    .C(_1040_),
    .Y(_1196_));
 sg13g2_a21o_1 _3709_ (.A2(net595),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .B1(_1196_),
    .X(_0115_));
 sg13g2_nor3_1 _3710_ (.A(net32),
    .B(net594),
    .C(_1144_),
    .Y(_1197_));
 sg13g2_a21oi_1 _3711_ (.A1(_1458_),
    .A2(net594),
    .Y(_0116_),
    .B1(_1197_));
 sg13g2_nand2_1 _3712_ (.Y(_1198_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .B(net595));
 sg13g2_a21oi_1 _3713_ (.A1(_0808_),
    .A2(_0820_),
    .Y(_1199_),
    .B1(_0845_));
 sg13g2_a21o_1 _3714_ (.A2(_1199_),
    .A1(_0850_),
    .B1(_1048_),
    .X(_1200_));
 sg13g2_nor3_1 _3715_ (.A(net19),
    .B(net580),
    .C(_1200_),
    .Y(_1201_));
 sg13g2_o21ai_1 _3716_ (.B1(net645),
    .Y(_1202_),
    .A1(net576),
    .A2(_0898_));
 sg13g2_o21ai_1 _3717_ (.B1(_1198_),
    .Y(_0117_),
    .A1(_1201_),
    .A2(_1202_));
 sg13g2_a21oi_1 _3718_ (.A1(_1975_),
    .A2(_1053_),
    .Y(_1203_),
    .B1(net595));
 sg13g2_a22oi_1 _3719_ (.Y(_1204_),
    .B1(_0921_),
    .B2(_1203_),
    .A2(net595),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ));
 sg13g2_inv_1 _3720_ (.Y(_0118_),
    .A(_1204_));
 sg13g2_nor2_1 _3721_ (.A(net594),
    .B(_1059_),
    .Y(_1205_));
 sg13g2_a22oi_1 _3722_ (.Y(_0119_),
    .B1(_1102_),
    .B2(_1205_),
    .A2(net594),
    .A1(_1472_));
 sg13g2_nand3b_1 _3723_ (.B(net643),
    .C(_1112_),
    .Y(_1206_),
    .A_N(_1133_));
 sg13g2_o21ai_1 _3724_ (.B1(_1206_),
    .Y(_0120_),
    .A1(_1477_),
    .A2(net643));
 sg13g2_nor2_1 _3725_ (.A(net595),
    .B(_1068_),
    .Y(_1207_));
 sg13g2_a22oi_1 _3726_ (.Y(_0121_),
    .B1(_1114_),
    .B2(_1207_),
    .A2(net595),
    .A1(_1485_));
 sg13g2_nor2_1 _3727_ (.A(net594),
    .B(_1194_),
    .Y(_1208_));
 sg13g2_a22oi_1 _3728_ (.Y(_0122_),
    .B1(_1125_),
    .B2(_1208_),
    .A2(net594),
    .A1(_1494_));
 sg13g2_nor2_1 _3729_ (.A(net594),
    .B(_0836_),
    .Y(_1209_));
 sg13g2_nor2_2 _3730_ (.A(net650),
    .B(_1209_),
    .Y(_1210_));
 sg13g2_inv_4 _3731_ (.A(net556),
    .Y(_1211_));
 sg13g2_nor3_1 _3732_ (.A(_1040_),
    .B(_1041_),
    .C(net556),
    .Y(_1212_));
 sg13g2_a21o_1 _3733_ (.A2(net556),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .B1(_1212_),
    .X(_0123_));
 sg13g2_nor3_1 _3734_ (.A(_1184_),
    .B(_1185_),
    .C(net556),
    .Y(_1213_));
 sg13g2_a21o_1 _3735_ (.A2(net556),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .B1(_1213_),
    .X(_0124_));
 sg13g2_nor2_1 _3736_ (.A(_1050_),
    .B(net556),
    .Y(_1214_));
 sg13g2_a22oi_1 _3737_ (.Y(_0125_),
    .B1(_1214_),
    .B2(_1049_),
    .A2(net556),
    .A1(_1449_));
 sg13g2_nand3_1 _3738_ (.B(_1055_),
    .C(_1211_),
    .A(_1054_),
    .Y(_1215_));
 sg13g2_o21ai_1 _3739_ (.B1(_1215_),
    .Y(_0126_),
    .A1(_1442_),
    .A2(_1211_));
 sg13g2_mux2_1 _3740_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .A1(_1188_),
    .S(_1211_),
    .X(_0127_));
 sg13g2_nor3_1 _3741_ (.A(_1133_),
    .B(_1134_),
    .C(net556),
    .Y(_1216_));
 sg13g2_a21o_1 _3742_ (.A2(_1210_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ),
    .B1(_1216_),
    .X(_0128_));
 sg13g2_nor3_1 _3743_ (.A(_1002_),
    .B(_1068_),
    .C(_1210_),
    .Y(_1217_));
 sg13g2_a21oi_1 _3744_ (.A1(_1484_),
    .A2(_1210_),
    .Y(_0129_),
    .B1(_1217_));
 sg13g2_mux2_1 _3745_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .A1(_1195_),
    .S(_1211_),
    .X(_0130_));
 sg13g2_o21ai_1 _3746_ (.B1(net656),
    .Y(_1218_),
    .A1(net575),
    .A2(_0860_));
 sg13g2_nand2b_1 _3747_ (.Y(_1219_),
    .B(_0844_),
    .A_N(_0857_));
 sg13g2_a21o_1 _3748_ (.A2(_0856_),
    .A1(_0744_),
    .B1(_1219_),
    .X(_1220_));
 sg13g2_nor3_1 _3749_ (.A(net9),
    .B(net581),
    .C(_1039_),
    .Y(_1221_));
 sg13g2_a21oi_1 _3750_ (.A1(_1220_),
    .A2(_1221_),
    .Y(_1222_),
    .B1(_1218_));
 sg13g2_a21o_1 _3751_ (.A2(net601),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .B1(_1222_),
    .X(_0131_));
 sg13g2_nand2b_1 _3752_ (.Y(_1223_),
    .B(_0871_),
    .A_N(_0857_));
 sg13g2_nand3_1 _3753_ (.B(_0873_),
    .C(_1223_),
    .A(_0844_),
    .Y(_1224_));
 sg13g2_o21ai_1 _3754_ (.B1(_1045_),
    .Y(_1225_),
    .A1(net10),
    .A2(net666));
 sg13g2_nand3b_1 _3755_ (.B(_1224_),
    .C(_1225_),
    .Y(_1226_),
    .A_N(_1144_));
 sg13g2_mux2_1 _3756_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .A1(_1226_),
    .S(net655),
    .X(_0132_));
 sg13g2_o21ai_1 _3757_ (.B1(_0844_),
    .Y(_1227_),
    .A1(_0873_),
    .A2(_0894_));
 sg13g2_a21oi_1 _3758_ (.A1(_0873_),
    .A2(_0894_),
    .Y(_1228_),
    .B1(_1227_));
 sg13g2_nor3_1 _3759_ (.A(net11),
    .B(net599),
    .C(_1228_),
    .Y(_1229_));
 sg13g2_a22oi_1 _3760_ (.Y(_0133_),
    .B1(_0899_),
    .B2(_1229_),
    .A2(net599),
    .A1(_1448_));
 sg13g2_o21ai_1 _3761_ (.B1(_0916_),
    .Y(_1230_),
    .A1(_0873_),
    .A2(_0894_));
 sg13g2_and3_1 _3762_ (.X(_1231_),
    .A(_0844_),
    .B(_0918_),
    .C(_1230_));
 sg13g2_o21ai_1 _3763_ (.B1(net580),
    .Y(_1232_),
    .A1(net655),
    .A2(_0924_));
 sg13g2_nor2_1 _3764_ (.A(_0920_),
    .B(_1232_),
    .Y(_1233_));
 sg13g2_nor4_1 _3765_ (.A(net12),
    .B(net599),
    .C(_1231_),
    .D(_1233_),
    .Y(_1234_));
 sg13g2_a21oi_1 _3766_ (.A1(_1441_),
    .A2(net600),
    .Y(_0134_),
    .B1(_1234_));
 sg13g2_and2_1 _3767_ (.A(_0918_),
    .B(net552),
    .X(_1235_));
 sg13g2_nor3_1 _3768_ (.A(net574),
    .B(_0955_),
    .C(_1235_),
    .Y(_1236_));
 sg13g2_nor3_1 _3769_ (.A(net13),
    .B(net599),
    .C(_1236_),
    .Y(_1237_));
 sg13g2_a22oi_1 _3770_ (.Y(_0135_),
    .B1(_1102_),
    .B2(_1237_),
    .A2(net598),
    .A1(_1471_));
 sg13g2_xnor2_1 _3771_ (.Y(_1238_),
    .A(_0955_),
    .B(_0969_));
 sg13g2_nor2_1 _3772_ (.A(net574),
    .B(_1238_),
    .Y(_1239_));
 sg13g2_nor3_1 _3773_ (.A(net14),
    .B(net598),
    .C(_1239_),
    .Y(_1240_));
 sg13g2_a22oi_1 _3774_ (.Y(_0136_),
    .B1(_0984_),
    .B2(_1240_),
    .A2(net598),
    .A1(_1476_));
 sg13g2_a21oi_1 _3775_ (.A1(_0955_),
    .A2(_0969_),
    .Y(_1241_),
    .B1(_0994_));
 sg13g2_nor3_1 _3776_ (.A(net574),
    .B(_0997_),
    .C(_1241_),
    .Y(_1242_));
 sg13g2_nor3_1 _3777_ (.A(net15),
    .B(net599),
    .C(_1242_),
    .Y(_1243_));
 sg13g2_a22oi_1 _3778_ (.Y(_0137_),
    .B1(_1114_),
    .B2(_1243_),
    .A2(net601),
    .A1(_1483_));
 sg13g2_xor2_1 _3779_ (.B(_1020_),
    .A(_0997_),
    .X(_1244_));
 sg13g2_nand2b_1 _3780_ (.Y(_1245_),
    .B(net655),
    .A_N(net16));
 sg13g2_a221oi_1 _3781_ (.B2(_0633_),
    .C1(_1074_),
    .B1(_1245_),
    .A1(net661),
    .Y(_1246_),
    .A2(_1244_));
 sg13g2_or2_1 _3782_ (.X(_1247_),
    .B(_1246_),
    .A(net579));
 sg13g2_and2_1 _3783_ (.A(net655),
    .B(_1125_),
    .X(_1248_));
 sg13g2_a22oi_1 _3784_ (.Y(_0138_),
    .B1(_1247_),
    .B2(_1248_),
    .A2(net598),
    .A1(_1493_));
 sg13g2_nor3_1 _3785_ (.A(net600),
    .B(_1040_),
    .C(_1041_),
    .Y(_1249_));
 sg13g2_a21o_1 _3786_ (.A2(net600),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .B1(_1249_),
    .X(_0139_));
 sg13g2_nor3_1 _3787_ (.A(net600),
    .B(_1184_),
    .C(_1185_),
    .Y(_1250_));
 sg13g2_a21o_1 _3788_ (.A2(net600),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .B1(_1250_),
    .X(_0140_));
 sg13g2_nor3_1 _3789_ (.A(net600),
    .B(_1050_),
    .C(_1200_),
    .Y(_1251_));
 sg13g2_a22oi_1 _3790_ (.Y(_0141_),
    .B1(_1049_),
    .B2(_1251_),
    .A2(net600),
    .A1(_1447_));
 sg13g2_and2_1 _3791_ (.A(net656),
    .B(_1055_),
    .X(_1252_));
 sg13g2_a22oi_1 _3792_ (.Y(_1253_),
    .B1(_1054_),
    .B2(_1252_),
    .A2(net600),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ));
 sg13g2_inv_1 _3793_ (.Y(_0142_),
    .A(_1253_));
 sg13g2_nor3_1 _3794_ (.A(net598),
    .B(_0952_),
    .C(_1188_),
    .Y(_1254_));
 sg13g2_a21oi_1 _3795_ (.A1(_1470_),
    .A2(net599),
    .Y(_0143_),
    .B1(_1254_));
 sg13g2_nor3_1 _3796_ (.A(net598),
    .B(_1133_),
    .C(_1134_),
    .Y(_1255_));
 sg13g2_a21o_1 _3797_ (.A2(net599),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .B1(_1255_),
    .X(_0144_));
 sg13g2_nor3_1 _3798_ (.A(net601),
    .B(_1002_),
    .C(_1071_),
    .Y(_1256_));
 sg13g2_a21oi_1 _3799_ (.A1(_1482_),
    .A2(net601),
    .Y(_0145_),
    .B1(_1256_));
 sg13g2_nor3_1 _3800_ (.A(net598),
    .B(_1033_),
    .C(_1195_),
    .Y(_1257_));
 sg13g2_a21oi_1 _3801_ (.A1(_1492_),
    .A2(net598),
    .Y(_0146_),
    .B1(_1257_));
 sg13g2_nor2_1 _3802_ (.A(net608),
    .B(_1038_),
    .Y(_1258_));
 sg13g2_nor3_1 _3803_ (.A(net9),
    .B(_1138_),
    .C(_1258_),
    .Y(_1259_));
 sg13g2_nor3_1 _3804_ (.A(net605),
    .B(_0861_),
    .C(_1259_),
    .Y(_1260_));
 sg13g2_a21o_1 _3805_ (.A2(net604),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ),
    .B1(_1260_),
    .X(_0147_));
 sg13g2_nor2_1 _3806_ (.A(net10),
    .B(_1086_),
    .Y(_1261_));
 sg13g2_a221oi_1 _3807_ (.B2(_1261_),
    .C1(net603),
    .B1(_0884_),
    .A1(net577),
    .Y(_1262_),
    .A2(_0874_));
 sg13g2_a21o_1 _3808_ (.A2(net604),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ),
    .B1(_1262_),
    .X(_0148_));
 sg13g2_nor2_1 _3809_ (.A(net11),
    .B(net603),
    .Y(_1263_));
 sg13g2_a22oi_1 _3810_ (.Y(_0149_),
    .B1(_0901_),
    .B2(_1263_),
    .A2(net603),
    .A1(_1446_));
 sg13g2_nand2_1 _3811_ (.Y(_1264_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .B(net604));
 sg13g2_nand2_1 _3812_ (.Y(_1265_),
    .A(net607),
    .B(_0921_));
 sg13g2_nand2_1 _3813_ (.Y(_1266_),
    .A(net604),
    .B(_0935_));
 sg13g2_nand2b_1 _3814_ (.Y(_1267_),
    .B(net607),
    .A_N(net12));
 sg13g2_a221oi_1 _3815_ (.B2(_0633_),
    .C1(_0929_),
    .B1(_1267_),
    .A1(_0933_),
    .Y(_1268_),
    .A2(_1266_));
 sg13g2_o21ai_1 _3816_ (.B1(_1264_),
    .Y(_0150_),
    .A1(_1265_),
    .A2(_1268_));
 sg13g2_nor2_1 _3817_ (.A(net13),
    .B(net603),
    .Y(_1269_));
 sg13g2_a22oi_1 _3818_ (.Y(_0151_),
    .B1(_1103_),
    .B2(_1269_),
    .A2(net603),
    .A1(_1469_));
 sg13g2_nand2_1 _3819_ (.Y(_1270_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .B(net602));
 sg13g2_nand2_1 _3820_ (.Y(_1271_),
    .A(net606),
    .B(_1112_));
 sg13g2_a21oi_1 _3821_ (.A1(net602),
    .A2(_0975_),
    .Y(_1272_),
    .B1(net583));
 sg13g2_or3_1 _3822_ (.A(net14),
    .B(net661),
    .C(net602),
    .X(_1273_));
 sg13g2_a221oi_1 _3823_ (.B2(_0633_),
    .C1(_1109_),
    .B1(_1273_),
    .A1(_0973_),
    .Y(_1274_),
    .A2(_1272_));
 sg13g2_o21ai_1 _3824_ (.B1(_1270_),
    .Y(_0152_),
    .A1(_1271_),
    .A2(_1274_));
 sg13g2_nor3_1 _3825_ (.A(net15),
    .B(net605),
    .C(_1117_),
    .Y(_1275_));
 sg13g2_a22oi_1 _3826_ (.Y(_0153_),
    .B1(_1114_),
    .B2(_1275_),
    .A2(net605),
    .A1(_1481_));
 sg13g2_nand2_1 _3827_ (.Y(_1276_),
    .A(net585),
    .B(_1027_));
 sg13g2_nor2b_1 _3828_ (.A(net16),
    .B_N(_0687_),
    .Y(_1277_));
 sg13g2_nor3_1 _3829_ (.A(net578),
    .B(_1173_),
    .C(_1277_),
    .Y(_1278_));
 sg13g2_a21oi_1 _3830_ (.A1(_1276_),
    .A2(_1278_),
    .Y(_1279_),
    .B1(net602));
 sg13g2_a22oi_1 _3831_ (.Y(_0154_),
    .B1(_1125_),
    .B2(_1279_),
    .A2(net602),
    .A1(_1491_));
 sg13g2_or2_1 _3832_ (.X(_1280_),
    .B(\sap_3_inst.reg_file.array_serializer_inst.state[1] ),
    .A(\sap_3_inst.reg_file.array_serializer_inst.state[0] ));
 sg13g2_inv_1 _3833_ (.Y(_0155_),
    .A(net764));
 sg13g2_nand2b_2 _3834_ (.Y(_1281_),
    .B(\sap_3_inst.reg_file.array_serializer_inst.state[0] ),
    .A_N(\sap_3_inst.reg_file.array_serializer_inst.state[1] ));
 sg13g2_nor2b_2 _3835_ (.A(\sap_3_inst.reg_file.array_serializer_inst.state[0] ),
    .B_N(\sap_3_inst.reg_file.array_serializer_inst.state[1] ),
    .Y(_1282_));
 sg13g2_nand3_1 _3836_ (.B(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .C(net769),
    .A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .Y(_1283_));
 sg13g2_nand2_1 _3837_ (.Y(_1284_),
    .A(_1282_),
    .B(_1283_));
 sg13g2_nand2_1 _3838_ (.Y(_0156_),
    .A(_1281_),
    .B(_1284_));
 sg13g2_nor2_1 _3839_ (.A(net769),
    .B(_1282_),
    .Y(_1285_));
 sg13g2_a21oi_1 _3840_ (.A1(net769),
    .A2(_0156_),
    .Y(_0157_),
    .B1(_1285_));
 sg13g2_a21oi_1 _3841_ (.A1(net769),
    .A2(_0156_),
    .Y(_1286_),
    .B1(net72));
 sg13g2_nand2_1 _3842_ (.Y(_1287_),
    .A(net63),
    .B(_1281_));
 sg13g2_nand3_1 _3843_ (.B(net769),
    .C(_1282_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .Y(_1288_));
 sg13g2_o21ai_1 _3844_ (.B1(_1281_),
    .Y(_1289_),
    .A1(net63),
    .A2(_1288_));
 sg13g2_nor2_1 _3845_ (.A(_1286_),
    .B(_1289_),
    .Y(_0158_));
 sg13g2_nand2_1 _3846_ (.Y(_0159_),
    .A(_1287_),
    .B(_1288_));
 sg13g2_a21o_1 _3847_ (.A2(regFile_serial_start),
    .A1(net75),
    .B1(_0155_),
    .X(_0160_));
 sg13g2_nor2_1 _3848_ (.A(net66),
    .B(_0156_),
    .Y(_1290_));
 sg13g2_nor2b_1 _3849_ (.A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[0] ),
    .B_N(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .Y(_1291_));
 sg13g2_mux4_1 _3850_ (.S0(net769),
    .A0(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[1] ),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[2] ),
    .A2(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[3] ),
    .A3(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[4] ),
    .S1(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .X(_1292_));
 sg13g2_nand2b_1 _3851_ (.Y(_1293_),
    .B(net769),
    .A_N(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[6] ));
 sg13g2_o21ai_1 _3852_ (.B1(_1293_),
    .Y(_1294_),
    .A1(net769),
    .A2(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[5] ));
 sg13g2_o21ai_1 _3853_ (.B1(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .Y(_1295_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .A2(_1294_));
 sg13g2_a21oi_1 _3854_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[7] ),
    .A2(_1291_),
    .Y(_1296_),
    .B1(_1295_));
 sg13g2_nor2b_1 _3855_ (.A(_1296_),
    .B_N(_1282_),
    .Y(_1297_));
 sg13g2_o21ai_1 _3856_ (.B1(_1297_),
    .Y(_1298_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .A2(_1292_));
 sg13g2_o21ai_1 _3857_ (.B1(_1284_),
    .Y(_1299_),
    .A1(net48),
    .A2(_1281_));
 sg13g2_a21oi_1 _3858_ (.A1(_1298_),
    .A2(_1299_),
    .Y(_0161_),
    .B1(_1290_));
 sg13g2_nand2b_2 _3859_ (.Y(_1300_),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .A_N(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ));
 sg13g2_or2_1 _3860_ (.X(_1301_),
    .B(_1300_),
    .A(_1497_));
 sg13g2_nor2_2 _3861_ (.A(net768),
    .B(_1301_),
    .Y(_1302_));
 sg13g2_nand2b_2 _3862_ (.Y(_1303_),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .A_N(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ));
 sg13g2_or2_1 _3863_ (.X(_1304_),
    .B(_1303_),
    .A(_1497_));
 sg13g2_nor2_2 _3864_ (.A(net768),
    .B(_1304_),
    .Y(_1305_));
 sg13g2_nor4_2 _3865_ (.A(_1497_),
    .B(net768),
    .C(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .Y(_1306_),
    .D(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ));
 sg13g2_nand2_2 _3866_ (.Y(_1307_),
    .A(_1497_),
    .B(net768));
 sg13g2_nor2_2 _3867_ (.A(_1300_),
    .B(_1307_),
    .Y(_1308_));
 sg13g2_nor4_1 _3868_ (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .C(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .D(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .Y(_1309_));
 sg13g2_a21o_2 _3869_ (.A2(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .B1(_1309_),
    .X(_1310_));
 sg13g2_nor3_2 _3870_ (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .B(net768),
    .C(_1303_),
    .Y(_1311_));
 sg13g2_nor3_2 _3871_ (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .B(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .C(_1307_),
    .Y(_1312_));
 sg13g2_nor2_2 _3872_ (.A(_1498_),
    .B(_1301_),
    .Y(_1313_));
 sg13g2_nor2_1 _3873_ (.A(_1498_),
    .B(_1304_),
    .Y(_1314_));
 sg13g2_nor4_1 _3874_ (.A(_1497_),
    .B(_1498_),
    .C(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .D(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .Y(_1315_));
 sg13g2_nor2_2 _3875_ (.A(_1303_),
    .B(_1307_),
    .Y(_1316_));
 sg13g2_nor3_2 _3876_ (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .B(net768),
    .C(_1300_),
    .Y(_1317_));
 sg13g2_a22oi_1 _3877_ (.Y(_1318_),
    .B1(_1308_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ),
    .A2(_1305_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ));
 sg13g2_a22oi_1 _3878_ (.Y(_1319_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .A2(_1306_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ));
 sg13g2_a22oi_1 _3879_ (.Y(_1320_),
    .B1(_1311_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .A2(_1302_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ));
 sg13g2_a22oi_1 _3880_ (.Y(_1321_),
    .B1(net761),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .A2(_1312_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ));
 sg13g2_nand4_1 _3881_ (.B(_1319_),
    .C(_1320_),
    .A(_1318_),
    .Y(_1322_),
    .D(_1321_));
 sg13g2_a21oi_1 _3882_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .A2(_1317_),
    .Y(_1323_),
    .B1(net762));
 sg13g2_nand2b_1 _3883_ (.Y(_1324_),
    .B(_1323_),
    .A_N(_1322_));
 sg13g2_a221oi_1 _3884_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .C1(_1324_),
    .B1(net721),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .Y(_1325_),
    .A2(_1313_));
 sg13g2_a21o_1 _3885_ (.A2(net762),
    .A1(_1460_),
    .B1(net765),
    .X(_1326_));
 sg13g2_nand2_1 _3886_ (.Y(_1327_),
    .A(net48),
    .B(net764));
 sg13g2_o21ai_1 _3887_ (.B1(_1327_),
    .Y(_0162_),
    .A1(_1325_),
    .A2(_1326_));
 sg13g2_a22oi_1 _3888_ (.Y(_1328_),
    .B1(_1313_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .A2(_1308_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ));
 sg13g2_a21oi_1 _3889_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .A2(_1305_),
    .Y(_1329_),
    .B1(net762));
 sg13g2_a22oi_1 _3890_ (.Y(_1330_),
    .B1(_1312_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .A2(_1311_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ));
 sg13g2_a22oi_1 _3891_ (.Y(_1331_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .A2(net721),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ));
 sg13g2_a22oi_1 _3892_ (.Y(_1332_),
    .B1(net761),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .A2(_1302_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ));
 sg13g2_nand4_1 _3893_ (.B(_1330_),
    .C(_1331_),
    .A(_1329_),
    .Y(_1333_),
    .D(_1332_));
 sg13g2_a221oi_1 _3894_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .C1(_1333_),
    .B1(_1317_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .Y(_1334_),
    .A2(_1306_));
 sg13g2_a221oi_1 _3895_ (.B2(_1334_),
    .C1(net765),
    .B1(_1328_),
    .A1(_1457_),
    .Y(_1335_),
    .A2(net762));
 sg13g2_a21o_1 _3896_ (.A2(net764),
    .A1(net53),
    .B1(_1335_),
    .X(_0163_));
 sg13g2_a22oi_1 _3897_ (.Y(_1336_),
    .B1(_1317_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .A2(_1302_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ));
 sg13g2_a22oi_1 _3898_ (.Y(_1337_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .A2(_1311_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ));
 sg13g2_a21oi_1 _3899_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .A2(_1308_),
    .Y(_1338_),
    .B1(net762));
 sg13g2_a22oi_1 _3900_ (.Y(_1339_),
    .B1(net761),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ),
    .A2(net721),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ));
 sg13g2_a22oi_1 _3901_ (.Y(_1340_),
    .B1(_1313_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .A2(_1305_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ));
 sg13g2_nand4_1 _3902_ (.B(_1338_),
    .C(_1339_),
    .A(_1337_),
    .Y(_1341_),
    .D(_1340_));
 sg13g2_a221oi_1 _3903_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .C1(_1341_),
    .B1(_1312_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .Y(_1342_),
    .A2(_1306_));
 sg13g2_a221oi_1 _3904_ (.B2(_1342_),
    .C1(net765),
    .B1(_1336_),
    .A1(_1444_),
    .Y(_1343_),
    .A2(net762));
 sg13g2_a21o_1 _3905_ (.A2(net764),
    .A1(net54),
    .B1(_1343_),
    .X(_0164_));
 sg13g2_a22oi_1 _3906_ (.Y(_1344_),
    .B1(_1317_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .A2(_1312_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ));
 sg13g2_a21oi_1 _3907_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .A2(_1316_),
    .Y(_1345_),
    .B1(net762));
 sg13g2_a22oi_1 _3908_ (.Y(_1346_),
    .B1(_1313_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .A2(_1311_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ));
 sg13g2_a22oi_1 _3909_ (.Y(_1347_),
    .B1(net761),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .A2(net721),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ));
 sg13g2_a22oi_1 _3910_ (.Y(_1348_),
    .B1(_1306_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .A2(_1302_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ));
 sg13g2_nand4_1 _3911_ (.B(_1346_),
    .C(_1347_),
    .A(_1345_),
    .Y(_1349_),
    .D(_1348_));
 sg13g2_a221oi_1 _3912_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .C1(_1349_),
    .B1(_1308_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .Y(_1350_),
    .A2(_1305_));
 sg13g2_a221oi_1 _3913_ (.B2(_1350_),
    .C1(net764),
    .B1(_1344_),
    .A1(_1440_),
    .Y(_1351_),
    .A2(net762));
 sg13g2_a21o_1 _3914_ (.A2(net764),
    .A1(net51),
    .B1(_1351_),
    .X(_0165_));
 sg13g2_a22oi_1 _3915_ (.Y(_1352_),
    .B1(net761),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .A2(_1305_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ));
 sg13g2_a22oi_1 _3916_ (.Y(_1353_),
    .B1(net721),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .A2(_1308_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ));
 sg13g2_a22oi_1 _3917_ (.Y(_1354_),
    .B1(_1317_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .A2(_1312_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ));
 sg13g2_a21oi_1 _3918_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .A2(_1302_),
    .Y(_1355_),
    .B1(net763));
 sg13g2_a22oi_1 _3919_ (.Y(_1356_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .A2(_1311_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ));
 sg13g2_nand4_1 _3920_ (.B(_1354_),
    .C(_1355_),
    .A(_1352_),
    .Y(_1357_),
    .D(_1356_));
 sg13g2_a221oi_1 _3921_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .C1(_1357_),
    .B1(_1313_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .Y(_1358_),
    .A2(_1306_));
 sg13g2_a221oi_1 _3922_ (.B2(_1358_),
    .C1(net765),
    .B1(_1353_),
    .A1(_1468_),
    .Y(_1359_),
    .A2(net763));
 sg13g2_a21o_1 _3923_ (.A2(net764),
    .A1(net49),
    .B1(_1359_),
    .X(_0166_));
 sg13g2_a22oi_1 _3924_ (.Y(_1360_),
    .B1(_1308_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .A2(_1306_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ));
 sg13g2_a22oi_1 _3925_ (.Y(_1361_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .A2(net721),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ));
 sg13g2_a21oi_1 _3926_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .A2(net761),
    .Y(_1362_),
    .B1(net763));
 sg13g2_a22oi_1 _3927_ (.Y(_1363_),
    .B1(_1313_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .A2(_1311_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ));
 sg13g2_a22oi_1 _3928_ (.Y(_1364_),
    .B1(_1305_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .A2(_1302_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ));
 sg13g2_nand4_1 _3929_ (.B(_1362_),
    .C(_1363_),
    .A(_1361_),
    .Y(_1365_),
    .D(_1364_));
 sg13g2_a221oi_1 _3930_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .C1(_1365_),
    .B1(_1317_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .Y(_1366_),
    .A2(_1312_));
 sg13g2_a221oi_1 _3931_ (.B2(_1366_),
    .C1(net765),
    .B1(_1360_),
    .A1(_1475_),
    .Y(_1367_),
    .A2(net763));
 sg13g2_a21o_1 _3932_ (.A2(net764),
    .A1(net55),
    .B1(_1367_),
    .X(_0167_));
 sg13g2_a21oi_1 _3933_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .A2(_1311_),
    .Y(_1368_),
    .B1(net763));
 sg13g2_a22oi_1 _3934_ (.Y(_1369_),
    .B1(_1315_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .A2(_1306_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ));
 sg13g2_a22oi_1 _3935_ (.Y(_1370_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .A2(_1313_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ));
 sg13g2_a22oi_1 _3936_ (.Y(_1371_),
    .B1(_1317_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .A2(_1308_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ));
 sg13g2_a22oi_1 _3937_ (.Y(_1372_),
    .B1(_1305_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .A2(_1302_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ));
 sg13g2_nand4_1 _3938_ (.B(_1370_),
    .C(_1371_),
    .A(_1368_),
    .Y(_1373_),
    .D(_1372_));
 sg13g2_a221oi_1 _3939_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .C1(_1373_),
    .B1(_1314_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .Y(_1374_),
    .A2(_1312_));
 sg13g2_a221oi_1 _3940_ (.B2(_1374_),
    .C1(net765),
    .B1(_1369_),
    .A1(_1479_),
    .Y(_1375_),
    .A2(_1310_));
 sg13g2_a21o_1 _3941_ (.A2(_1280_),
    .A1(net50),
    .B1(_1375_),
    .X(_0168_));
 sg13g2_a22oi_1 _3942_ (.Y(_1376_),
    .B1(net761),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .A2(_1306_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ));
 sg13g2_a22oi_1 _3943_ (.Y(_1377_),
    .B1(_1316_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .A2(_1312_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ));
 sg13g2_a21oi_1 _3944_ (.A1(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .A2(_1317_),
    .Y(_1378_),
    .B1(net763));
 sg13g2_a22oi_1 _3945_ (.Y(_1379_),
    .B1(_1313_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .A2(_1305_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ));
 sg13g2_a22oi_1 _3946_ (.Y(_1380_),
    .B1(_1311_),
    .B2(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .A2(_1302_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ));
 sg13g2_nand4_1 _3947_ (.B(_1377_),
    .C(_1378_),
    .A(_1376_),
    .Y(_1381_),
    .D(_1380_));
 sg13g2_a221oi_1 _3948_ (.B2(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .C1(_1381_),
    .B1(net721),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ),
    .Y(_1382_),
    .A2(_1308_));
 sg13g2_a221oi_1 _3949_ (.B2(_1382_),
    .C1(net765),
    .B1(_1379_),
    .A1(_1490_),
    .Y(_1383_),
    .A2(net763));
 sg13g2_a21o_1 _3950_ (.A2(_1280_),
    .A1(net52),
    .B1(_1383_),
    .X(_0169_));
 sg13g2_nor3_1 _3951_ (.A(net604),
    .B(_1040_),
    .C(_1041_),
    .Y(_1384_));
 sg13g2_a21o_1 _3952_ (.A2(net604),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .B1(_1384_),
    .X(_0170_));
 sg13g2_mux2_1 _3953_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .A1(_1047_),
    .S(net609),
    .X(_0171_));
 sg13g2_a21oi_1 _3954_ (.A1(net580),
    .A2(_0906_),
    .Y(_1385_),
    .B1(net604));
 sg13g2_nand2b_1 _3955_ (.Y(_1386_),
    .B(_1385_),
    .A_N(_1201_));
 sg13g2_o21ai_1 _3956_ (.B1(_1386_),
    .Y(_0172_),
    .A1(_1445_),
    .A2(net608));
 sg13g2_mux2_1 _3957_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .A1(_1130_),
    .S(net608),
    .X(_0173_));
 sg13g2_mux2_1 _3958_ (.A0(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .A1(_1188_),
    .S(net607),
    .X(_0174_));
 sg13g2_nand2_1 _3959_ (.Y(_1387_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .B(net602));
 sg13g2_o21ai_1 _3960_ (.B1(_1387_),
    .Y(_0175_),
    .A1(net603),
    .A2(_1190_));
 sg13g2_nor3_1 _3961_ (.A(net604),
    .B(_1002_),
    .C(_1068_),
    .Y(_1388_));
 sg13g2_a21oi_1 _3962_ (.A1(_1480_),
    .A2(net605),
    .Y(_0176_),
    .B1(_1388_));
 sg13g2_nor3_1 _3963_ (.A(net602),
    .B(_1025_),
    .C(_1075_),
    .Y(_1389_));
 sg13g2_a21o_1 _3964_ (.A2(net602),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .B1(_1389_),
    .X(_0177_));
 sg13g2_nand3_1 _3965_ (.B(_0299_),
    .C(_0301_),
    .A(net683),
    .Y(_1390_));
 sg13g2_nand2b_1 _3966_ (.Y(_1391_),
    .B(_1390_),
    .A_N(_1845_));
 sg13g2_nand2b_1 _3967_ (.Y(_1392_),
    .B(net617),
    .A_N(net664));
 sg13g2_nand2_1 _3968_ (.Y(_1393_),
    .A(_1938_),
    .B(_0315_));
 sg13g2_nand3_1 _3969_ (.B(_1392_),
    .C(_1393_),
    .A(_0311_),
    .Y(_1394_));
 sg13g2_mux2_1 _3970_ (.A0(_0321_),
    .A1(net759),
    .S(net664),
    .X(_1395_));
 sg13g2_nor2_1 _3971_ (.A(net549),
    .B(_1395_),
    .Y(_1396_));
 sg13g2_a21oi_1 _3972_ (.A1(_1462_),
    .A2(net549),
    .Y(_0178_),
    .B1(_1396_));
 sg13g2_mux2_1 _3973_ (.A0(_0358_),
    .A1(net758),
    .S(net664),
    .X(_1397_));
 sg13g2_mux2_1 _3974_ (.A0(_1397_),
    .A1(\sap_3_inst.alu.act[1] ),
    .S(net549),
    .X(_0179_));
 sg13g2_mux2_1 _3975_ (.A0(_0391_),
    .A1(net755),
    .S(net663),
    .X(_1398_));
 sg13g2_mux2_1 _3976_ (.A0(_1398_),
    .A1(\sap_3_inst.alu.act[2] ),
    .S(net548),
    .X(_0180_));
 sg13g2_nor2_1 _3977_ (.A(_0431_),
    .B(net664),
    .Y(_1399_));
 sg13g2_a21oi_1 _3978_ (.A1(net753),
    .A2(net663),
    .Y(_1400_),
    .B1(_1399_));
 sg13g2_nand2_1 _3979_ (.Y(_1401_),
    .A(\sap_3_inst.alu.act[3] ),
    .B(net548));
 sg13g2_o21ai_1 _3980_ (.B1(_1401_),
    .Y(_0181_),
    .A1(net548),
    .A2(_1400_));
 sg13g2_mux2_1 _3981_ (.A0(_0458_),
    .A1(net750),
    .S(net663),
    .X(_1402_));
 sg13g2_mux2_1 _3982_ (.A0(_1402_),
    .A1(\sap_3_inst.alu.act[4] ),
    .S(net548),
    .X(_0182_));
 sg13g2_mux2_1 _3983_ (.A0(_0488_),
    .A1(net748),
    .S(net663),
    .X(_1403_));
 sg13g2_mux2_1 _3984_ (.A0(_1403_),
    .A1(\sap_3_inst.alu.act[5] ),
    .S(net548),
    .X(_0183_));
 sg13g2_nor2_1 _3985_ (.A(_0510_),
    .B(net663),
    .Y(_1404_));
 sg13g2_a21oi_1 _3986_ (.A1(net746),
    .A2(net663),
    .Y(_1405_),
    .B1(_1404_));
 sg13g2_nand2_1 _3987_ (.Y(_1406_),
    .A(\sap_3_inst.alu.act[6] ),
    .B(net548));
 sg13g2_o21ai_1 _3988_ (.B1(_1406_),
    .Y(_0184_),
    .A1(net548),
    .A2(_1405_));
 sg13g2_nand2_1 _3989_ (.Y(_1407_),
    .A(\sap_3_inst.alu.act[7] ),
    .B(net548));
 sg13g2_nor2_1 _3990_ (.A(_0542_),
    .B(net663),
    .Y(_1408_));
 sg13g2_a21oi_1 _3991_ (.A1(net744),
    .A2(net663),
    .Y(_1409_),
    .B1(_1408_));
 sg13g2_o21ai_1 _3992_ (.B1(_1407_),
    .Y(_0185_),
    .A1(net549),
    .A2(_1409_));
 sg13g2_nor2_2 _3993_ (.A(\u_ser.state[0] ),
    .B(_1433_),
    .Y(_1410_));
 sg13g2_nand2_1 _3994_ (.Y(_1411_),
    .A(\u_ser.bit_pos[1] ),
    .B(net767));
 sg13g2_nand2_1 _3995_ (.Y(_1412_),
    .A(_1410_),
    .B(_1411_));
 sg13g2_o21ai_1 _3996_ (.B1(_1410_),
    .Y(_1413_),
    .A1(_1434_),
    .A2(_1411_));
 sg13g2_o21ai_1 _3997_ (.B1(_1413_),
    .Y(_0187_),
    .A1(_1432_),
    .A2(\u_ser.state[1] ));
 sg13g2_nand3b_1 _3998_ (.B(\u_ser.shadow_reg[7] ),
    .C(\u_ser.bit_pos[1] ),
    .Y(_1414_),
    .A_N(net767));
 sg13g2_nand2b_1 _3999_ (.Y(_1415_),
    .B(net767),
    .A_N(\u_ser.shadow_reg[6] ));
 sg13g2_o21ai_1 _4000_ (.B1(_1415_),
    .Y(_1416_),
    .A1(\u_ser.bit_pos[0] ),
    .A2(\u_ser.shadow_reg[5] ));
 sg13g2_o21ai_1 _4001_ (.B1(_1414_),
    .Y(_1417_),
    .A1(\u_ser.bit_pos[1] ),
    .A2(_1416_));
 sg13g2_nand3_1 _4002_ (.B(_1410_),
    .C(_1417_),
    .A(\u_ser.bit_pos[2] ),
    .Y(_1418_));
 sg13g2_mux4_1 _4003_ (.S0(net767),
    .A0(\u_ser.shadow_reg[1] ),
    .A1(\u_ser.shadow_reg[2] ),
    .A2(\u_ser.shadow_reg[3] ),
    .A3(\u_ser.shadow_reg[4] ),
    .S1(\u_ser.bit_pos[1] ),
    .X(_1419_));
 sg13g2_nand3_1 _4004_ (.B(_1410_),
    .C(_1419_),
    .A(_1434_),
    .Y(_1420_));
 sg13g2_o21ai_1 _4005_ (.B1(\u_ser.shadow_reg[0] ),
    .Y(_1421_),
    .A1(\u_ser.state[0] ),
    .A2(_1433_));
 sg13g2_nand4_1 _4006_ (.B(_1418_),
    .C(_1420_),
    .A(_0187_),
    .Y(_1422_),
    .D(_1421_));
 sg13g2_o21ai_1 _4007_ (.B1(_1422_),
    .Y(_1423_),
    .A1(net77),
    .A2(_0187_));
 sg13g2_inv_1 _4008_ (.Y(_0188_),
    .A(_1423_));
 sg13g2_a21o_1 _4009_ (.A2(net68),
    .A1(\u_ser.state[1] ),
    .B1(net766),
    .X(_0189_));
 sg13g2_nor2_2 _4010_ (.A(_1435_),
    .B(_1288_),
    .Y(_1424_));
 sg13g2_xnor2_1 _4011_ (.Y(_0190_),
    .A(_1497_),
    .B(_1424_));
 sg13g2_nand3_1 _4012_ (.B(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .C(_1424_),
    .A(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .Y(_1425_));
 sg13g2_a21o_1 _4013_ (.A2(_1424_),
    .A1(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .B1(net768),
    .X(_1426_));
 sg13g2_and2_1 _4014_ (.A(_1425_),
    .B(_1426_),
    .X(_0191_));
 sg13g2_a22oi_1 _4015_ (.Y(_1427_),
    .B1(_1425_),
    .B2(net79),
    .A2(_1424_),
    .A1(net761));
 sg13g2_inv_1 _4016_ (.Y(_0192_),
    .A(_1427_));
 sg13g2_a22oi_1 _4017_ (.Y(_1428_),
    .B1(_1425_),
    .B2(net78),
    .A2(_1424_),
    .A1(net721));
 sg13g2_inv_1 _4018_ (.Y(_0193_),
    .A(_1428_));
 sg13g2_nor2_1 _4019_ (.A(net767),
    .B(_1410_),
    .Y(_1429_));
 sg13g2_a21oi_1 _4020_ (.A1(net767),
    .A2(_0187_),
    .Y(_0194_),
    .B1(_1429_));
 sg13g2_a21oi_1 _4021_ (.A1(net767),
    .A2(_0187_),
    .Y(_1430_),
    .B1(net71));
 sg13g2_a21oi_1 _4022_ (.A1(_1412_),
    .A2(_0187_),
    .Y(_0195_),
    .B1(_1430_));
 sg13g2_nand3_1 _4023_ (.B(net767),
    .C(_1410_),
    .A(\u_ser.bit_pos[1] ),
    .Y(_1431_));
 sg13g2_a22oi_1 _4024_ (.Y(_0196_),
    .B1(_1434_),
    .B2(_1431_),
    .A2(_1433_),
    .A1(net58));
 sg13g2_inv_1 _4026__4 (.Y(net38),
    .A(\clknet_leaf_2_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4027__5 (.Y(net39),
    .A(\clknet_leaf_2_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4028__6 (.Y(net40),
    .A(\clknet_leaf_0_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4029__7 (.Y(net41),
    .A(\clknet_leaf_0_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4030__8 (.Y(net42),
    .A(\clknet_leaf_3_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4031__9 (.Y(net43),
    .A(\clknet_leaf_3_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4032__10 (.Y(net44),
    .A(\clknet_leaf_1_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4033__11 (.Y(net45),
    .A(\clknet_leaf_1_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4034__12 (.Y(net46),
    .A(\clknet_leaf_1_sap_3_inst.alu.clk ));
 sg13g2_inv_1 _4035__13 (.Y(net47),
    .A(\clknet_leaf_1_sap_3_inst.alu.clk ));
 sg13g2_buf_8 clkbuf_regs_0_clk_div_two (.A(\sap_3_inst.alu.clk ),
    .X(\sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4036_ (.RESET_B(net783),
    .D(_0018_),
    .Q(\u_ser.shadow_reg[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _4037_ (.RESET_B(net784),
    .D(_0019_),
    .Q(\u_ser.shadow_reg[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _4038_ (.RESET_B(net784),
    .D(_0020_),
    .Q(\u_ser.shadow_reg[2] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4039_ (.RESET_B(net784),
    .D(_0021_),
    .Q(\u_ser.shadow_reg[3] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _4040_ (.RESET_B(net788),
    .D(_0022_),
    .Q(\u_ser.shadow_reg[4] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4041_ (.RESET_B(net788),
    .D(_0023_),
    .Q(\u_ser.shadow_reg[5] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4042_ (.RESET_B(net788),
    .D(_0024_),
    .Q(\u_ser.shadow_reg[6] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4043_ (.RESET_B(net788),
    .D(_0025_),
    .Q(\u_ser.shadow_reg[7] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4044_ (.RESET_B(net786),
    .D(_0026_),
    .Q(\sap_3_inst.alu.flags[0] ),
    .CLK(net36));
 sg13g2_dfrbpq_1 _4045_ (.RESET_B(net783),
    .D(_0027_),
    .Q(\sap_3_inst.alu.flags[1] ),
    .CLK(net37));
 sg13g2_dfrbpq_1 _4046_ (.RESET_B(net786),
    .D(_0028_),
    .Q(\sap_3_inst.alu.flags[2] ),
    .CLK(net38));
 sg13g2_dfrbpq_1 _4047_ (.RESET_B(net786),
    .D(_0029_),
    .Q(\sap_3_inst.alu.flags[3] ),
    .CLK(net39));
 sg13g2_dfrbpq_2 _4048_ (.RESET_B(net770),
    .D(_0002_),
    .Q(\sap_3_inst.controller.stage[0] ),
    .CLK(net40));
 sg13g2_dfrbpq_2 _4049_ (.RESET_B(net772),
    .D(_0003_),
    .Q(\sap_3_inst.controller.stage[1] ),
    .CLK(net41));
 sg13g2_dfrbpq_2 _4050_ (.RESET_B(net772),
    .D(_0004_),
    .Q(\sap_3_inst.controller.stage[2] ),
    .CLK(net42));
 sg13g2_dfrbpq_2 _4051_ (.RESET_B(net772),
    .D(_0005_),
    .Q(\sap_3_inst.controller.stage[3] ),
    .CLK(net43));
 sg13g2_dfrbpq_1 _4052_ (.RESET_B(net787),
    .D(_0030_),
    .Q(\sap_3_inst.alu.flags[4] ),
    .CLK(net44));
 sg13g2_dfrbpq_1 _4053_ (.RESET_B(net787),
    .D(_0031_),
    .Q(\sap_3_inst.alu.flags[5] ),
    .CLK(net45));
 sg13g2_dfrbpq_1 _4054_ (.RESET_B(net793),
    .D(_0032_),
    .Q(\sap_3_inst.alu.flags[6] ),
    .CLK(net46));
 sg13g2_dfrbpq_1 _4055_ (.RESET_B(net799),
    .D(_0033_),
    .Q(\sap_3_inst.alu.flags[7] ),
    .CLK(net47));
 sg13g2_dfrbpq_1 _4056_ (.RESET_B(net785),
    .D(_0034_),
    .Q(\sap_3_inst.alu.acc[0] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4057_ (.RESET_B(net784),
    .D(_0035_),
    .Q(\sap_3_inst.alu.acc[1] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4058_ (.RESET_B(net790),
    .D(_0036_),
    .Q(\sap_3_inst.alu.acc[2] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4059_ (.RESET_B(net789),
    .D(_0037_),
    .Q(\sap_3_inst.alu.acc[3] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4060_ (.RESET_B(net790),
    .D(_0038_),
    .Q(\sap_3_inst.alu.acc[4] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4061_ (.RESET_B(net790),
    .D(_0039_),
    .Q(\sap_3_inst.alu.acc[5] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4062_ (.RESET_B(net791),
    .D(_0040_),
    .Q(\sap_3_inst.alu.acc[6] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4063_ (.RESET_B(net791),
    .D(_0041_),
    .Q(\sap_3_inst.alu.acc[7] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4064_ (.RESET_B(net783),
    .D(_0042_),
    .Q(\sap_3_inst.out[0] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4065_ (.RESET_B(net783),
    .D(_0043_),
    .Q(\sap_3_inst.out[1] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4066_ (.RESET_B(net784),
    .D(_0044_),
    .Q(\sap_3_inst.out[2] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4067_ (.RESET_B(net784),
    .D(_0045_),
    .Q(\sap_3_inst.out[3] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4068_ (.RESET_B(net789),
    .D(_0046_),
    .Q(\sap_3_inst.out[4] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4069_ (.RESET_B(net789),
    .D(_0047_),
    .Q(\sap_3_inst.out[5] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4070_ (.RESET_B(net789),
    .D(_0048_),
    .Q(\sap_3_inst.out[6] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4071_ (.RESET_B(net788),
    .D(_0049_),
    .Q(\sap_3_inst.out[7] ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4072_ (.RESET_B(net787),
    .D(_0050_),
    .Q(\sap_3_inst.alu.carry ),
    .CLK(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4073_ (.RESET_B(net785),
    .D(_0051_),
    .Q(\sap_3_inst.alu.tmp[0] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4074_ (.RESET_B(net785),
    .D(_0052_),
    .Q(\sap_3_inst.alu.tmp[1] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4075_ (.RESET_B(net789),
    .D(_0053_),
    .Q(\sap_3_inst.alu.tmp[2] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4076_ (.RESET_B(net789),
    .D(_0054_),
    .Q(\sap_3_inst.alu.tmp[3] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4077_ (.RESET_B(net790),
    .D(_0055_),
    .Q(\sap_3_inst.alu.tmp[4] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4078_ (.RESET_B(net791),
    .D(_0056_),
    .Q(\sap_3_inst.alu.tmp[5] ),
    .CLK(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4079_ (.RESET_B(net791),
    .D(_0057_),
    .Q(\sap_3_inst.alu.tmp[6] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4080_ (.RESET_B(net791),
    .D(_0058_),
    .Q(\sap_3_inst.alu.tmp[7] ),
    .CLK(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4081_ (.RESET_B(net770),
    .D(_0059_),
    .Q(\sap_3_inst.controller.opcode[0] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4082_ (.RESET_B(net785),
    .D(_0060_),
    .Q(\sap_3_inst.controller.opcode[1] ),
    .CLK(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4083_ (.RESET_B(net770),
    .D(_0061_),
    .Q(\sap_3_inst.controller.opcode[2] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4084_ (.RESET_B(net770),
    .D(_0062_),
    .Q(\sap_3_inst.controller.opcode[3] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4085_ (.RESET_B(net770),
    .D(_0063_),
    .Q(\sap_3_inst.controller.opcode[4] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4086_ (.RESET_B(net771),
    .D(_0064_),
    .Q(\sap_3_inst.controller.opcode[5] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4087_ (.RESET_B(net770),
    .D(_0065_),
    .Q(\sap_3_inst.controller.opcode[6] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4088_ (.RESET_B(net772),
    .D(_0066_),
    .Q(\sap_3_inst.controller.opcode[7] ),
    .CLK(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4089_ (.RESET_B(net782),
    .D(_0067_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][0] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4090_ (.RESET_B(net778),
    .D(_0068_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][1] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4091_ (.RESET_B(net774),
    .D(_0069_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][2] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4092_ (.RESET_B(net782),
    .D(_0070_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][3] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4093_ (.RESET_B(net774),
    .D(_0071_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][4] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4094_ (.RESET_B(net778),
    .D(_0072_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][5] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4095_ (.RESET_B(net780),
    .D(_0073_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][6] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4096_ (.RESET_B(net775),
    .D(_0074_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[0][7] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4097_ (.RESET_B(net797),
    .D(_0075_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][0] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4098_ (.RESET_B(net786),
    .D(_0076_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][1] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4099_ (.RESET_B(net786),
    .D(_0077_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][2] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4100_ (.RESET_B(net793),
    .D(_0078_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][3] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4101_ (.RESET_B(net776),
    .D(_0079_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][4] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4102_ (.RESET_B(net776),
    .D(_0080_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][5] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4103_ (.RESET_B(net797),
    .D(_0081_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][6] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4104_ (.RESET_B(net775),
    .D(_0082_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[1][7] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4105_ (.RESET_B(net795),
    .D(_0083_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][0] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4106_ (.RESET_B(net770),
    .D(_0084_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4107_ (.RESET_B(net771),
    .D(_0085_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][2] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4108_ (.RESET_B(net782),
    .D(_0086_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][3] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4109_ (.RESET_B(net774),
    .D(_0087_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][4] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4110_ (.RESET_B(net776),
    .D(_0088_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][5] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4111_ (.RESET_B(net780),
    .D(_0089_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][6] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4112_ (.RESET_B(net775),
    .D(_0090_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[2][7] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4113_ (.RESET_B(net796),
    .D(_0091_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][0] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4114_ (.RESET_B(net793),
    .D(_0092_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][1] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4115_ (.RESET_B(net795),
    .D(_0093_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][2] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4116_ (.RESET_B(net793),
    .D(_0094_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][3] ),
    .CLK(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4117_ (.RESET_B(net776),
    .D(_0095_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][4] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4118_ (.RESET_B(net776),
    .D(_0096_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][5] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4119_ (.RESET_B(net796),
    .D(_0097_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][6] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4120_ (.RESET_B(net775),
    .D(_0098_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[3][7] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4121_ (.RESET_B(net795),
    .D(_0099_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][0] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4122_ (.RESET_B(net773),
    .D(_0100_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][1] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4123_ (.RESET_B(net771),
    .D(_0101_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][2] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4124_ (.RESET_B(net782),
    .D(_0102_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][3] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4125_ (.RESET_B(net774),
    .D(_0103_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][4] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4126_ (.RESET_B(net777),
    .D(_0104_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][5] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4127_ (.RESET_B(net780),
    .D(_0105_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][6] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4128_ (.RESET_B(net775),
    .D(_0106_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[4][7] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4129_ (.RESET_B(net796),
    .D(_0107_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][0] ),
    .CLK(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4130_ (.RESET_B(net773),
    .D(_0108_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][1] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4131_ (.RESET_B(net786),
    .D(_0109_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][2] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4132_ (.RESET_B(net795),
    .D(_0110_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][3] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4133_ (.RESET_B(net779),
    .D(_0111_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][4] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4134_ (.RESET_B(net779),
    .D(_0112_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][5] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4135_ (.RESET_B(net796),
    .D(_0113_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][6] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4136_ (.RESET_B(net779),
    .D(_0114_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[5][7] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4137_ (.RESET_B(net796),
    .D(_0115_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][0] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4138_ (.RESET_B(net773),
    .D(_0116_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][1] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4139_ (.RESET_B(net773),
    .D(_0117_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][2] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4140_ (.RESET_B(net795),
    .D(_0118_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][3] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4141_ (.RESET_B(net774),
    .D(_0119_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][4] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4142_ (.RESET_B(net776),
    .D(_0120_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][5] ),
    .CLK(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4143_ (.RESET_B(net780),
    .D(_0121_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][6] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4144_ (.RESET_B(net777),
    .D(_0122_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[6][7] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4145_ (.RESET_B(net796),
    .D(_0123_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][0] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4146_ (.RESET_B(net773),
    .D(_0124_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][1] ),
    .CLK(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4147_ (.RESET_B(net793),
    .D(_0125_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][2] ),
    .CLK(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4148_ (.RESET_B(net795),
    .D(_0126_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][3] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4149_ (.RESET_B(net779),
    .D(_0127_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][4] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4150_ (.RESET_B(net779),
    .D(_0128_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][5] ),
    .CLK(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4151_ (.RESET_B(net780),
    .D(_0129_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][6] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4152_ (.RESET_B(net779),
    .D(_0130_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[7][7] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4153_ (.RESET_B(net795),
    .D(_0131_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][0] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4154_ (.RESET_B(net770),
    .D(_0132_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][1] ),
    .CLK(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4155_ (.RESET_B(net774),
    .D(_0133_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][2] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4156_ (.RESET_B(net782),
    .D(_0134_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][3] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4157_ (.RESET_B(net774),
    .D(_0135_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][4] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4158_ (.RESET_B(net775),
    .D(_0136_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][5] ),
    .CLK(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4159_ (.RESET_B(net781),
    .D(_0137_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][6] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4160_ (.RESET_B(net775),
    .D(_0138_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[8][7] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4161_ (.RESET_B(net796),
    .D(_0139_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][0] ),
    .CLK(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4162_ (.RESET_B(net786),
    .D(_0140_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][1] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4163_ (.RESET_B(net786),
    .D(_0141_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][2] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4164_ (.RESET_B(net794),
    .D(_0142_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][3] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4165_ (.RESET_B(net779),
    .D(_0143_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][4] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4166_ (.RESET_B(net776),
    .D(_0144_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][5] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4167_ (.RESET_B(net780),
    .D(_0145_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][6] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4168_ (.RESET_B(net776),
    .D(_0146_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[9][7] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4169_ (.RESET_B(net795),
    .D(_0147_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][0] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4170_ (.RESET_B(net773),
    .D(_0148_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][1] ),
    .CLK(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4171_ (.RESET_B(net771),
    .D(_0149_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][2] ),
    .CLK(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4172_ (.RESET_B(net782),
    .D(_0150_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][3] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4173_ (.RESET_B(net774),
    .D(_0151_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][4] ),
    .CLK(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4174_ (.RESET_B(net777),
    .D(_0152_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][5] ),
    .CLK(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4175_ (.RESET_B(net780),
    .D(_0153_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][6] ),
    .CLK(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4176_ (.RESET_B(net777),
    .D(_0154_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[10][7] ),
    .CLK(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4177_ (.RESET_B(net799),
    .D(_0155_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.state[0] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _4178_ (.RESET_B(net799),
    .D(_0156_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.state[1] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4179_ (.RESET_B(net799),
    .D(net81),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[0] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _4180_ (.RESET_B(net799),
    .D(net73),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _4181_ (.RESET_B(net799),
    .D(net64),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4182_ (.RESET_B(net799),
    .D(net76),
    .Q(regFile_serial_start),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _4183_ (.RESET_B(net799),
    .D(net67),
    .Q(regFile_serial),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _4184_ (.RESET_B(net794),
    .D(_0162_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[0] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _4185_ (.RESET_B(net793),
    .D(_0163_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[1] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4186_ (.RESET_B(net793),
    .D(_0164_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[2] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _4187_ (.RESET_B(net794),
    .D(_0165_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[3] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _4188_ (.RESET_B(net794),
    .D(_0166_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[4] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _4189_ (.RESET_B(net800),
    .D(_0167_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[5] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _4190_ (.RESET_B(net797),
    .D(_0168_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[6] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _4191_ (.RESET_B(net800),
    .D(_0169_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[7] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _4192_ (.RESET_B(net796),
    .D(_0170_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][0] ),
    .CLK(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4193_ (.RESET_B(net787),
    .D(_0171_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][1] ),
    .CLK(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4194_ (.RESET_B(net773),
    .D(_0172_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][2] ),
    .CLK(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4195_ (.RESET_B(net793),
    .D(_0173_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][3] ),
    .CLK(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4196_ (.RESET_B(net781),
    .D(_0174_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][4] ),
    .CLK(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4197_ (.RESET_B(net779),
    .D(_0175_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][5] ),
    .CLK(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4198_ (.RESET_B(net780),
    .D(_0176_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][6] ),
    .CLK(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4199_ (.RESET_B(net775),
    .D(_0177_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.data[11][7] ),
    .CLK(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4200_ (.RESET_B(net785),
    .D(net35),
    .Q(clk_div_out),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _4201_ (.RESET_B(net788),
    .D(_0178_),
    .Q(\sap_3_inst.alu.act[0] ),
    .CLK(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4202_ (.RESET_B(net788),
    .D(_0179_),
    .Q(\sap_3_inst.alu.act[1] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4203_ (.RESET_B(net789),
    .D(_0180_),
    .Q(\sap_3_inst.alu.act[2] ),
    .CLK(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4204_ (.RESET_B(net789),
    .D(_0181_),
    .Q(\sap_3_inst.alu.act[3] ),
    .CLK(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4205_ (.RESET_B(net790),
    .D(_0182_),
    .Q(\sap_3_inst.alu.act[4] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4206_ (.RESET_B(net790),
    .D(_0183_),
    .Q(\sap_3_inst.alu.act[5] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_1 _4207_ (.RESET_B(net790),
    .D(_0184_),
    .Q(\sap_3_inst.alu.act[6] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4208_ (.RESET_B(net790),
    .D(_0185_),
    .Q(\sap_3_inst.alu.act[7] ),
    .CLK(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dfrbpq_2 _4209_ (.RESET_B(net783),
    .D(net766),
    .Q(\u_ser.state[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _4210_ (.RESET_B(net783),
    .D(_0187_),
    .Q(\u_ser.state[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _4211_ (.RESET_B(net783),
    .D(_0188_),
    .Q(sap_3_outputReg_serial),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _4212_ (.RESET_B(net783),
    .D(net69),
    .Q(sap_3_outputReg_start_sync),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _4213_ (.RESET_B(net797),
    .D(_0190_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _4214_ (.RESET_B(net797),
    .D(_0191_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _4215_ (.RESET_B(net797),
    .D(_0192_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _4216_ (.RESET_B(net797),
    .D(_0193_),
    .Q(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _4217_ (.RESET_B(net788),
    .D(_0194_),
    .Q(\u_ser.bit_pos[0] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _4218_ (.RESET_B(net784),
    .D(_0195_),
    .Q(\u_ser.bit_pos[1] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _4219_ (.RESET_B(net784),
    .D(net59),
    .Q(\u_ser.bit_pos[2] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_tielo heichips25_template_34 (.L_LO(net34));
 sg13g2_inv_1 _2076__1 (.Y(net35),
    .A(clknet_1_0__leaf_clk_div_out));
 sg13g2_buf_1 _4222_ (.A(mem_ram_we),
    .X(net25));
 sg13g2_buf_1 _4223_ (.A(mem_mar_we),
    .X(net26));
 sg13g2_buf_1 _4224_ (.A(sap_3_outputReg_serial),
    .X(net27));
 sg13g2_buf_1 _4225_ (.A(sap_3_outputReg_start_sync),
    .X(net28));
 sg13g2_buf_8 _4226_ (.A(regFile_serial),
    .X(net29));
 sg13g2_buf_8 _4227_ (.A(regFile_serial_start),
    .X(net30));
 sg13g2_lgcp_1 \sap_3_inst.clock.clock_gate_inst  (.GATE(_0001_),
    .CLK(clknet_1_1__leaf_clk_div_out),
    .GCLK(\sap_3_inst.alu.clk ));
 sg13g2_buf_8 fanout542 (.A(net542),
    .X(net24));
 sg13g2_buf_8 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_8 fanout544 (.A(_0331_),
    .X(net544));
 sg13g2_buf_8 fanout545 (.A(net545),
    .X(net19));
 sg13g2_buf_8 fanout546 (.A(_1975_),
    .X(net546));
 sg13g2_buf_8 fanout547 (.A(_1878_),
    .X(net547));
 sg13g2_buf_8 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_8 fanout549 (.A(_1394_),
    .X(net549));
 sg13g2_buf_8 fanout550 (.A(_1126_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_1126_),
    .X(net551));
 sg13g2_buf_8 fanout552 (.A(_0944_),
    .X(net552));
 sg13g2_buf_8 fanout553 (.A(_0751_),
    .X(net553));
 sg13g2_buf_8 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_8 fanout555 (.A(_0319_),
    .X(net555));
 sg13g2_buf_8 fanout556 (.A(_1210_),
    .X(net556));
 sg13g2_buf_8 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_8 fanout558 (.A(_1037_),
    .X(net558));
 sg13g2_buf_8 fanout559 (.A(net560),
    .X(net559));
 sg13g2_buf_8 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_8 fanout561 (.A(_0796_),
    .X(net561));
 sg13g2_buf_8 fanout562 (.A(_0716_),
    .X(net562));
 sg13g2_buf_8 fanout563 (.A(_0330_),
    .X(net563));
 sg13g2_buf_8 fanout564 (.A(_2007_),
    .X(net564));
 sg13g2_buf_8 fanout565 (.A(net567),
    .X(net565));
 sg13g2_buf_1 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_8 fanout567 (.A(_1673_),
    .X(net567));
 sg13g2_buf_8 fanout568 (.A(_1139_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_1139_),
    .X(net569));
 sg13g2_buf_8 fanout570 (.A(_1077_),
    .X(net570));
 sg13g2_buf_8 fanout571 (.A(_0837_),
    .X(net571));
 sg13g2_buf_8 fanout572 (.A(_0339_),
    .X(net572));
 sg13g2_buf_8 fanout573 (.A(_0338_),
    .X(net573));
 sg13g2_buf_8 fanout574 (.A(_0845_),
    .X(net574));
 sg13g2_buf_8 fanout575 (.A(_0843_),
    .X(net575));
 sg13g2_buf_8 fanout576 (.A(_0843_),
    .X(net576));
 sg13g2_buf_8 fanout577 (.A(net582),
    .X(net577));
 sg13g2_buf_8 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_8 fanout579 (.A(net582),
    .X(net579));
 sg13g2_buf_8 fanout580 (.A(net582),
    .X(net580));
 sg13g2_buf_1 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_8 fanout582 (.A(_0842_),
    .X(net582));
 sg13g2_buf_8 fanout583 (.A(_0830_),
    .X(net583));
 sg13g2_buf_8 fanout584 (.A(net586),
    .X(net584));
 sg13g2_buf_1 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_8 fanout586 (.A(_0829_),
    .X(net586));
 sg13g2_buf_8 fanout587 (.A(_0740_),
    .X(net587));
 sg13g2_buf_8 fanout588 (.A(_0740_),
    .X(net588));
 sg13g2_buf_8 fanout589 (.A(net591),
    .X(net589));
 sg13g2_buf_8 fanout590 (.A(net591),
    .X(net590));
 sg13g2_buf_8 fanout591 (.A(_0739_),
    .X(net591));
 sg13g2_buf_8 fanout592 (.A(_0738_),
    .X(net592));
 sg13g2_buf_1 fanout593 (.A(_0738_),
    .X(net593));
 sg13g2_buf_8 fanout594 (.A(_0734_),
    .X(net594));
 sg13g2_buf_8 fanout595 (.A(_0734_),
    .X(net595));
 sg13g2_buf_8 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_8 fanout597 (.A(_0727_),
    .X(net597));
 sg13g2_buf_8 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_8 fanout599 (.A(_0724_),
    .X(net599));
 sg13g2_buf_8 fanout600 (.A(_0724_),
    .X(net600));
 sg13g2_buf_1 fanout601 (.A(_0724_),
    .X(net601));
 sg13g2_buf_8 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_8 fanout603 (.A(_0722_),
    .X(net603));
 sg13g2_buf_8 fanout604 (.A(_0722_),
    .X(net604));
 sg13g2_buf_1 fanout605 (.A(_0722_),
    .X(net605));
 sg13g2_buf_8 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_8 fanout607 (.A(_0721_),
    .X(net607));
 sg13g2_buf_8 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_8 fanout609 (.A(_0721_),
    .X(net609));
 sg13g2_buf_8 fanout610 (.A(_0715_),
    .X(net610));
 sg13g2_buf_8 fanout611 (.A(_0715_),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(net613),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_8 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_8 fanout615 (.A(_0714_),
    .X(net615));
 sg13g2_buf_8 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_8 fanout617 (.A(_0310_),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(_1949_),
    .X(net618));
 sg13g2_buf_8 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_8 fanout620 (.A(_1803_),
    .X(net620));
 sg13g2_buf_8 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_8 fanout622 (.A(_1802_),
    .X(net622));
 sg13g2_buf_8 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_8 fanout624 (.A(_1801_),
    .X(net624));
 sg13g2_buf_8 fanout625 (.A(net626),
    .X(net625));
 sg13g2_buf_8 fanout626 (.A(_1800_),
    .X(net626));
 sg13g2_buf_8 fanout627 (.A(net628),
    .X(net627));
 sg13g2_buf_8 fanout628 (.A(_1799_),
    .X(net628));
 sg13g2_buf_8 fanout629 (.A(net630),
    .X(net629));
 sg13g2_buf_8 fanout630 (.A(_1798_),
    .X(net630));
 sg13g2_buf_8 fanout631 (.A(net632),
    .X(net631));
 sg13g2_buf_8 fanout632 (.A(_1797_),
    .X(net632));
 sg13g2_buf_8 fanout633 (.A(net634),
    .X(net633));
 sg13g2_buf_8 fanout634 (.A(_1796_),
    .X(net634));
 sg13g2_buf_8 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_8 fanout636 (.A(_1795_),
    .X(net636));
 sg13g2_buf_8 fanout637 (.A(_1794_),
    .X(net637));
 sg13g2_buf_8 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_8 fanout639 (.A(_1794_),
    .X(net639));
 sg13g2_buf_8 fanout640 (.A(net642),
    .X(net640));
 sg13g2_buf_8 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_8 fanout642 (.A(_0737_),
    .X(net642));
 sg13g2_buf_8 fanout643 (.A(net645),
    .X(net643));
 sg13g2_buf_1 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_8 fanout645 (.A(_0733_),
    .X(net645));
 sg13g2_buf_8 fanout646 (.A(net648),
    .X(net646));
 sg13g2_buf_1 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_8 fanout648 (.A(_0732_),
    .X(net648));
 sg13g2_buf_8 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_8 fanout650 (.A(_0729_),
    .X(net650));
 sg13g2_buf_8 fanout651 (.A(net652),
    .X(net651));
 sg13g2_buf_8 fanout652 (.A(net654),
    .X(net652));
 sg13g2_buf_8 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_8 fanout654 (.A(_0726_),
    .X(net654));
 sg13g2_buf_8 fanout655 (.A(net658),
    .X(net655));
 sg13g2_buf_8 fanout656 (.A(net658),
    .X(net656));
 sg13g2_buf_1 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_8 fanout658 (.A(_0723_),
    .X(net658));
 sg13g2_buf_8 fanout659 (.A(_0712_),
    .X(net659));
 sg13g2_buf_8 fanout660 (.A(_0625_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_0625_),
    .X(net661));
 sg13g2_buf_8 fanout662 (.A(_1746_),
    .X(net662));
 sg13g2_buf_8 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_8 fanout664 (.A(_1391_),
    .X(net664));
 sg13g2_buf_8 fanout665 (.A(_0671_),
    .X(net665));
 sg13g2_buf_8 fanout666 (.A(_0632_),
    .X(net666));
 sg13g2_buf_8 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_8 fanout668 (.A(_0585_),
    .X(net668));
 sg13g2_buf_8 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_8 fanout670 (.A(_0314_),
    .X(net670));
 sg13g2_buf_8 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_8 fanout672 (.A(_1947_),
    .X(net672));
 sg13g2_buf_8 fanout673 (.A(_0260_),
    .X(net673));
 sg13g2_buf_8 fanout674 (.A(_0260_),
    .X(net674));
 sg13g2_buf_8 fanout675 (.A(_1857_),
    .X(net675));
 sg13g2_buf_1 fanout676 (.A(_1857_),
    .X(net676));
 sg13g2_buf_8 fanout677 (.A(net679),
    .X(net677));
 sg13g2_buf_1 fanout678 (.A(net679),
    .X(net678));
 sg13g2_buf_8 fanout679 (.A(_1753_),
    .X(net679));
 sg13g2_buf_8 fanout680 (.A(net681),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_1617_),
    .X(net681));
 sg13g2_buf_8 fanout682 (.A(_1714_),
    .X(net682));
 sg13g2_buf_1 fanout683 (.A(_1714_),
    .X(net683));
 sg13g2_buf_8 fanout684 (.A(_1674_),
    .X(net684));
 sg13g2_buf_8 fanout685 (.A(_1674_),
    .X(net685));
 sg13g2_buf_8 fanout686 (.A(_1582_),
    .X(net686));
 sg13g2_buf_8 fanout687 (.A(net688),
    .X(net687));
 sg13g2_buf_8 fanout688 (.A(_1558_),
    .X(net688));
 sg13g2_buf_8 fanout689 (.A(_1552_),
    .X(net689));
 sg13g2_buf_1 fanout690 (.A(_1552_),
    .X(net690));
 sg13g2_buf_8 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_8 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_8 fanout693 (.A(_1532_),
    .X(net693));
 sg13g2_buf_8 fanout694 (.A(_1530_),
    .X(net694));
 sg13g2_buf_8 fanout695 (.A(_1530_),
    .X(net695));
 sg13g2_buf_8 fanout696 (.A(net701),
    .X(net696));
 sg13g2_buf_1 fanout697 (.A(net701),
    .X(net697));
 sg13g2_buf_8 fanout698 (.A(net701),
    .X(net698));
 sg13g2_buf_1 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_8 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_1529_),
    .X(net701));
 sg13g2_buf_8 fanout702 (.A(_1513_),
    .X(net702));
 sg13g2_buf_1 fanout703 (.A(_1513_),
    .X(net703));
 sg13g2_buf_8 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_8 fanout705 (.A(_1624_),
    .X(net705));
 sg13g2_buf_8 fanout706 (.A(_1611_),
    .X(net706));
 sg13g2_buf_8 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_8 fanout708 (.A(_1603_),
    .X(net708));
 sg13g2_buf_8 fanout709 (.A(_1565_),
    .X(net709));
 sg13g2_buf_8 fanout710 (.A(_1556_),
    .X(net710));
 sg13g2_buf_8 fanout711 (.A(_1531_),
    .X(net711));
 sg13g2_buf_8 fanout712 (.A(_1514_),
    .X(net712));
 sg13g2_buf_8 fanout713 (.A(_1512_),
    .X(net713));
 sg13g2_buf_8 fanout714 (.A(_1501_),
    .X(net714));
 sg13g2_buf_1 fanout715 (.A(_1501_),
    .X(net715));
 sg13g2_buf_8 fanout716 (.A(\sap_3_inst.controller.stage[3] ),
    .X(net716));
 sg13g2_buf_8 fanout717 (.A(\sap_3_inst.controller.stage[2] ),
    .X(net717));
 sg13g2_buf_8 fanout718 (.A(\sap_3_inst.controller.stage[1] ),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(\sap_3_inst.controller.stage[0] ),
    .X(net719));
 sg13g2_buf_8 fanout720 (.A(\sap_3_inst.alu.flags[1] ),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(_1314_),
    .X(net721));
 sg13g2_buf_8 fanout722 (.A(_1524_),
    .X(net722));
 sg13g2_buf_8 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_8 fanout724 (.A(_1505_),
    .X(net724));
 sg13g2_buf_8 fanout725 (.A(\sap_3_inst.controller.opcode[7] ),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(\sap_3_inst.controller.opcode[7] ),
    .X(net726));
 sg13g2_buf_8 fanout727 (.A(\sap_3_inst.controller.opcode[6] ),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(\sap_3_inst.controller.opcode[6] ),
    .X(net728));
 sg13g2_buf_8 fanout729 (.A(\sap_3_inst.controller.opcode[5] ),
    .X(net729));
 sg13g2_buf_8 fanout730 (.A(\sap_3_inst.controller.opcode[5] ),
    .X(net730));
 sg13g2_buf_8 fanout731 (.A(net732),
    .X(net731));
 sg13g2_buf_8 fanout732 (.A(\sap_3_inst.controller.opcode[4] ),
    .X(net732));
 sg13g2_buf_8 fanout733 (.A(net734),
    .X(net733));
 sg13g2_buf_8 fanout734 (.A(\sap_3_inst.controller.opcode[3] ),
    .X(net734));
 sg13g2_buf_8 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_8 fanout736 (.A(\sap_3_inst.controller.opcode[3] ),
    .X(net736));
 sg13g2_buf_8 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_8 fanout738 (.A(\sap_3_inst.controller.opcode[2] ),
    .X(net738));
 sg13g2_buf_8 fanout739 (.A(\sap_3_inst.controller.opcode[1] ),
    .X(net739));
 sg13g2_buf_8 fanout740 (.A(\sap_3_inst.controller.opcode[1] ),
    .X(net740));
 sg13g2_buf_8 fanout741 (.A(net742),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(\sap_3_inst.controller.opcode[0] ),
    .X(net742));
 sg13g2_buf_8 fanout743 (.A(net744),
    .X(net743));
 sg13g2_buf_8 fanout744 (.A(\sap_3_inst.alu.acc[7] ),
    .X(net744));
 sg13g2_buf_8 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_8 fanout746 (.A(\sap_3_inst.alu.acc[6] ),
    .X(net746));
 sg13g2_buf_8 fanout747 (.A(net749),
    .X(net747));
 sg13g2_buf_1 fanout748 (.A(net749),
    .X(net748));
 sg13g2_buf_8 fanout749 (.A(\sap_3_inst.alu.acc[5] ),
    .X(net749));
 sg13g2_buf_8 fanout750 (.A(net751),
    .X(net750));
 sg13g2_buf_8 fanout751 (.A(net752),
    .X(net751));
 sg13g2_buf_8 fanout752 (.A(\sap_3_inst.alu.acc[4] ),
    .X(net752));
 sg13g2_buf_8 fanout753 (.A(net754),
    .X(net753));
 sg13g2_buf_8 fanout754 (.A(\sap_3_inst.alu.acc[3] ),
    .X(net754));
 sg13g2_buf_8 fanout755 (.A(net756),
    .X(net755));
 sg13g2_buf_8 fanout756 (.A(\sap_3_inst.alu.acc[2] ),
    .X(net756));
 sg13g2_buf_8 fanout757 (.A(\sap_3_inst.alu.acc[1] ),
    .X(net757));
 sg13g2_buf_1 fanout758 (.A(\sap_3_inst.alu.acc[1] ),
    .X(net758));
 sg13g2_buf_8 fanout759 (.A(net760),
    .X(net759));
 sg13g2_buf_8 fanout760 (.A(\sap_3_inst.alu.acc[0] ),
    .X(net760));
 sg13g2_buf_8 fanout761 (.A(_1315_),
    .X(net761));
 sg13g2_buf_8 fanout762 (.A(net763),
    .X(net762));
 sg13g2_buf_8 fanout763 (.A(_1310_),
    .X(net763));
 sg13g2_buf_8 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_8 fanout765 (.A(_1280_),
    .X(net765));
 sg13g2_buf_8 fanout766 (.A(_0186_),
    .X(net766));
 sg13g2_buf_8 fanout767 (.A(\u_ser.bit_pos[0] ),
    .X(net767));
 sg13g2_buf_8 fanout768 (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[1] ),
    .X(net768));
 sg13g2_buf_8 fanout769 (.A(net80),
    .X(net769));
 sg13g2_buf_8 fanout770 (.A(net772),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_8 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_8 fanout773 (.A(net801),
    .X(net773));
 sg13g2_buf_8 fanout774 (.A(net778),
    .X(net774));
 sg13g2_buf_8 fanout775 (.A(net777),
    .X(net775));
 sg13g2_buf_8 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_8 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_8 fanout778 (.A(net801),
    .X(net778));
 sg13g2_buf_8 fanout779 (.A(net781),
    .X(net779));
 sg13g2_buf_8 fanout780 (.A(net781),
    .X(net780));
 sg13g2_buf_8 fanout781 (.A(net782),
    .X(net781));
 sg13g2_buf_8 fanout782 (.A(net801),
    .X(net782));
 sg13g2_buf_8 fanout783 (.A(net785),
    .X(net783));
 sg13g2_buf_8 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_8 fanout785 (.A(net792),
    .X(net785));
 sg13g2_buf_8 fanout786 (.A(net792),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(net792),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(net792),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(net792),
    .X(net789));
 sg13g2_buf_8 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_8 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(net801),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(net798),
    .X(net793));
 sg13g2_buf_1 fanout794 (.A(net798),
    .X(net794));
 sg13g2_buf_8 fanout795 (.A(net798),
    .X(net795));
 sg13g2_buf_8 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_8 fanout797 (.A(net798),
    .X(net797));
 sg13g2_buf_8 fanout798 (.A(net800),
    .X(net798));
 sg13g2_buf_8 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_8 fanout800 (.A(net801),
    .X(net800));
 sg13g2_buf_8 fanout801 (.A(rst_n),
    .X(net801));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[0]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[1]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[2]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[3]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[4]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[5]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[6]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[7]));
 sg13g2_buf_1 output17 (.A(net31),
    .X(uio_out[0]));
 sg13g2_buf_1 output18 (.A(net32),
    .X(uio_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[7]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[0]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[1]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[2]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[3]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[4]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[5]));
 sg13g2_buf_2 fanout31 (.A(net17),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(net18),
    .X(net32));
 sg13g2_tielo heichips25_template_33 (.L_LO(net33));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkbuf_0_clk_div_out (.A(clk_div_out),
    .X(clknet_0_clk_div_out));
 sg13g2_buf_8 clkbuf_1_0__f_clk_div_out (.A(clknet_0_clk_div_out),
    .X(clknet_1_0__leaf_clk_div_out));
 sg13g2_buf_8 clkbuf_1_1__f_clk_div_out (.A(clknet_0_clk_div_out),
    .X(clknet_1_1__leaf_clk_div_out));
 sg13g2_buf_1 clkload7 (.A(clknet_1_0__leaf_clk_div_out));
 sg13g2_buf_8 \clkbuf_leaf_0_sap_3_inst.alu.clk  (.A(\clknet_1_0__leaf_sap_3_inst.alu.clk ),
    .X(\clknet_leaf_0_sap_3_inst.alu.clk ));
 sg13g2_buf_8 \clkbuf_leaf_1_sap_3_inst.alu.clk  (.A(\clknet_1_1__leaf_sap_3_inst.alu.clk ),
    .X(\clknet_leaf_1_sap_3_inst.alu.clk ));
 sg13g2_buf_8 \clkbuf_leaf_2_sap_3_inst.alu.clk  (.A(\clknet_1_1__leaf_sap_3_inst.alu.clk ),
    .X(\clknet_leaf_2_sap_3_inst.alu.clk ));
 sg13g2_buf_8 \clkbuf_leaf_3_sap_3_inst.alu.clk  (.A(\clknet_1_0__leaf_sap_3_inst.alu.clk ),
    .X(\clknet_leaf_3_sap_3_inst.alu.clk ));
 sg13g2_buf_8 \clkbuf_0_sap_3_inst.alu.clk  (.A(\sap_3_inst.alu.clk ),
    .X(\clknet_0_sap_3_inst.alu.clk ));
 sg13g2_buf_8 \clkbuf_1_0__f_sap_3_inst.alu.clk  (.A(\clknet_0_sap_3_inst.alu.clk ),
    .X(\clknet_1_0__leaf_sap_3_inst.alu.clk ));
 sg13g2_buf_8 \clkbuf_1_1__f_sap_3_inst.alu.clk  (.A(\clknet_0_sap_3_inst.alu.clk ),
    .X(\clknet_1_1__leaf_sap_3_inst.alu.clk ));
 sg13g2_buf_8 \clkbuf_0_sap_3_inst.alu.clk_regs  (.A(\sap_3_inst.alu.clk_regs ),
    .X(\clknet_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_0_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_0_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_1_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_1_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_2_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_2_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_3_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_3_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_4_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_4_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_5_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_5_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_6_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_6_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_7_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_7_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_8_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_8_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_9_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_9_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_10_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_10_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_11_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_11_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_12_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_12_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_13_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_13_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_14_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_14_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_4_15_0_sap_3_inst.alu.clk_regs  (.A(\clknet_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_4_15_0_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_0__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_0_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_0__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_1__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_0_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_2__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_1_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_2__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_3__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_1_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_4__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_2_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_4__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_5__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_2_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_6__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_3_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_7__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_3_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_7__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_8__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_4_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_8__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_9__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_4_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_10__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_5_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_11__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_5_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_11__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_12__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_6_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_12__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_13__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_6_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_14__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_7_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_14__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_15__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_7_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_15__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_16__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_8_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_16__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_17__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_8_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_18__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_9_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_19__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_9_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_19__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_20__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_10_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_20__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_21__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_10_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_22__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_11_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_22__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_23__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_11_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_24__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_12_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_24__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_25__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_12_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_26__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_13_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_26__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_27__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_13_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_27__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_28__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_14_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_28__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_29__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_14_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_30__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_15_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_30__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_8 \clkbuf_5_31__f_sap_3_inst.alu.clk_regs  (.A(\clknet_4_15_0_sap_3_inst.alu.clk_regs ),
    .X(\clknet_5_31__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_inv_1 clkload8 (.A(\clknet_5_1__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_inv_1 clkload9 (.A(\clknet_5_3__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_inv_1 clkload10 (.A(\clknet_5_5__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_1 clkload11 (.A(\clknet_5_6__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_inv_1 clkload12 (.A(\clknet_5_9__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_1 clkload13 (.A(\clknet_5_10__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_inv_1 clkload14 (.A(\clknet_5_13__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_inv_1 clkload15 (.A(\clknet_5_17__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_1 clkload16 (.A(\clknet_5_18__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_inv_1 clkload17 (.A(\clknet_5_21__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_buf_1 clkload18 (.A(\clknet_5_23__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_inv_1 clkload19 (.A(\clknet_5_25__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_inv_1 clkload20 (.A(\clknet_5_29__leaf_sap_3_inst.alu.clk_regs ));
 sg13g2_dlygate4sd3_1 hold1 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[0] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold2 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[4] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold3 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[6] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold4 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[3] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold5 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[7] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold6 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[1] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold7 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[2] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold8 (.A(\sap_3_inst.reg_file.array_serializer_inst.shadow_reg[5] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_ser.shadow_reg[6] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_ser.shadow_reg[3] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_ser.state[0] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0196_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_ser.shadow_reg[7] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_ser.shadow_reg[1] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u_ser.shadow_reg[2] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold16 (.A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[2] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0159_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_ser.shadow_reg[5] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold19 (.A(regFile_serial),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0161_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold21 (.A(sap_3_outputReg_start_sync),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0189_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_ser.shadow_reg[0] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u_ser.bit_pos[1] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold25 (.A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[1] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0158_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_ser.shadow_reg[4] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold28 (.A(\sap_3_inst.reg_file.array_serializer_inst.state[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0160_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold30 (.A(sap_3_outputReg_serial),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold31 (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[3] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold32 (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[2] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold33 (.A(\sap_3_inst.reg_file.array_serializer_inst.bit_pos[0] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0157_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold35 (.A(\sap_3_inst.reg_file.array_serializer_inst.word_index[0] ),
    .X(net82));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_fill_2 FILLER_0_21 ();
 sg13g2_fill_1 FILLER_0_23 ();
 sg13g2_decap_8 FILLER_0_29 ();
 sg13g2_decap_8 FILLER_0_36 ();
 sg13g2_decap_8 FILLER_0_43 ();
 sg13g2_decap_8 FILLER_0_50 ();
 sg13g2_decap_8 FILLER_0_57 ();
 sg13g2_decap_8 FILLER_0_64 ();
 sg13g2_fill_2 FILLER_0_71 ();
 sg13g2_fill_1 FILLER_0_73 ();
 sg13g2_decap_8 FILLER_0_89 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_fill_2 FILLER_0_110 ();
 sg13g2_fill_1 FILLER_0_112 ();
 sg13g2_fill_1 FILLER_0_117 ();
 sg13g2_decap_4 FILLER_0_123 ();
 sg13g2_decap_8 FILLER_0_132 ();
 sg13g2_fill_1 FILLER_0_139 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_fill_2 FILLER_0_282 ();
 sg13g2_fill_2 FILLER_0_311 ();
 sg13g2_fill_1 FILLER_0_338 ();
 sg13g2_fill_1 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_435 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_decap_8 FILLER_0_449 ();
 sg13g2_decap_8 FILLER_0_456 ();
 sg13g2_decap_8 FILLER_0_463 ();
 sg13g2_decap_8 FILLER_0_470 ();
 sg13g2_decap_8 FILLER_0_477 ();
 sg13g2_decap_8 FILLER_0_484 ();
 sg13g2_decap_8 FILLER_0_491 ();
 sg13g2_decap_8 FILLER_0_498 ();
 sg13g2_decap_8 FILLER_0_505 ();
 sg13g2_decap_8 FILLER_0_512 ();
 sg13g2_decap_8 FILLER_0_519 ();
 sg13g2_decap_8 FILLER_0_526 ();
 sg13g2_decap_8 FILLER_0_533 ();
 sg13g2_decap_8 FILLER_0_540 ();
 sg13g2_decap_8 FILLER_0_547 ();
 sg13g2_decap_8 FILLER_0_554 ();
 sg13g2_decap_8 FILLER_0_561 ();
 sg13g2_decap_8 FILLER_0_568 ();
 sg13g2_decap_8 FILLER_0_575 ();
 sg13g2_decap_8 FILLER_0_582 ();
 sg13g2_decap_8 FILLER_0_589 ();
 sg13g2_decap_8 FILLER_0_596 ();
 sg13g2_decap_8 FILLER_0_603 ();
 sg13g2_decap_8 FILLER_0_610 ();
 sg13g2_decap_8 FILLER_0_617 ();
 sg13g2_decap_8 FILLER_0_624 ();
 sg13g2_decap_8 FILLER_0_631 ();
 sg13g2_decap_8 FILLER_0_638 ();
 sg13g2_decap_8 FILLER_0_645 ();
 sg13g2_decap_8 FILLER_0_652 ();
 sg13g2_decap_8 FILLER_0_659 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_8 FILLER_0_673 ();
 sg13g2_decap_8 FILLER_0_680 ();
 sg13g2_decap_8 FILLER_0_687 ();
 sg13g2_decap_8 FILLER_0_694 ();
 sg13g2_decap_8 FILLER_0_701 ();
 sg13g2_decap_8 FILLER_0_708 ();
 sg13g2_decap_8 FILLER_0_715 ();
 sg13g2_decap_8 FILLER_0_722 ();
 sg13g2_decap_8 FILLER_0_729 ();
 sg13g2_decap_8 FILLER_0_736 ();
 sg13g2_decap_8 FILLER_0_743 ();
 sg13g2_decap_8 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_757 ();
 sg13g2_decap_8 FILLER_0_764 ();
 sg13g2_decap_8 FILLER_0_771 ();
 sg13g2_decap_8 FILLER_0_778 ();
 sg13g2_decap_8 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_decap_8 FILLER_0_799 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_8 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_820 ();
 sg13g2_decap_8 FILLER_0_827 ();
 sg13g2_decap_8 FILLER_0_834 ();
 sg13g2_decap_8 FILLER_0_841 ();
 sg13g2_decap_8 FILLER_0_848 ();
 sg13g2_decap_8 FILLER_0_855 ();
 sg13g2_decap_8 FILLER_0_862 ();
 sg13g2_decap_8 FILLER_0_869 ();
 sg13g2_decap_8 FILLER_0_876 ();
 sg13g2_decap_8 FILLER_0_883 ();
 sg13g2_decap_8 FILLER_0_890 ();
 sg13g2_decap_8 FILLER_0_897 ();
 sg13g2_decap_8 FILLER_0_904 ();
 sg13g2_decap_8 FILLER_0_911 ();
 sg13g2_decap_8 FILLER_0_918 ();
 sg13g2_decap_8 FILLER_0_925 ();
 sg13g2_decap_8 FILLER_0_932 ();
 sg13g2_decap_8 FILLER_0_939 ();
 sg13g2_decap_8 FILLER_0_946 ();
 sg13g2_decap_8 FILLER_0_953 ();
 sg13g2_decap_8 FILLER_0_960 ();
 sg13g2_decap_8 FILLER_0_967 ();
 sg13g2_decap_8 FILLER_0_974 ();
 sg13g2_decap_8 FILLER_0_981 ();
 sg13g2_decap_8 FILLER_0_988 ();
 sg13g2_decap_8 FILLER_0_995 ();
 sg13g2_decap_8 FILLER_0_1002 ();
 sg13g2_decap_8 FILLER_0_1009 ();
 sg13g2_decap_8 FILLER_0_1016 ();
 sg13g2_decap_4 FILLER_0_1023 ();
 sg13g2_fill_2 FILLER_0_1027 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_7 ();
 sg13g2_fill_1 FILLER_1_9 ();
 sg13g2_fill_2 FILLER_1_33 ();
 sg13g2_decap_4 FILLER_1_39 ();
 sg13g2_fill_1 FILLER_1_43 ();
 sg13g2_decap_4 FILLER_1_54 ();
 sg13g2_fill_1 FILLER_1_66 ();
 sg13g2_fill_2 FILLER_1_78 ();
 sg13g2_decap_4 FILLER_1_93 ();
 sg13g2_fill_2 FILLER_1_107 ();
 sg13g2_fill_1 FILLER_1_109 ();
 sg13g2_decap_4 FILLER_1_134 ();
 sg13g2_decap_8 FILLER_1_155 ();
 sg13g2_fill_2 FILLER_1_185 ();
 sg13g2_fill_2 FILLER_1_214 ();
 sg13g2_fill_2 FILLER_1_258 ();
 sg13g2_fill_1 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_443 ();
 sg13g2_decap_8 FILLER_1_450 ();
 sg13g2_decap_8 FILLER_1_457 ();
 sg13g2_decap_8 FILLER_1_464 ();
 sg13g2_decap_8 FILLER_1_471 ();
 sg13g2_decap_8 FILLER_1_478 ();
 sg13g2_decap_8 FILLER_1_485 ();
 sg13g2_decap_8 FILLER_1_492 ();
 sg13g2_decap_8 FILLER_1_499 ();
 sg13g2_decap_8 FILLER_1_506 ();
 sg13g2_decap_8 FILLER_1_513 ();
 sg13g2_decap_8 FILLER_1_520 ();
 sg13g2_decap_8 FILLER_1_527 ();
 sg13g2_decap_8 FILLER_1_534 ();
 sg13g2_decap_8 FILLER_1_541 ();
 sg13g2_decap_8 FILLER_1_548 ();
 sg13g2_decap_8 FILLER_1_555 ();
 sg13g2_decap_8 FILLER_1_562 ();
 sg13g2_decap_8 FILLER_1_569 ();
 sg13g2_decap_8 FILLER_1_576 ();
 sg13g2_decap_8 FILLER_1_583 ();
 sg13g2_decap_8 FILLER_1_590 ();
 sg13g2_decap_8 FILLER_1_597 ();
 sg13g2_decap_8 FILLER_1_604 ();
 sg13g2_decap_8 FILLER_1_611 ();
 sg13g2_decap_8 FILLER_1_618 ();
 sg13g2_decap_8 FILLER_1_625 ();
 sg13g2_decap_8 FILLER_1_632 ();
 sg13g2_decap_8 FILLER_1_639 ();
 sg13g2_decap_8 FILLER_1_646 ();
 sg13g2_decap_8 FILLER_1_653 ();
 sg13g2_decap_8 FILLER_1_660 ();
 sg13g2_decap_8 FILLER_1_667 ();
 sg13g2_decap_8 FILLER_1_674 ();
 sg13g2_decap_8 FILLER_1_681 ();
 sg13g2_decap_8 FILLER_1_688 ();
 sg13g2_decap_8 FILLER_1_695 ();
 sg13g2_decap_8 FILLER_1_702 ();
 sg13g2_decap_8 FILLER_1_709 ();
 sg13g2_decap_8 FILLER_1_716 ();
 sg13g2_decap_8 FILLER_1_723 ();
 sg13g2_decap_8 FILLER_1_730 ();
 sg13g2_decap_8 FILLER_1_737 ();
 sg13g2_decap_8 FILLER_1_744 ();
 sg13g2_decap_8 FILLER_1_751 ();
 sg13g2_decap_8 FILLER_1_758 ();
 sg13g2_decap_8 FILLER_1_765 ();
 sg13g2_decap_8 FILLER_1_772 ();
 sg13g2_decap_8 FILLER_1_779 ();
 sg13g2_decap_8 FILLER_1_786 ();
 sg13g2_decap_8 FILLER_1_793 ();
 sg13g2_decap_8 FILLER_1_800 ();
 sg13g2_decap_8 FILLER_1_807 ();
 sg13g2_decap_8 FILLER_1_814 ();
 sg13g2_decap_8 FILLER_1_821 ();
 sg13g2_decap_8 FILLER_1_828 ();
 sg13g2_decap_8 FILLER_1_835 ();
 sg13g2_decap_8 FILLER_1_842 ();
 sg13g2_decap_8 FILLER_1_849 ();
 sg13g2_decap_8 FILLER_1_856 ();
 sg13g2_decap_8 FILLER_1_863 ();
 sg13g2_decap_8 FILLER_1_870 ();
 sg13g2_decap_8 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_1_884 ();
 sg13g2_decap_8 FILLER_1_891 ();
 sg13g2_decap_8 FILLER_1_898 ();
 sg13g2_decap_8 FILLER_1_905 ();
 sg13g2_decap_8 FILLER_1_912 ();
 sg13g2_decap_8 FILLER_1_919 ();
 sg13g2_decap_8 FILLER_1_926 ();
 sg13g2_decap_8 FILLER_1_933 ();
 sg13g2_decap_8 FILLER_1_940 ();
 sg13g2_decap_8 FILLER_1_947 ();
 sg13g2_decap_8 FILLER_1_954 ();
 sg13g2_decap_8 FILLER_1_961 ();
 sg13g2_decap_8 FILLER_1_968 ();
 sg13g2_decap_8 FILLER_1_975 ();
 sg13g2_decap_8 FILLER_1_982 ();
 sg13g2_decap_8 FILLER_1_989 ();
 sg13g2_decap_8 FILLER_1_996 ();
 sg13g2_decap_8 FILLER_1_1003 ();
 sg13g2_decap_8 FILLER_1_1010 ();
 sg13g2_decap_8 FILLER_1_1017 ();
 sg13g2_decap_4 FILLER_1_1024 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_fill_1 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_30 ();
 sg13g2_fill_1 FILLER_2_37 ();
 sg13g2_fill_1 FILLER_2_80 ();
 sg13g2_fill_1 FILLER_2_91 ();
 sg13g2_fill_2 FILLER_2_96 ();
 sg13g2_decap_4 FILLER_2_122 ();
 sg13g2_decap_4 FILLER_2_131 ();
 sg13g2_fill_1 FILLER_2_135 ();
 sg13g2_fill_2 FILLER_2_141 ();
 sg13g2_fill_1 FILLER_2_143 ();
 sg13g2_decap_4 FILLER_2_147 ();
 sg13g2_fill_1 FILLER_2_172 ();
 sg13g2_fill_1 FILLER_2_208 ();
 sg13g2_fill_1 FILLER_2_256 ();
 sg13g2_fill_1 FILLER_2_284 ();
 sg13g2_fill_1 FILLER_2_360 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_decap_8 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_882 ();
 sg13g2_decap_8 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_decap_8 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_924 ();
 sg13g2_decap_8 FILLER_2_931 ();
 sg13g2_decap_8 FILLER_2_938 ();
 sg13g2_decap_8 FILLER_2_945 ();
 sg13g2_decap_8 FILLER_2_952 ();
 sg13g2_decap_8 FILLER_2_959 ();
 sg13g2_decap_8 FILLER_2_966 ();
 sg13g2_decap_8 FILLER_2_973 ();
 sg13g2_decap_8 FILLER_2_980 ();
 sg13g2_decap_8 FILLER_2_987 ();
 sg13g2_decap_8 FILLER_2_994 ();
 sg13g2_decap_8 FILLER_2_1001 ();
 sg13g2_decap_8 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1015 ();
 sg13g2_decap_8 FILLER_2_1022 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_fill_2 FILLER_3_11 ();
 sg13g2_fill_1 FILLER_3_13 ();
 sg13g2_decap_8 FILLER_3_23 ();
 sg13g2_fill_2 FILLER_3_30 ();
 sg13g2_fill_2 FILLER_3_58 ();
 sg13g2_decap_8 FILLER_3_64 ();
 sg13g2_decap_4 FILLER_3_71 ();
 sg13g2_fill_1 FILLER_3_75 ();
 sg13g2_decap_8 FILLER_3_92 ();
 sg13g2_decap_4 FILLER_3_99 ();
 sg13g2_fill_1 FILLER_3_103 ();
 sg13g2_fill_1 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_115 ();
 sg13g2_decap_8 FILLER_3_122 ();
 sg13g2_decap_8 FILLER_3_129 ();
 sg13g2_decap_8 FILLER_3_136 ();
 sg13g2_decap_4 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_152 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_fill_1 FILLER_3_211 ();
 sg13g2_fill_2 FILLER_3_362 ();
 sg13g2_fill_1 FILLER_3_364 ();
 sg13g2_fill_1 FILLER_3_380 ();
 sg13g2_fill_2 FILLER_3_400 ();
 sg13g2_fill_1 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_3_444 ();
 sg13g2_decap_8 FILLER_3_451 ();
 sg13g2_decap_8 FILLER_3_458 ();
 sg13g2_decap_8 FILLER_3_465 ();
 sg13g2_decap_8 FILLER_3_472 ();
 sg13g2_decap_8 FILLER_3_479 ();
 sg13g2_decap_8 FILLER_3_486 ();
 sg13g2_decap_8 FILLER_3_493 ();
 sg13g2_decap_8 FILLER_3_500 ();
 sg13g2_decap_8 FILLER_3_507 ();
 sg13g2_decap_8 FILLER_3_514 ();
 sg13g2_decap_8 FILLER_3_521 ();
 sg13g2_decap_8 FILLER_3_528 ();
 sg13g2_decap_8 FILLER_3_535 ();
 sg13g2_decap_8 FILLER_3_542 ();
 sg13g2_decap_8 FILLER_3_549 ();
 sg13g2_decap_8 FILLER_3_556 ();
 sg13g2_decap_8 FILLER_3_563 ();
 sg13g2_decap_8 FILLER_3_570 ();
 sg13g2_decap_8 FILLER_3_577 ();
 sg13g2_decap_8 FILLER_3_584 ();
 sg13g2_decap_8 FILLER_3_591 ();
 sg13g2_decap_8 FILLER_3_598 ();
 sg13g2_decap_8 FILLER_3_605 ();
 sg13g2_decap_8 FILLER_3_612 ();
 sg13g2_decap_8 FILLER_3_619 ();
 sg13g2_decap_8 FILLER_3_626 ();
 sg13g2_decap_8 FILLER_3_633 ();
 sg13g2_decap_8 FILLER_3_640 ();
 sg13g2_decap_8 FILLER_3_647 ();
 sg13g2_decap_8 FILLER_3_654 ();
 sg13g2_decap_8 FILLER_3_661 ();
 sg13g2_decap_8 FILLER_3_668 ();
 sg13g2_decap_8 FILLER_3_675 ();
 sg13g2_decap_8 FILLER_3_682 ();
 sg13g2_decap_8 FILLER_3_689 ();
 sg13g2_decap_8 FILLER_3_696 ();
 sg13g2_decap_8 FILLER_3_703 ();
 sg13g2_decap_8 FILLER_3_710 ();
 sg13g2_decap_8 FILLER_3_717 ();
 sg13g2_decap_8 FILLER_3_724 ();
 sg13g2_decap_8 FILLER_3_731 ();
 sg13g2_decap_8 FILLER_3_738 ();
 sg13g2_decap_8 FILLER_3_745 ();
 sg13g2_decap_8 FILLER_3_752 ();
 sg13g2_decap_8 FILLER_3_759 ();
 sg13g2_decap_8 FILLER_3_766 ();
 sg13g2_decap_8 FILLER_3_773 ();
 sg13g2_decap_8 FILLER_3_780 ();
 sg13g2_decap_8 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_794 ();
 sg13g2_decap_8 FILLER_3_801 ();
 sg13g2_decap_8 FILLER_3_808 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_decap_8 FILLER_3_829 ();
 sg13g2_decap_8 FILLER_3_836 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_850 ();
 sg13g2_decap_8 FILLER_3_857 ();
 sg13g2_decap_8 FILLER_3_864 ();
 sg13g2_decap_8 FILLER_3_871 ();
 sg13g2_decap_8 FILLER_3_878 ();
 sg13g2_decap_8 FILLER_3_885 ();
 sg13g2_decap_8 FILLER_3_892 ();
 sg13g2_decap_8 FILLER_3_899 ();
 sg13g2_decap_8 FILLER_3_906 ();
 sg13g2_decap_8 FILLER_3_913 ();
 sg13g2_decap_8 FILLER_3_920 ();
 sg13g2_decap_8 FILLER_3_927 ();
 sg13g2_decap_8 FILLER_3_934 ();
 sg13g2_decap_8 FILLER_3_941 ();
 sg13g2_decap_8 FILLER_3_948 ();
 sg13g2_decap_8 FILLER_3_955 ();
 sg13g2_decap_8 FILLER_3_962 ();
 sg13g2_decap_8 FILLER_3_969 ();
 sg13g2_decap_8 FILLER_3_976 ();
 sg13g2_decap_8 FILLER_3_983 ();
 sg13g2_decap_8 FILLER_3_990 ();
 sg13g2_decap_8 FILLER_3_997 ();
 sg13g2_decap_8 FILLER_3_1004 ();
 sg13g2_decap_8 FILLER_3_1011 ();
 sg13g2_decap_8 FILLER_3_1018 ();
 sg13g2_decap_4 FILLER_3_1025 ();
 sg13g2_fill_1 FILLER_4_34 ();
 sg13g2_decap_8 FILLER_4_55 ();
 sg13g2_fill_1 FILLER_4_62 ();
 sg13g2_fill_1 FILLER_4_67 ();
 sg13g2_fill_2 FILLER_4_72 ();
 sg13g2_fill_2 FILLER_4_79 ();
 sg13g2_fill_1 FILLER_4_81 ();
 sg13g2_decap_8 FILLER_4_87 ();
 sg13g2_fill_1 FILLER_4_94 ();
 sg13g2_decap_4 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_121 ();
 sg13g2_fill_2 FILLER_4_147 ();
 sg13g2_fill_2 FILLER_4_167 ();
 sg13g2_fill_1 FILLER_4_210 ();
 sg13g2_fill_1 FILLER_4_337 ();
 sg13g2_fill_1 FILLER_4_402 ();
 sg13g2_fill_2 FILLER_4_447 ();
 sg13g2_fill_1 FILLER_4_449 ();
 sg13g2_decap_8 FILLER_4_453 ();
 sg13g2_decap_8 FILLER_4_460 ();
 sg13g2_decap_8 FILLER_4_467 ();
 sg13g2_decap_8 FILLER_4_474 ();
 sg13g2_decap_8 FILLER_4_481 ();
 sg13g2_decap_8 FILLER_4_488 ();
 sg13g2_decap_8 FILLER_4_495 ();
 sg13g2_decap_8 FILLER_4_502 ();
 sg13g2_decap_8 FILLER_4_509 ();
 sg13g2_decap_8 FILLER_4_516 ();
 sg13g2_decap_8 FILLER_4_523 ();
 sg13g2_decap_8 FILLER_4_530 ();
 sg13g2_decap_8 FILLER_4_537 ();
 sg13g2_decap_8 FILLER_4_544 ();
 sg13g2_decap_8 FILLER_4_551 ();
 sg13g2_decap_8 FILLER_4_558 ();
 sg13g2_decap_8 FILLER_4_565 ();
 sg13g2_decap_8 FILLER_4_572 ();
 sg13g2_decap_8 FILLER_4_579 ();
 sg13g2_decap_8 FILLER_4_586 ();
 sg13g2_decap_8 FILLER_4_593 ();
 sg13g2_decap_8 FILLER_4_600 ();
 sg13g2_decap_8 FILLER_4_607 ();
 sg13g2_decap_8 FILLER_4_614 ();
 sg13g2_decap_8 FILLER_4_621 ();
 sg13g2_decap_8 FILLER_4_628 ();
 sg13g2_decap_8 FILLER_4_635 ();
 sg13g2_decap_8 FILLER_4_642 ();
 sg13g2_decap_8 FILLER_4_649 ();
 sg13g2_decap_8 FILLER_4_656 ();
 sg13g2_decap_8 FILLER_4_663 ();
 sg13g2_decap_8 FILLER_4_670 ();
 sg13g2_decap_8 FILLER_4_677 ();
 sg13g2_decap_8 FILLER_4_684 ();
 sg13g2_decap_8 FILLER_4_691 ();
 sg13g2_decap_8 FILLER_4_698 ();
 sg13g2_decap_8 FILLER_4_705 ();
 sg13g2_decap_8 FILLER_4_712 ();
 sg13g2_decap_8 FILLER_4_719 ();
 sg13g2_decap_8 FILLER_4_726 ();
 sg13g2_decap_8 FILLER_4_733 ();
 sg13g2_decap_8 FILLER_4_740 ();
 sg13g2_decap_8 FILLER_4_747 ();
 sg13g2_decap_8 FILLER_4_754 ();
 sg13g2_decap_8 FILLER_4_761 ();
 sg13g2_decap_8 FILLER_4_768 ();
 sg13g2_decap_8 FILLER_4_775 ();
 sg13g2_decap_8 FILLER_4_782 ();
 sg13g2_decap_8 FILLER_4_789 ();
 sg13g2_decap_8 FILLER_4_796 ();
 sg13g2_decap_8 FILLER_4_803 ();
 sg13g2_decap_8 FILLER_4_810 ();
 sg13g2_decap_8 FILLER_4_817 ();
 sg13g2_decap_8 FILLER_4_824 ();
 sg13g2_decap_8 FILLER_4_831 ();
 sg13g2_decap_8 FILLER_4_838 ();
 sg13g2_decap_8 FILLER_4_845 ();
 sg13g2_decap_8 FILLER_4_852 ();
 sg13g2_decap_8 FILLER_4_859 ();
 sg13g2_decap_8 FILLER_4_866 ();
 sg13g2_decap_8 FILLER_4_873 ();
 sg13g2_decap_8 FILLER_4_880 ();
 sg13g2_decap_8 FILLER_4_887 ();
 sg13g2_decap_8 FILLER_4_894 ();
 sg13g2_decap_8 FILLER_4_901 ();
 sg13g2_decap_8 FILLER_4_908 ();
 sg13g2_decap_8 FILLER_4_915 ();
 sg13g2_decap_8 FILLER_4_922 ();
 sg13g2_decap_8 FILLER_4_929 ();
 sg13g2_decap_8 FILLER_4_936 ();
 sg13g2_decap_8 FILLER_4_943 ();
 sg13g2_decap_8 FILLER_4_950 ();
 sg13g2_decap_8 FILLER_4_957 ();
 sg13g2_decap_8 FILLER_4_964 ();
 sg13g2_decap_8 FILLER_4_971 ();
 sg13g2_decap_8 FILLER_4_978 ();
 sg13g2_decap_8 FILLER_4_985 ();
 sg13g2_decap_8 FILLER_4_992 ();
 sg13g2_decap_8 FILLER_4_999 ();
 sg13g2_decap_8 FILLER_4_1006 ();
 sg13g2_decap_8 FILLER_4_1013 ();
 sg13g2_decap_8 FILLER_4_1020 ();
 sg13g2_fill_2 FILLER_4_1027 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_4 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_20 ();
 sg13g2_decap_8 FILLER_5_27 ();
 sg13g2_fill_2 FILLER_5_34 ();
 sg13g2_fill_1 FILLER_5_36 ();
 sg13g2_fill_2 FILLER_5_62 ();
 sg13g2_fill_1 FILLER_5_69 ();
 sg13g2_decap_4 FILLER_5_83 ();
 sg13g2_fill_1 FILLER_5_87 ();
 sg13g2_fill_2 FILLER_5_93 ();
 sg13g2_decap_4 FILLER_5_109 ();
 sg13g2_fill_2 FILLER_5_113 ();
 sg13g2_fill_1 FILLER_5_126 ();
 sg13g2_fill_2 FILLER_5_140 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_fill_2 FILLER_5_149 ();
 sg13g2_fill_2 FILLER_5_157 ();
 sg13g2_fill_1 FILLER_5_159 ();
 sg13g2_fill_1 FILLER_5_168 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_fill_1 FILLER_5_213 ();
 sg13g2_fill_2 FILLER_5_311 ();
 sg13g2_fill_2 FILLER_5_438 ();
 sg13g2_decap_8 FILLER_5_460 ();
 sg13g2_decap_8 FILLER_5_467 ();
 sg13g2_decap_8 FILLER_5_474 ();
 sg13g2_decap_8 FILLER_5_481 ();
 sg13g2_decap_8 FILLER_5_488 ();
 sg13g2_decap_8 FILLER_5_495 ();
 sg13g2_decap_8 FILLER_5_502 ();
 sg13g2_decap_8 FILLER_5_509 ();
 sg13g2_decap_8 FILLER_5_516 ();
 sg13g2_decap_8 FILLER_5_523 ();
 sg13g2_decap_8 FILLER_5_530 ();
 sg13g2_decap_8 FILLER_5_537 ();
 sg13g2_decap_8 FILLER_5_544 ();
 sg13g2_decap_8 FILLER_5_551 ();
 sg13g2_decap_8 FILLER_5_558 ();
 sg13g2_decap_8 FILLER_5_565 ();
 sg13g2_decap_8 FILLER_5_572 ();
 sg13g2_decap_8 FILLER_5_579 ();
 sg13g2_decap_8 FILLER_5_586 ();
 sg13g2_decap_8 FILLER_5_593 ();
 sg13g2_decap_8 FILLER_5_600 ();
 sg13g2_decap_8 FILLER_5_607 ();
 sg13g2_decap_8 FILLER_5_614 ();
 sg13g2_decap_8 FILLER_5_621 ();
 sg13g2_decap_8 FILLER_5_628 ();
 sg13g2_decap_8 FILLER_5_635 ();
 sg13g2_decap_8 FILLER_5_642 ();
 sg13g2_decap_8 FILLER_5_649 ();
 sg13g2_decap_8 FILLER_5_656 ();
 sg13g2_decap_8 FILLER_5_663 ();
 sg13g2_decap_8 FILLER_5_670 ();
 sg13g2_decap_8 FILLER_5_677 ();
 sg13g2_decap_8 FILLER_5_684 ();
 sg13g2_decap_8 FILLER_5_691 ();
 sg13g2_decap_8 FILLER_5_698 ();
 sg13g2_decap_8 FILLER_5_705 ();
 sg13g2_decap_8 FILLER_5_712 ();
 sg13g2_decap_8 FILLER_5_719 ();
 sg13g2_decap_8 FILLER_5_726 ();
 sg13g2_decap_8 FILLER_5_733 ();
 sg13g2_decap_8 FILLER_5_740 ();
 sg13g2_decap_8 FILLER_5_747 ();
 sg13g2_decap_8 FILLER_5_754 ();
 sg13g2_decap_8 FILLER_5_761 ();
 sg13g2_decap_8 FILLER_5_768 ();
 sg13g2_decap_8 FILLER_5_775 ();
 sg13g2_decap_8 FILLER_5_782 ();
 sg13g2_decap_8 FILLER_5_789 ();
 sg13g2_decap_8 FILLER_5_796 ();
 sg13g2_decap_8 FILLER_5_803 ();
 sg13g2_decap_8 FILLER_5_810 ();
 sg13g2_decap_8 FILLER_5_817 ();
 sg13g2_decap_8 FILLER_5_824 ();
 sg13g2_decap_8 FILLER_5_831 ();
 sg13g2_decap_8 FILLER_5_838 ();
 sg13g2_decap_8 FILLER_5_845 ();
 sg13g2_decap_8 FILLER_5_852 ();
 sg13g2_decap_8 FILLER_5_859 ();
 sg13g2_decap_8 FILLER_5_866 ();
 sg13g2_decap_8 FILLER_5_873 ();
 sg13g2_decap_8 FILLER_5_880 ();
 sg13g2_decap_8 FILLER_5_887 ();
 sg13g2_decap_8 FILLER_5_894 ();
 sg13g2_decap_8 FILLER_5_901 ();
 sg13g2_decap_8 FILLER_5_908 ();
 sg13g2_decap_8 FILLER_5_915 ();
 sg13g2_decap_8 FILLER_5_922 ();
 sg13g2_decap_8 FILLER_5_929 ();
 sg13g2_decap_8 FILLER_5_936 ();
 sg13g2_decap_8 FILLER_5_943 ();
 sg13g2_decap_8 FILLER_5_950 ();
 sg13g2_decap_8 FILLER_5_957 ();
 sg13g2_decap_8 FILLER_5_964 ();
 sg13g2_decap_8 FILLER_5_971 ();
 sg13g2_decap_8 FILLER_5_978 ();
 sg13g2_decap_8 FILLER_5_985 ();
 sg13g2_decap_8 FILLER_5_992 ();
 sg13g2_decap_8 FILLER_5_999 ();
 sg13g2_decap_8 FILLER_5_1006 ();
 sg13g2_decap_8 FILLER_5_1013 ();
 sg13g2_decap_8 FILLER_5_1020 ();
 sg13g2_fill_2 FILLER_5_1027 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_fill_2 FILLER_6_27 ();
 sg13g2_fill_1 FILLER_6_29 ();
 sg13g2_decap_4 FILLER_6_36 ();
 sg13g2_fill_2 FILLER_6_57 ();
 sg13g2_decap_8 FILLER_6_83 ();
 sg13g2_fill_2 FILLER_6_90 ();
 sg13g2_fill_1 FILLER_6_92 ();
 sg13g2_fill_2 FILLER_6_132 ();
 sg13g2_fill_1 FILLER_6_142 ();
 sg13g2_fill_1 FILLER_6_182 ();
 sg13g2_fill_2 FILLER_6_198 ();
 sg13g2_fill_2 FILLER_6_301 ();
 sg13g2_fill_1 FILLER_6_349 ();
 sg13g2_fill_2 FILLER_6_381 ();
 sg13g2_fill_1 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_484 ();
 sg13g2_decap_8 FILLER_6_491 ();
 sg13g2_decap_8 FILLER_6_498 ();
 sg13g2_decap_8 FILLER_6_505 ();
 sg13g2_decap_8 FILLER_6_512 ();
 sg13g2_decap_8 FILLER_6_519 ();
 sg13g2_decap_8 FILLER_6_526 ();
 sg13g2_decap_8 FILLER_6_533 ();
 sg13g2_decap_8 FILLER_6_540 ();
 sg13g2_decap_8 FILLER_6_547 ();
 sg13g2_decap_8 FILLER_6_554 ();
 sg13g2_decap_8 FILLER_6_561 ();
 sg13g2_decap_8 FILLER_6_568 ();
 sg13g2_decap_8 FILLER_6_575 ();
 sg13g2_decap_8 FILLER_6_582 ();
 sg13g2_decap_8 FILLER_6_589 ();
 sg13g2_decap_8 FILLER_6_596 ();
 sg13g2_decap_8 FILLER_6_603 ();
 sg13g2_decap_8 FILLER_6_610 ();
 sg13g2_decap_8 FILLER_6_617 ();
 sg13g2_decap_8 FILLER_6_624 ();
 sg13g2_decap_8 FILLER_6_631 ();
 sg13g2_decap_8 FILLER_6_638 ();
 sg13g2_decap_8 FILLER_6_645 ();
 sg13g2_decap_8 FILLER_6_652 ();
 sg13g2_decap_8 FILLER_6_659 ();
 sg13g2_decap_8 FILLER_6_666 ();
 sg13g2_decap_8 FILLER_6_673 ();
 sg13g2_decap_8 FILLER_6_680 ();
 sg13g2_decap_8 FILLER_6_687 ();
 sg13g2_decap_8 FILLER_6_694 ();
 sg13g2_decap_8 FILLER_6_701 ();
 sg13g2_decap_8 FILLER_6_708 ();
 sg13g2_decap_8 FILLER_6_715 ();
 sg13g2_decap_8 FILLER_6_722 ();
 sg13g2_decap_8 FILLER_6_729 ();
 sg13g2_decap_8 FILLER_6_736 ();
 sg13g2_decap_8 FILLER_6_743 ();
 sg13g2_decap_8 FILLER_6_750 ();
 sg13g2_decap_8 FILLER_6_757 ();
 sg13g2_decap_8 FILLER_6_764 ();
 sg13g2_decap_8 FILLER_6_771 ();
 sg13g2_decap_8 FILLER_6_778 ();
 sg13g2_decap_8 FILLER_6_785 ();
 sg13g2_decap_8 FILLER_6_792 ();
 sg13g2_decap_8 FILLER_6_799 ();
 sg13g2_decap_8 FILLER_6_806 ();
 sg13g2_decap_8 FILLER_6_813 ();
 sg13g2_decap_8 FILLER_6_820 ();
 sg13g2_decap_8 FILLER_6_827 ();
 sg13g2_decap_8 FILLER_6_834 ();
 sg13g2_decap_8 FILLER_6_841 ();
 sg13g2_decap_8 FILLER_6_848 ();
 sg13g2_decap_8 FILLER_6_855 ();
 sg13g2_decap_8 FILLER_6_862 ();
 sg13g2_decap_8 FILLER_6_869 ();
 sg13g2_decap_8 FILLER_6_876 ();
 sg13g2_decap_8 FILLER_6_883 ();
 sg13g2_decap_8 FILLER_6_890 ();
 sg13g2_decap_8 FILLER_6_897 ();
 sg13g2_decap_8 FILLER_6_904 ();
 sg13g2_decap_8 FILLER_6_911 ();
 sg13g2_decap_8 FILLER_6_918 ();
 sg13g2_decap_8 FILLER_6_925 ();
 sg13g2_decap_8 FILLER_6_932 ();
 sg13g2_decap_8 FILLER_6_939 ();
 sg13g2_decap_8 FILLER_6_946 ();
 sg13g2_decap_8 FILLER_6_953 ();
 sg13g2_decap_8 FILLER_6_960 ();
 sg13g2_decap_8 FILLER_6_967 ();
 sg13g2_decap_8 FILLER_6_974 ();
 sg13g2_decap_8 FILLER_6_981 ();
 sg13g2_decap_8 FILLER_6_988 ();
 sg13g2_decap_8 FILLER_6_995 ();
 sg13g2_decap_8 FILLER_6_1002 ();
 sg13g2_decap_8 FILLER_6_1009 ();
 sg13g2_decap_8 FILLER_6_1016 ();
 sg13g2_decap_4 FILLER_6_1023 ();
 sg13g2_fill_2 FILLER_6_1027 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_16 ();
 sg13g2_fill_1 FILLER_7_18 ();
 sg13g2_fill_2 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_41 ();
 sg13g2_fill_1 FILLER_7_47 ();
 sg13g2_decap_8 FILLER_7_53 ();
 sg13g2_decap_8 FILLER_7_60 ();
 sg13g2_decap_4 FILLER_7_67 ();
 sg13g2_fill_2 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_102 ();
 sg13g2_decap_4 FILLER_7_109 ();
 sg13g2_fill_1 FILLER_7_139 ();
 sg13g2_fill_2 FILLER_7_162 ();
 sg13g2_fill_1 FILLER_7_164 ();
 sg13g2_fill_2 FILLER_7_181 ();
 sg13g2_fill_1 FILLER_7_183 ();
 sg13g2_fill_2 FILLER_7_213 ();
 sg13g2_fill_2 FILLER_7_227 ();
 sg13g2_fill_1 FILLER_7_229 ();
 sg13g2_fill_2 FILLER_7_334 ();
 sg13g2_fill_1 FILLER_7_439 ();
 sg13g2_fill_2 FILLER_7_473 ();
 sg13g2_fill_1 FILLER_7_475 ();
 sg13g2_decap_8 FILLER_7_503 ();
 sg13g2_decap_8 FILLER_7_510 ();
 sg13g2_decap_8 FILLER_7_517 ();
 sg13g2_decap_8 FILLER_7_524 ();
 sg13g2_decap_8 FILLER_7_531 ();
 sg13g2_decap_8 FILLER_7_538 ();
 sg13g2_decap_8 FILLER_7_545 ();
 sg13g2_decap_8 FILLER_7_552 ();
 sg13g2_decap_8 FILLER_7_559 ();
 sg13g2_decap_8 FILLER_7_566 ();
 sg13g2_decap_8 FILLER_7_573 ();
 sg13g2_decap_8 FILLER_7_580 ();
 sg13g2_decap_8 FILLER_7_587 ();
 sg13g2_decap_8 FILLER_7_594 ();
 sg13g2_decap_8 FILLER_7_601 ();
 sg13g2_decap_8 FILLER_7_608 ();
 sg13g2_decap_8 FILLER_7_615 ();
 sg13g2_decap_8 FILLER_7_622 ();
 sg13g2_decap_8 FILLER_7_629 ();
 sg13g2_decap_8 FILLER_7_636 ();
 sg13g2_decap_8 FILLER_7_643 ();
 sg13g2_decap_8 FILLER_7_650 ();
 sg13g2_decap_8 FILLER_7_657 ();
 sg13g2_decap_8 FILLER_7_664 ();
 sg13g2_decap_8 FILLER_7_671 ();
 sg13g2_decap_8 FILLER_7_678 ();
 sg13g2_decap_8 FILLER_7_685 ();
 sg13g2_decap_8 FILLER_7_692 ();
 sg13g2_decap_8 FILLER_7_699 ();
 sg13g2_decap_8 FILLER_7_706 ();
 sg13g2_decap_8 FILLER_7_713 ();
 sg13g2_decap_8 FILLER_7_720 ();
 sg13g2_decap_8 FILLER_7_727 ();
 sg13g2_decap_8 FILLER_7_734 ();
 sg13g2_decap_8 FILLER_7_741 ();
 sg13g2_decap_8 FILLER_7_748 ();
 sg13g2_decap_8 FILLER_7_755 ();
 sg13g2_decap_8 FILLER_7_762 ();
 sg13g2_decap_8 FILLER_7_769 ();
 sg13g2_decap_8 FILLER_7_776 ();
 sg13g2_decap_8 FILLER_7_783 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_8 FILLER_7_797 ();
 sg13g2_decap_8 FILLER_7_804 ();
 sg13g2_decap_8 FILLER_7_811 ();
 sg13g2_decap_8 FILLER_7_818 ();
 sg13g2_decap_8 FILLER_7_825 ();
 sg13g2_decap_8 FILLER_7_832 ();
 sg13g2_decap_8 FILLER_7_839 ();
 sg13g2_decap_8 FILLER_7_846 ();
 sg13g2_decap_8 FILLER_7_853 ();
 sg13g2_decap_8 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_7_867 ();
 sg13g2_decap_8 FILLER_7_874 ();
 sg13g2_decap_8 FILLER_7_881 ();
 sg13g2_decap_8 FILLER_7_888 ();
 sg13g2_decap_8 FILLER_7_895 ();
 sg13g2_decap_8 FILLER_7_902 ();
 sg13g2_decap_8 FILLER_7_909 ();
 sg13g2_decap_8 FILLER_7_916 ();
 sg13g2_decap_8 FILLER_7_923 ();
 sg13g2_decap_8 FILLER_7_930 ();
 sg13g2_decap_8 FILLER_7_937 ();
 sg13g2_decap_8 FILLER_7_944 ();
 sg13g2_decap_8 FILLER_7_951 ();
 sg13g2_decap_8 FILLER_7_958 ();
 sg13g2_decap_8 FILLER_7_965 ();
 sg13g2_decap_8 FILLER_7_972 ();
 sg13g2_decap_8 FILLER_7_979 ();
 sg13g2_decap_8 FILLER_7_986 ();
 sg13g2_decap_8 FILLER_7_993 ();
 sg13g2_decap_8 FILLER_7_1000 ();
 sg13g2_decap_8 FILLER_7_1007 ();
 sg13g2_decap_8 FILLER_7_1014 ();
 sg13g2_decap_8 FILLER_7_1021 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_fill_2 FILLER_8_8 ();
 sg13g2_fill_2 FILLER_8_23 ();
 sg13g2_decap_4 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_46 ();
 sg13g2_fill_1 FILLER_8_64 ();
 sg13g2_fill_2 FILLER_8_79 ();
 sg13g2_decap_8 FILLER_8_87 ();
 sg13g2_decap_8 FILLER_8_94 ();
 sg13g2_decap_8 FILLER_8_101 ();
 sg13g2_fill_2 FILLER_8_108 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_fill_1 FILLER_8_122 ();
 sg13g2_fill_1 FILLER_8_186 ();
 sg13g2_fill_2 FILLER_8_233 ();
 sg13g2_fill_1 FILLER_8_235 ();
 sg13g2_fill_2 FILLER_8_262 ();
 sg13g2_fill_2 FILLER_8_384 ();
 sg13g2_fill_2 FILLER_8_391 ();
 sg13g2_fill_1 FILLER_8_441 ();
 sg13g2_fill_1 FILLER_8_460 ();
 sg13g2_decap_8 FILLER_8_503 ();
 sg13g2_decap_8 FILLER_8_510 ();
 sg13g2_decap_8 FILLER_8_517 ();
 sg13g2_decap_8 FILLER_8_524 ();
 sg13g2_decap_8 FILLER_8_531 ();
 sg13g2_decap_8 FILLER_8_538 ();
 sg13g2_decap_8 FILLER_8_545 ();
 sg13g2_decap_8 FILLER_8_552 ();
 sg13g2_decap_8 FILLER_8_559 ();
 sg13g2_decap_8 FILLER_8_566 ();
 sg13g2_decap_8 FILLER_8_573 ();
 sg13g2_decap_8 FILLER_8_580 ();
 sg13g2_decap_8 FILLER_8_587 ();
 sg13g2_decap_8 FILLER_8_594 ();
 sg13g2_decap_8 FILLER_8_601 ();
 sg13g2_decap_8 FILLER_8_608 ();
 sg13g2_decap_8 FILLER_8_615 ();
 sg13g2_decap_8 FILLER_8_622 ();
 sg13g2_decap_8 FILLER_8_629 ();
 sg13g2_decap_8 FILLER_8_636 ();
 sg13g2_decap_8 FILLER_8_643 ();
 sg13g2_decap_8 FILLER_8_650 ();
 sg13g2_decap_8 FILLER_8_657 ();
 sg13g2_decap_8 FILLER_8_664 ();
 sg13g2_decap_8 FILLER_8_671 ();
 sg13g2_decap_8 FILLER_8_678 ();
 sg13g2_decap_8 FILLER_8_685 ();
 sg13g2_decap_8 FILLER_8_692 ();
 sg13g2_decap_8 FILLER_8_699 ();
 sg13g2_decap_8 FILLER_8_706 ();
 sg13g2_decap_8 FILLER_8_713 ();
 sg13g2_decap_8 FILLER_8_720 ();
 sg13g2_decap_8 FILLER_8_727 ();
 sg13g2_decap_8 FILLER_8_734 ();
 sg13g2_decap_8 FILLER_8_741 ();
 sg13g2_decap_8 FILLER_8_748 ();
 sg13g2_decap_8 FILLER_8_755 ();
 sg13g2_decap_8 FILLER_8_762 ();
 sg13g2_decap_8 FILLER_8_769 ();
 sg13g2_decap_8 FILLER_8_776 ();
 sg13g2_decap_8 FILLER_8_783 ();
 sg13g2_decap_8 FILLER_8_790 ();
 sg13g2_decap_8 FILLER_8_797 ();
 sg13g2_decap_8 FILLER_8_804 ();
 sg13g2_decap_8 FILLER_8_811 ();
 sg13g2_decap_8 FILLER_8_818 ();
 sg13g2_decap_8 FILLER_8_825 ();
 sg13g2_decap_8 FILLER_8_832 ();
 sg13g2_decap_8 FILLER_8_839 ();
 sg13g2_decap_8 FILLER_8_846 ();
 sg13g2_decap_8 FILLER_8_853 ();
 sg13g2_decap_8 FILLER_8_860 ();
 sg13g2_decap_8 FILLER_8_867 ();
 sg13g2_decap_8 FILLER_8_874 ();
 sg13g2_decap_8 FILLER_8_881 ();
 sg13g2_decap_8 FILLER_8_888 ();
 sg13g2_decap_8 FILLER_8_895 ();
 sg13g2_decap_8 FILLER_8_902 ();
 sg13g2_decap_8 FILLER_8_909 ();
 sg13g2_decap_8 FILLER_8_916 ();
 sg13g2_decap_8 FILLER_8_923 ();
 sg13g2_decap_8 FILLER_8_930 ();
 sg13g2_decap_8 FILLER_8_937 ();
 sg13g2_decap_8 FILLER_8_944 ();
 sg13g2_decap_8 FILLER_8_951 ();
 sg13g2_decap_8 FILLER_8_958 ();
 sg13g2_decap_8 FILLER_8_965 ();
 sg13g2_decap_8 FILLER_8_972 ();
 sg13g2_decap_8 FILLER_8_979 ();
 sg13g2_decap_8 FILLER_8_986 ();
 sg13g2_decap_8 FILLER_8_993 ();
 sg13g2_decap_8 FILLER_8_1000 ();
 sg13g2_decap_8 FILLER_8_1007 ();
 sg13g2_decap_8 FILLER_8_1014 ();
 sg13g2_decap_8 FILLER_8_1021 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_fill_2 FILLER_9_4 ();
 sg13g2_fill_1 FILLER_9_6 ();
 sg13g2_fill_2 FILLER_9_40 ();
 sg13g2_fill_1 FILLER_9_51 ();
 sg13g2_decap_4 FILLER_9_80 ();
 sg13g2_decap_4 FILLER_9_92 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_fill_2 FILLER_9_123 ();
 sg13g2_fill_1 FILLER_9_153 ();
 sg13g2_fill_2 FILLER_9_163 ();
 sg13g2_fill_1 FILLER_9_165 ();
 sg13g2_fill_1 FILLER_9_188 ();
 sg13g2_fill_2 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_205 ();
 sg13g2_fill_2 FILLER_9_212 ();
 sg13g2_fill_1 FILLER_9_214 ();
 sg13g2_fill_1 FILLER_9_220 ();
 sg13g2_fill_2 FILLER_9_298 ();
 sg13g2_fill_1 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_384 ();
 sg13g2_fill_1 FILLER_9_415 ();
 sg13g2_fill_2 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_9_488 ();
 sg13g2_decap_8 FILLER_9_495 ();
 sg13g2_decap_8 FILLER_9_502 ();
 sg13g2_decap_8 FILLER_9_509 ();
 sg13g2_decap_8 FILLER_9_516 ();
 sg13g2_decap_8 FILLER_9_523 ();
 sg13g2_decap_8 FILLER_9_530 ();
 sg13g2_decap_8 FILLER_9_537 ();
 sg13g2_decap_8 FILLER_9_544 ();
 sg13g2_decap_8 FILLER_9_551 ();
 sg13g2_decap_8 FILLER_9_558 ();
 sg13g2_decap_8 FILLER_9_565 ();
 sg13g2_decap_8 FILLER_9_572 ();
 sg13g2_decap_8 FILLER_9_579 ();
 sg13g2_decap_8 FILLER_9_586 ();
 sg13g2_decap_8 FILLER_9_593 ();
 sg13g2_decap_8 FILLER_9_600 ();
 sg13g2_decap_8 FILLER_9_607 ();
 sg13g2_decap_8 FILLER_9_614 ();
 sg13g2_decap_8 FILLER_9_621 ();
 sg13g2_decap_8 FILLER_9_628 ();
 sg13g2_decap_8 FILLER_9_635 ();
 sg13g2_decap_8 FILLER_9_642 ();
 sg13g2_decap_8 FILLER_9_649 ();
 sg13g2_decap_8 FILLER_9_656 ();
 sg13g2_decap_8 FILLER_9_663 ();
 sg13g2_decap_8 FILLER_9_670 ();
 sg13g2_decap_8 FILLER_9_677 ();
 sg13g2_decap_8 FILLER_9_684 ();
 sg13g2_decap_8 FILLER_9_691 ();
 sg13g2_decap_8 FILLER_9_698 ();
 sg13g2_decap_8 FILLER_9_705 ();
 sg13g2_decap_8 FILLER_9_712 ();
 sg13g2_decap_8 FILLER_9_719 ();
 sg13g2_decap_8 FILLER_9_726 ();
 sg13g2_decap_8 FILLER_9_733 ();
 sg13g2_decap_8 FILLER_9_740 ();
 sg13g2_decap_8 FILLER_9_747 ();
 sg13g2_decap_8 FILLER_9_754 ();
 sg13g2_decap_8 FILLER_9_761 ();
 sg13g2_decap_8 FILLER_9_768 ();
 sg13g2_decap_8 FILLER_9_775 ();
 sg13g2_decap_8 FILLER_9_782 ();
 sg13g2_decap_8 FILLER_9_789 ();
 sg13g2_decap_8 FILLER_9_796 ();
 sg13g2_decap_8 FILLER_9_803 ();
 sg13g2_decap_8 FILLER_9_810 ();
 sg13g2_decap_8 FILLER_9_817 ();
 sg13g2_decap_8 FILLER_9_824 ();
 sg13g2_decap_8 FILLER_9_831 ();
 sg13g2_decap_8 FILLER_9_838 ();
 sg13g2_decap_8 FILLER_9_845 ();
 sg13g2_decap_8 FILLER_9_852 ();
 sg13g2_decap_8 FILLER_9_859 ();
 sg13g2_decap_8 FILLER_9_866 ();
 sg13g2_decap_8 FILLER_9_873 ();
 sg13g2_decap_8 FILLER_9_880 ();
 sg13g2_decap_8 FILLER_9_887 ();
 sg13g2_decap_8 FILLER_9_894 ();
 sg13g2_decap_8 FILLER_9_901 ();
 sg13g2_decap_8 FILLER_9_908 ();
 sg13g2_decap_8 FILLER_9_915 ();
 sg13g2_decap_8 FILLER_9_922 ();
 sg13g2_decap_8 FILLER_9_929 ();
 sg13g2_decap_8 FILLER_9_936 ();
 sg13g2_decap_8 FILLER_9_943 ();
 sg13g2_decap_8 FILLER_9_950 ();
 sg13g2_decap_8 FILLER_9_957 ();
 sg13g2_decap_8 FILLER_9_964 ();
 sg13g2_decap_8 FILLER_9_971 ();
 sg13g2_decap_8 FILLER_9_978 ();
 sg13g2_decap_8 FILLER_9_985 ();
 sg13g2_decap_8 FILLER_9_992 ();
 sg13g2_decap_8 FILLER_9_999 ();
 sg13g2_decap_8 FILLER_9_1006 ();
 sg13g2_decap_8 FILLER_9_1013 ();
 sg13g2_decap_8 FILLER_9_1020 ();
 sg13g2_fill_2 FILLER_9_1027 ();
 sg13g2_fill_1 FILLER_10_32 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_fill_1 FILLER_10_64 ();
 sg13g2_fill_2 FILLER_10_120 ();
 sg13g2_fill_1 FILLER_10_122 ();
 sg13g2_fill_2 FILLER_10_133 ();
 sg13g2_fill_2 FILLER_10_154 ();
 sg13g2_fill_2 FILLER_10_166 ();
 sg13g2_fill_1 FILLER_10_168 ();
 sg13g2_fill_1 FILLER_10_174 ();
 sg13g2_fill_2 FILLER_10_188 ();
 sg13g2_fill_1 FILLER_10_190 ();
 sg13g2_fill_2 FILLER_10_213 ();
 sg13g2_fill_2 FILLER_10_261 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_312 ();
 sg13g2_fill_1 FILLER_10_353 ();
 sg13g2_fill_2 FILLER_10_391 ();
 sg13g2_fill_1 FILLER_10_441 ();
 sg13g2_fill_1 FILLER_10_450 ();
 sg13g2_decap_8 FILLER_10_503 ();
 sg13g2_decap_8 FILLER_10_510 ();
 sg13g2_decap_8 FILLER_10_517 ();
 sg13g2_decap_8 FILLER_10_524 ();
 sg13g2_decap_8 FILLER_10_531 ();
 sg13g2_decap_8 FILLER_10_538 ();
 sg13g2_decap_8 FILLER_10_545 ();
 sg13g2_decap_8 FILLER_10_552 ();
 sg13g2_decap_8 FILLER_10_559 ();
 sg13g2_decap_8 FILLER_10_566 ();
 sg13g2_decap_8 FILLER_10_573 ();
 sg13g2_decap_8 FILLER_10_580 ();
 sg13g2_decap_8 FILLER_10_587 ();
 sg13g2_decap_8 FILLER_10_594 ();
 sg13g2_decap_8 FILLER_10_601 ();
 sg13g2_decap_8 FILLER_10_608 ();
 sg13g2_decap_8 FILLER_10_615 ();
 sg13g2_decap_8 FILLER_10_622 ();
 sg13g2_decap_8 FILLER_10_629 ();
 sg13g2_decap_8 FILLER_10_636 ();
 sg13g2_decap_8 FILLER_10_643 ();
 sg13g2_decap_8 FILLER_10_650 ();
 sg13g2_decap_8 FILLER_10_657 ();
 sg13g2_decap_8 FILLER_10_664 ();
 sg13g2_decap_8 FILLER_10_671 ();
 sg13g2_decap_8 FILLER_10_678 ();
 sg13g2_decap_8 FILLER_10_685 ();
 sg13g2_decap_8 FILLER_10_692 ();
 sg13g2_decap_8 FILLER_10_699 ();
 sg13g2_decap_8 FILLER_10_706 ();
 sg13g2_decap_8 FILLER_10_713 ();
 sg13g2_decap_8 FILLER_10_720 ();
 sg13g2_decap_8 FILLER_10_727 ();
 sg13g2_decap_8 FILLER_10_734 ();
 sg13g2_decap_8 FILLER_10_741 ();
 sg13g2_decap_8 FILLER_10_748 ();
 sg13g2_decap_8 FILLER_10_755 ();
 sg13g2_decap_8 FILLER_10_762 ();
 sg13g2_decap_8 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_776 ();
 sg13g2_decap_8 FILLER_10_783 ();
 sg13g2_decap_8 FILLER_10_790 ();
 sg13g2_decap_8 FILLER_10_797 ();
 sg13g2_decap_8 FILLER_10_804 ();
 sg13g2_decap_8 FILLER_10_811 ();
 sg13g2_decap_8 FILLER_10_818 ();
 sg13g2_decap_8 FILLER_10_825 ();
 sg13g2_decap_8 FILLER_10_832 ();
 sg13g2_decap_8 FILLER_10_839 ();
 sg13g2_decap_8 FILLER_10_846 ();
 sg13g2_decap_8 FILLER_10_853 ();
 sg13g2_decap_8 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_10_867 ();
 sg13g2_decap_8 FILLER_10_874 ();
 sg13g2_decap_8 FILLER_10_881 ();
 sg13g2_decap_8 FILLER_10_888 ();
 sg13g2_decap_8 FILLER_10_895 ();
 sg13g2_decap_8 FILLER_10_902 ();
 sg13g2_decap_8 FILLER_10_909 ();
 sg13g2_decap_8 FILLER_10_916 ();
 sg13g2_decap_8 FILLER_10_923 ();
 sg13g2_decap_8 FILLER_10_930 ();
 sg13g2_decap_8 FILLER_10_937 ();
 sg13g2_decap_8 FILLER_10_944 ();
 sg13g2_decap_8 FILLER_10_951 ();
 sg13g2_decap_8 FILLER_10_958 ();
 sg13g2_decap_8 FILLER_10_965 ();
 sg13g2_decap_8 FILLER_10_972 ();
 sg13g2_decap_8 FILLER_10_979 ();
 sg13g2_decap_8 FILLER_10_986 ();
 sg13g2_decap_8 FILLER_10_993 ();
 sg13g2_decap_8 FILLER_10_1000 ();
 sg13g2_decap_8 FILLER_10_1007 ();
 sg13g2_decap_8 FILLER_10_1014 ();
 sg13g2_decap_8 FILLER_10_1021 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_fill_1 FILLER_11_63 ();
 sg13g2_fill_2 FILLER_11_68 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_fill_1 FILLER_11_88 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_138 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_fill_1 FILLER_11_169 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_261 ();
 sg13g2_fill_2 FILLER_11_275 ();
 sg13g2_fill_2 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_450 ();
 sg13g2_fill_1 FILLER_11_465 ();
 sg13g2_decap_8 FILLER_11_501 ();
 sg13g2_decap_8 FILLER_11_508 ();
 sg13g2_decap_8 FILLER_11_515 ();
 sg13g2_decap_8 FILLER_11_522 ();
 sg13g2_decap_8 FILLER_11_529 ();
 sg13g2_decap_8 FILLER_11_536 ();
 sg13g2_decap_8 FILLER_11_543 ();
 sg13g2_decap_8 FILLER_11_550 ();
 sg13g2_decap_8 FILLER_11_557 ();
 sg13g2_decap_8 FILLER_11_564 ();
 sg13g2_decap_8 FILLER_11_571 ();
 sg13g2_decap_8 FILLER_11_578 ();
 sg13g2_decap_8 FILLER_11_585 ();
 sg13g2_decap_8 FILLER_11_592 ();
 sg13g2_decap_8 FILLER_11_599 ();
 sg13g2_decap_8 FILLER_11_606 ();
 sg13g2_decap_8 FILLER_11_613 ();
 sg13g2_decap_8 FILLER_11_620 ();
 sg13g2_decap_8 FILLER_11_627 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_662 ();
 sg13g2_decap_8 FILLER_11_669 ();
 sg13g2_decap_8 FILLER_11_676 ();
 sg13g2_decap_8 FILLER_11_683 ();
 sg13g2_decap_8 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_decap_8 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_decap_8 FILLER_11_739 ();
 sg13g2_decap_8 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_753 ();
 sg13g2_decap_8 FILLER_11_760 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_8 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_11_865 ();
 sg13g2_decap_8 FILLER_11_872 ();
 sg13g2_decap_8 FILLER_11_879 ();
 sg13g2_decap_8 FILLER_11_886 ();
 sg13g2_decap_8 FILLER_11_893 ();
 sg13g2_decap_8 FILLER_11_900 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_914 ();
 sg13g2_decap_8 FILLER_11_921 ();
 sg13g2_decap_8 FILLER_11_928 ();
 sg13g2_decap_8 FILLER_11_935 ();
 sg13g2_decap_8 FILLER_11_942 ();
 sg13g2_decap_8 FILLER_11_949 ();
 sg13g2_decap_8 FILLER_11_956 ();
 sg13g2_decap_8 FILLER_11_963 ();
 sg13g2_decap_8 FILLER_11_970 ();
 sg13g2_decap_8 FILLER_11_977 ();
 sg13g2_decap_8 FILLER_11_984 ();
 sg13g2_decap_8 FILLER_11_991 ();
 sg13g2_decap_8 FILLER_11_998 ();
 sg13g2_decap_8 FILLER_11_1005 ();
 sg13g2_decap_8 FILLER_11_1012 ();
 sg13g2_decap_8 FILLER_11_1019 ();
 sg13g2_fill_2 FILLER_11_1026 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_fill_2 FILLER_12_33 ();
 sg13g2_fill_2 FILLER_12_60 ();
 sg13g2_fill_1 FILLER_12_62 ();
 sg13g2_fill_2 FILLER_12_73 ();
 sg13g2_fill_1 FILLER_12_75 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_fill_2 FILLER_12_107 ();
 sg13g2_fill_1 FILLER_12_109 ();
 sg13g2_fill_2 FILLER_12_123 ();
 sg13g2_fill_1 FILLER_12_125 ();
 sg13g2_fill_2 FILLER_12_149 ();
 sg13g2_fill_1 FILLER_12_151 ();
 sg13g2_fill_2 FILLER_12_228 ();
 sg13g2_fill_1 FILLER_12_240 ();
 sg13g2_fill_2 FILLER_12_325 ();
 sg13g2_fill_1 FILLER_12_327 ();
 sg13g2_fill_2 FILLER_12_366 ();
 sg13g2_fill_2 FILLER_12_420 ();
 sg13g2_fill_1 FILLER_12_447 ();
 sg13g2_fill_1 FILLER_12_453 ();
 sg13g2_fill_1 FILLER_12_468 ();
 sg13g2_fill_1 FILLER_12_477 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_decap_8 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_12_868 ();
 sg13g2_decap_8 FILLER_12_875 ();
 sg13g2_decap_8 FILLER_12_882 ();
 sg13g2_decap_8 FILLER_12_889 ();
 sg13g2_decap_8 FILLER_12_896 ();
 sg13g2_decap_8 FILLER_12_903 ();
 sg13g2_decap_8 FILLER_12_910 ();
 sg13g2_decap_8 FILLER_12_917 ();
 sg13g2_decap_8 FILLER_12_924 ();
 sg13g2_decap_8 FILLER_12_931 ();
 sg13g2_decap_8 FILLER_12_938 ();
 sg13g2_decap_8 FILLER_12_945 ();
 sg13g2_decap_8 FILLER_12_952 ();
 sg13g2_decap_8 FILLER_12_959 ();
 sg13g2_decap_8 FILLER_12_966 ();
 sg13g2_decap_8 FILLER_12_973 ();
 sg13g2_decap_8 FILLER_12_980 ();
 sg13g2_decap_8 FILLER_12_987 ();
 sg13g2_decap_8 FILLER_12_994 ();
 sg13g2_decap_8 FILLER_12_1001 ();
 sg13g2_decap_8 FILLER_12_1008 ();
 sg13g2_decap_8 FILLER_12_1015 ();
 sg13g2_decap_8 FILLER_12_1022 ();
 sg13g2_fill_2 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_46 ();
 sg13g2_fill_2 FILLER_13_64 ();
 sg13g2_fill_1 FILLER_13_106 ();
 sg13g2_fill_2 FILLER_13_127 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_fill_2 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_181 ();
 sg13g2_fill_2 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_239 ();
 sg13g2_fill_2 FILLER_13_271 ();
 sg13g2_fill_2 FILLER_13_291 ();
 sg13g2_fill_1 FILLER_13_293 ();
 sg13g2_fill_2 FILLER_13_300 ();
 sg13g2_fill_1 FILLER_13_302 ();
 sg13g2_fill_1 FILLER_13_330 ();
 sg13g2_fill_1 FILLER_13_368 ();
 sg13g2_fill_1 FILLER_13_424 ();
 sg13g2_fill_1 FILLER_13_458 ();
 sg13g2_fill_1 FILLER_13_467 ();
 sg13g2_decap_8 FILLER_13_502 ();
 sg13g2_decap_8 FILLER_13_509 ();
 sg13g2_decap_8 FILLER_13_516 ();
 sg13g2_decap_8 FILLER_13_523 ();
 sg13g2_decap_8 FILLER_13_530 ();
 sg13g2_decap_8 FILLER_13_537 ();
 sg13g2_decap_8 FILLER_13_544 ();
 sg13g2_decap_8 FILLER_13_551 ();
 sg13g2_decap_8 FILLER_13_558 ();
 sg13g2_decap_8 FILLER_13_565 ();
 sg13g2_decap_8 FILLER_13_572 ();
 sg13g2_decap_8 FILLER_13_579 ();
 sg13g2_decap_8 FILLER_13_586 ();
 sg13g2_decap_8 FILLER_13_593 ();
 sg13g2_decap_8 FILLER_13_600 ();
 sg13g2_decap_8 FILLER_13_607 ();
 sg13g2_decap_8 FILLER_13_614 ();
 sg13g2_decap_8 FILLER_13_621 ();
 sg13g2_decap_8 FILLER_13_628 ();
 sg13g2_decap_8 FILLER_13_635 ();
 sg13g2_decap_8 FILLER_13_642 ();
 sg13g2_decap_8 FILLER_13_649 ();
 sg13g2_decap_8 FILLER_13_656 ();
 sg13g2_decap_8 FILLER_13_663 ();
 sg13g2_decap_8 FILLER_13_670 ();
 sg13g2_decap_8 FILLER_13_677 ();
 sg13g2_decap_8 FILLER_13_684 ();
 sg13g2_decap_8 FILLER_13_691 ();
 sg13g2_decap_8 FILLER_13_698 ();
 sg13g2_decap_8 FILLER_13_705 ();
 sg13g2_decap_8 FILLER_13_712 ();
 sg13g2_decap_8 FILLER_13_719 ();
 sg13g2_decap_8 FILLER_13_726 ();
 sg13g2_decap_8 FILLER_13_733 ();
 sg13g2_decap_8 FILLER_13_740 ();
 sg13g2_decap_8 FILLER_13_747 ();
 sg13g2_decap_8 FILLER_13_754 ();
 sg13g2_decap_8 FILLER_13_761 ();
 sg13g2_decap_8 FILLER_13_768 ();
 sg13g2_decap_8 FILLER_13_775 ();
 sg13g2_decap_8 FILLER_13_782 ();
 sg13g2_decap_8 FILLER_13_789 ();
 sg13g2_decap_8 FILLER_13_796 ();
 sg13g2_decap_8 FILLER_13_803 ();
 sg13g2_decap_8 FILLER_13_810 ();
 sg13g2_decap_8 FILLER_13_817 ();
 sg13g2_decap_8 FILLER_13_824 ();
 sg13g2_decap_8 FILLER_13_831 ();
 sg13g2_decap_8 FILLER_13_838 ();
 sg13g2_decap_8 FILLER_13_845 ();
 sg13g2_decap_8 FILLER_13_852 ();
 sg13g2_decap_8 FILLER_13_859 ();
 sg13g2_decap_8 FILLER_13_866 ();
 sg13g2_decap_8 FILLER_13_873 ();
 sg13g2_decap_8 FILLER_13_880 ();
 sg13g2_decap_8 FILLER_13_887 ();
 sg13g2_decap_8 FILLER_13_894 ();
 sg13g2_decap_8 FILLER_13_901 ();
 sg13g2_decap_8 FILLER_13_908 ();
 sg13g2_decap_8 FILLER_13_915 ();
 sg13g2_decap_8 FILLER_13_922 ();
 sg13g2_decap_8 FILLER_13_929 ();
 sg13g2_decap_8 FILLER_13_936 ();
 sg13g2_decap_8 FILLER_13_943 ();
 sg13g2_decap_8 FILLER_13_950 ();
 sg13g2_decap_8 FILLER_13_957 ();
 sg13g2_decap_8 FILLER_13_964 ();
 sg13g2_decap_8 FILLER_13_971 ();
 sg13g2_decap_8 FILLER_13_978 ();
 sg13g2_decap_8 FILLER_13_985 ();
 sg13g2_decap_8 FILLER_13_992 ();
 sg13g2_decap_8 FILLER_13_999 ();
 sg13g2_decap_8 FILLER_13_1006 ();
 sg13g2_decap_8 FILLER_13_1013 ();
 sg13g2_decap_8 FILLER_13_1020 ();
 sg13g2_fill_2 FILLER_13_1027 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_fill_2 FILLER_14_117 ();
 sg13g2_fill_1 FILLER_14_119 ();
 sg13g2_fill_2 FILLER_14_139 ();
 sg13g2_fill_1 FILLER_14_141 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_fill_2 FILLER_14_246 ();
 sg13g2_fill_1 FILLER_14_248 ();
 sg13g2_fill_2 FILLER_14_271 ();
 sg13g2_fill_1 FILLER_14_283 ();
 sg13g2_fill_2 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_337 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_fill_1 FILLER_14_354 ();
 sg13g2_fill_2 FILLER_14_369 ();
 sg13g2_fill_2 FILLER_14_400 ();
 sg13g2_fill_1 FILLER_14_407 ();
 sg13g2_fill_1 FILLER_14_415 ();
 sg13g2_fill_2 FILLER_14_421 ();
 sg13g2_fill_1 FILLER_14_423 ();
 sg13g2_fill_1 FILLER_14_460 ();
 sg13g2_decap_8 FILLER_14_488 ();
 sg13g2_decap_8 FILLER_14_495 ();
 sg13g2_decap_8 FILLER_14_502 ();
 sg13g2_decap_8 FILLER_14_509 ();
 sg13g2_decap_8 FILLER_14_516 ();
 sg13g2_decap_8 FILLER_14_523 ();
 sg13g2_decap_8 FILLER_14_530 ();
 sg13g2_decap_8 FILLER_14_537 ();
 sg13g2_decap_8 FILLER_14_544 ();
 sg13g2_decap_8 FILLER_14_551 ();
 sg13g2_decap_8 FILLER_14_558 ();
 sg13g2_decap_8 FILLER_14_565 ();
 sg13g2_decap_8 FILLER_14_572 ();
 sg13g2_decap_8 FILLER_14_579 ();
 sg13g2_decap_8 FILLER_14_586 ();
 sg13g2_decap_8 FILLER_14_593 ();
 sg13g2_decap_8 FILLER_14_600 ();
 sg13g2_decap_8 FILLER_14_607 ();
 sg13g2_decap_8 FILLER_14_614 ();
 sg13g2_decap_8 FILLER_14_621 ();
 sg13g2_decap_8 FILLER_14_628 ();
 sg13g2_decap_8 FILLER_14_635 ();
 sg13g2_decap_8 FILLER_14_642 ();
 sg13g2_decap_8 FILLER_14_649 ();
 sg13g2_decap_8 FILLER_14_656 ();
 sg13g2_decap_8 FILLER_14_663 ();
 sg13g2_decap_8 FILLER_14_670 ();
 sg13g2_decap_8 FILLER_14_677 ();
 sg13g2_decap_8 FILLER_14_684 ();
 sg13g2_decap_8 FILLER_14_691 ();
 sg13g2_decap_8 FILLER_14_698 ();
 sg13g2_decap_8 FILLER_14_705 ();
 sg13g2_decap_8 FILLER_14_712 ();
 sg13g2_decap_8 FILLER_14_719 ();
 sg13g2_decap_8 FILLER_14_726 ();
 sg13g2_decap_8 FILLER_14_733 ();
 sg13g2_decap_8 FILLER_14_740 ();
 sg13g2_decap_8 FILLER_14_747 ();
 sg13g2_decap_8 FILLER_14_754 ();
 sg13g2_decap_8 FILLER_14_761 ();
 sg13g2_decap_8 FILLER_14_768 ();
 sg13g2_decap_8 FILLER_14_775 ();
 sg13g2_decap_8 FILLER_14_782 ();
 sg13g2_decap_8 FILLER_14_789 ();
 sg13g2_decap_8 FILLER_14_796 ();
 sg13g2_decap_8 FILLER_14_803 ();
 sg13g2_decap_8 FILLER_14_810 ();
 sg13g2_decap_8 FILLER_14_817 ();
 sg13g2_decap_8 FILLER_14_824 ();
 sg13g2_decap_8 FILLER_14_831 ();
 sg13g2_decap_8 FILLER_14_838 ();
 sg13g2_decap_8 FILLER_14_845 ();
 sg13g2_decap_8 FILLER_14_852 ();
 sg13g2_decap_8 FILLER_14_859 ();
 sg13g2_decap_8 FILLER_14_866 ();
 sg13g2_decap_8 FILLER_14_873 ();
 sg13g2_decap_8 FILLER_14_880 ();
 sg13g2_decap_8 FILLER_14_887 ();
 sg13g2_decap_8 FILLER_14_894 ();
 sg13g2_decap_8 FILLER_14_901 ();
 sg13g2_decap_8 FILLER_14_908 ();
 sg13g2_decap_8 FILLER_14_915 ();
 sg13g2_decap_8 FILLER_14_922 ();
 sg13g2_decap_8 FILLER_14_929 ();
 sg13g2_decap_8 FILLER_14_936 ();
 sg13g2_decap_8 FILLER_14_943 ();
 sg13g2_decap_8 FILLER_14_950 ();
 sg13g2_decap_8 FILLER_14_957 ();
 sg13g2_decap_8 FILLER_14_964 ();
 sg13g2_decap_8 FILLER_14_971 ();
 sg13g2_decap_8 FILLER_14_978 ();
 sg13g2_decap_8 FILLER_14_985 ();
 sg13g2_decap_8 FILLER_14_992 ();
 sg13g2_decap_8 FILLER_14_999 ();
 sg13g2_decap_8 FILLER_14_1006 ();
 sg13g2_decap_8 FILLER_14_1013 ();
 sg13g2_decap_8 FILLER_14_1020 ();
 sg13g2_fill_2 FILLER_14_1027 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_57 ();
 sg13g2_fill_2 FILLER_15_106 ();
 sg13g2_fill_2 FILLER_15_115 ();
 sg13g2_fill_2 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_168 ();
 sg13g2_fill_1 FILLER_15_170 ();
 sg13g2_fill_1 FILLER_15_178 ();
 sg13g2_fill_1 FILLER_15_186 ();
 sg13g2_fill_1 FILLER_15_209 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_fill_1 FILLER_15_226 ();
 sg13g2_fill_2 FILLER_15_303 ();
 sg13g2_fill_2 FILLER_15_314 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_fill_2 FILLER_15_393 ();
 sg13g2_fill_2 FILLER_15_414 ();
 sg13g2_fill_2 FILLER_15_433 ();
 sg13g2_fill_1 FILLER_15_435 ();
 sg13g2_fill_2 FILLER_15_461 ();
 sg13g2_fill_1 FILLER_15_463 ();
 sg13g2_decap_8 FILLER_15_507 ();
 sg13g2_decap_8 FILLER_15_514 ();
 sg13g2_decap_8 FILLER_15_521 ();
 sg13g2_decap_8 FILLER_15_528 ();
 sg13g2_decap_8 FILLER_15_535 ();
 sg13g2_decap_8 FILLER_15_542 ();
 sg13g2_decap_8 FILLER_15_549 ();
 sg13g2_decap_8 FILLER_15_556 ();
 sg13g2_decap_8 FILLER_15_563 ();
 sg13g2_decap_8 FILLER_15_570 ();
 sg13g2_decap_8 FILLER_15_577 ();
 sg13g2_decap_8 FILLER_15_584 ();
 sg13g2_decap_8 FILLER_15_591 ();
 sg13g2_decap_8 FILLER_15_598 ();
 sg13g2_decap_8 FILLER_15_605 ();
 sg13g2_decap_8 FILLER_15_612 ();
 sg13g2_decap_8 FILLER_15_619 ();
 sg13g2_decap_8 FILLER_15_626 ();
 sg13g2_decap_8 FILLER_15_633 ();
 sg13g2_decap_8 FILLER_15_640 ();
 sg13g2_decap_8 FILLER_15_647 ();
 sg13g2_decap_8 FILLER_15_654 ();
 sg13g2_decap_8 FILLER_15_661 ();
 sg13g2_decap_8 FILLER_15_668 ();
 sg13g2_decap_8 FILLER_15_675 ();
 sg13g2_decap_8 FILLER_15_682 ();
 sg13g2_decap_8 FILLER_15_689 ();
 sg13g2_decap_8 FILLER_15_696 ();
 sg13g2_decap_8 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_710 ();
 sg13g2_decap_8 FILLER_15_717 ();
 sg13g2_decap_8 FILLER_15_724 ();
 sg13g2_decap_8 FILLER_15_731 ();
 sg13g2_decap_8 FILLER_15_738 ();
 sg13g2_decap_8 FILLER_15_745 ();
 sg13g2_decap_8 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_759 ();
 sg13g2_decap_8 FILLER_15_766 ();
 sg13g2_decap_8 FILLER_15_773 ();
 sg13g2_decap_8 FILLER_15_780 ();
 sg13g2_decap_8 FILLER_15_787 ();
 sg13g2_decap_8 FILLER_15_794 ();
 sg13g2_decap_8 FILLER_15_801 ();
 sg13g2_decap_8 FILLER_15_808 ();
 sg13g2_decap_8 FILLER_15_815 ();
 sg13g2_decap_8 FILLER_15_822 ();
 sg13g2_decap_8 FILLER_15_829 ();
 sg13g2_decap_8 FILLER_15_836 ();
 sg13g2_decap_8 FILLER_15_843 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_decap_8 FILLER_15_857 ();
 sg13g2_decap_8 FILLER_15_864 ();
 sg13g2_decap_8 FILLER_15_871 ();
 sg13g2_decap_8 FILLER_15_878 ();
 sg13g2_decap_8 FILLER_15_885 ();
 sg13g2_decap_8 FILLER_15_892 ();
 sg13g2_decap_8 FILLER_15_899 ();
 sg13g2_decap_8 FILLER_15_906 ();
 sg13g2_decap_8 FILLER_15_913 ();
 sg13g2_decap_8 FILLER_15_920 ();
 sg13g2_decap_8 FILLER_15_927 ();
 sg13g2_decap_8 FILLER_15_934 ();
 sg13g2_decap_8 FILLER_15_941 ();
 sg13g2_decap_8 FILLER_15_948 ();
 sg13g2_decap_8 FILLER_15_955 ();
 sg13g2_decap_8 FILLER_15_962 ();
 sg13g2_decap_8 FILLER_15_969 ();
 sg13g2_decap_8 FILLER_15_976 ();
 sg13g2_decap_8 FILLER_15_983 ();
 sg13g2_decap_8 FILLER_15_990 ();
 sg13g2_decap_8 FILLER_15_997 ();
 sg13g2_decap_8 FILLER_15_1004 ();
 sg13g2_decap_8 FILLER_15_1011 ();
 sg13g2_decap_8 FILLER_15_1018 ();
 sg13g2_decap_4 FILLER_15_1025 ();
 sg13g2_fill_1 FILLER_16_58 ();
 sg13g2_fill_2 FILLER_16_85 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_138 ();
 sg13g2_fill_1 FILLER_16_140 ();
 sg13g2_fill_1 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_171 ();
 sg13g2_fill_1 FILLER_16_173 ();
 sg13g2_fill_2 FILLER_16_193 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_fill_2 FILLER_16_329 ();
 sg13g2_fill_1 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_fill_1 FILLER_16_377 ();
 sg13g2_fill_1 FILLER_16_412 ();
 sg13g2_fill_2 FILLER_16_440 ();
 sg13g2_fill_1 FILLER_16_442 ();
 sg13g2_fill_1 FILLER_16_448 ();
 sg13g2_fill_2 FILLER_16_464 ();
 sg13g2_decap_8 FILLER_16_508 ();
 sg13g2_decap_8 FILLER_16_515 ();
 sg13g2_decap_8 FILLER_16_522 ();
 sg13g2_decap_8 FILLER_16_529 ();
 sg13g2_decap_8 FILLER_16_536 ();
 sg13g2_decap_8 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_550 ();
 sg13g2_decap_8 FILLER_16_557 ();
 sg13g2_decap_8 FILLER_16_564 ();
 sg13g2_decap_8 FILLER_16_571 ();
 sg13g2_decap_8 FILLER_16_578 ();
 sg13g2_decap_8 FILLER_16_585 ();
 sg13g2_decap_8 FILLER_16_592 ();
 sg13g2_decap_8 FILLER_16_599 ();
 sg13g2_decap_8 FILLER_16_606 ();
 sg13g2_decap_8 FILLER_16_613 ();
 sg13g2_decap_8 FILLER_16_620 ();
 sg13g2_decap_8 FILLER_16_627 ();
 sg13g2_decap_8 FILLER_16_634 ();
 sg13g2_decap_8 FILLER_16_641 ();
 sg13g2_decap_8 FILLER_16_648 ();
 sg13g2_decap_8 FILLER_16_655 ();
 sg13g2_decap_8 FILLER_16_662 ();
 sg13g2_decap_8 FILLER_16_669 ();
 sg13g2_decap_8 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_683 ();
 sg13g2_decap_8 FILLER_16_690 ();
 sg13g2_decap_8 FILLER_16_697 ();
 sg13g2_decap_8 FILLER_16_704 ();
 sg13g2_decap_8 FILLER_16_711 ();
 sg13g2_decap_8 FILLER_16_718 ();
 sg13g2_decap_8 FILLER_16_725 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_decap_8 FILLER_16_753 ();
 sg13g2_decap_8 FILLER_16_760 ();
 sg13g2_decap_8 FILLER_16_767 ();
 sg13g2_decap_8 FILLER_16_774 ();
 sg13g2_decap_8 FILLER_16_781 ();
 sg13g2_decap_8 FILLER_16_788 ();
 sg13g2_decap_8 FILLER_16_795 ();
 sg13g2_decap_8 FILLER_16_802 ();
 sg13g2_decap_8 FILLER_16_809 ();
 sg13g2_decap_8 FILLER_16_816 ();
 sg13g2_decap_8 FILLER_16_823 ();
 sg13g2_decap_8 FILLER_16_830 ();
 sg13g2_decap_8 FILLER_16_837 ();
 sg13g2_decap_8 FILLER_16_844 ();
 sg13g2_decap_8 FILLER_16_851 ();
 sg13g2_decap_8 FILLER_16_858 ();
 sg13g2_decap_8 FILLER_16_865 ();
 sg13g2_decap_8 FILLER_16_872 ();
 sg13g2_decap_8 FILLER_16_879 ();
 sg13g2_decap_8 FILLER_16_886 ();
 sg13g2_decap_8 FILLER_16_893 ();
 sg13g2_decap_8 FILLER_16_900 ();
 sg13g2_decap_8 FILLER_16_907 ();
 sg13g2_decap_8 FILLER_16_914 ();
 sg13g2_decap_8 FILLER_16_921 ();
 sg13g2_decap_8 FILLER_16_928 ();
 sg13g2_decap_8 FILLER_16_935 ();
 sg13g2_decap_8 FILLER_16_942 ();
 sg13g2_decap_8 FILLER_16_949 ();
 sg13g2_decap_8 FILLER_16_956 ();
 sg13g2_decap_8 FILLER_16_963 ();
 sg13g2_decap_8 FILLER_16_970 ();
 sg13g2_decap_8 FILLER_16_977 ();
 sg13g2_decap_8 FILLER_16_984 ();
 sg13g2_decap_8 FILLER_16_991 ();
 sg13g2_decap_8 FILLER_16_998 ();
 sg13g2_decap_8 FILLER_16_1005 ();
 sg13g2_decap_8 FILLER_16_1012 ();
 sg13g2_decap_8 FILLER_16_1019 ();
 sg13g2_fill_2 FILLER_16_1026 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_fill_2 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_75 ();
 sg13g2_fill_2 FILLER_17_89 ();
 sg13g2_fill_1 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_fill_2 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_fill_1 FILLER_17_337 ();
 sg13g2_fill_2 FILLER_17_351 ();
 sg13g2_fill_2 FILLER_17_405 ();
 sg13g2_fill_2 FILLER_17_460 ();
 sg13g2_fill_1 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_507 ();
 sg13g2_decap_8 FILLER_17_514 ();
 sg13g2_decap_8 FILLER_17_521 ();
 sg13g2_decap_8 FILLER_17_528 ();
 sg13g2_decap_8 FILLER_17_535 ();
 sg13g2_decap_8 FILLER_17_542 ();
 sg13g2_decap_8 FILLER_17_549 ();
 sg13g2_decap_8 FILLER_17_556 ();
 sg13g2_decap_8 FILLER_17_563 ();
 sg13g2_decap_8 FILLER_17_570 ();
 sg13g2_decap_8 FILLER_17_577 ();
 sg13g2_decap_8 FILLER_17_584 ();
 sg13g2_decap_8 FILLER_17_591 ();
 sg13g2_decap_8 FILLER_17_598 ();
 sg13g2_decap_8 FILLER_17_605 ();
 sg13g2_decap_8 FILLER_17_612 ();
 sg13g2_decap_8 FILLER_17_619 ();
 sg13g2_decap_8 FILLER_17_626 ();
 sg13g2_decap_8 FILLER_17_633 ();
 sg13g2_decap_8 FILLER_17_640 ();
 sg13g2_decap_8 FILLER_17_647 ();
 sg13g2_decap_8 FILLER_17_654 ();
 sg13g2_decap_8 FILLER_17_661 ();
 sg13g2_decap_8 FILLER_17_668 ();
 sg13g2_decap_8 FILLER_17_675 ();
 sg13g2_decap_8 FILLER_17_682 ();
 sg13g2_decap_8 FILLER_17_689 ();
 sg13g2_decap_8 FILLER_17_696 ();
 sg13g2_decap_8 FILLER_17_703 ();
 sg13g2_decap_8 FILLER_17_710 ();
 sg13g2_decap_8 FILLER_17_717 ();
 sg13g2_decap_8 FILLER_17_724 ();
 sg13g2_decap_8 FILLER_17_731 ();
 sg13g2_decap_8 FILLER_17_738 ();
 sg13g2_decap_8 FILLER_17_745 ();
 sg13g2_decap_8 FILLER_17_752 ();
 sg13g2_decap_8 FILLER_17_759 ();
 sg13g2_decap_8 FILLER_17_766 ();
 sg13g2_decap_8 FILLER_17_773 ();
 sg13g2_decap_8 FILLER_17_780 ();
 sg13g2_decap_8 FILLER_17_787 ();
 sg13g2_decap_8 FILLER_17_794 ();
 sg13g2_decap_8 FILLER_17_801 ();
 sg13g2_decap_8 FILLER_17_808 ();
 sg13g2_decap_8 FILLER_17_815 ();
 sg13g2_decap_8 FILLER_17_822 ();
 sg13g2_decap_8 FILLER_17_829 ();
 sg13g2_decap_8 FILLER_17_836 ();
 sg13g2_decap_8 FILLER_17_843 ();
 sg13g2_decap_8 FILLER_17_850 ();
 sg13g2_decap_8 FILLER_17_857 ();
 sg13g2_decap_8 FILLER_17_864 ();
 sg13g2_decap_8 FILLER_17_871 ();
 sg13g2_decap_8 FILLER_17_878 ();
 sg13g2_decap_8 FILLER_17_885 ();
 sg13g2_decap_8 FILLER_17_892 ();
 sg13g2_decap_8 FILLER_17_899 ();
 sg13g2_decap_8 FILLER_17_906 ();
 sg13g2_decap_8 FILLER_17_913 ();
 sg13g2_decap_8 FILLER_17_920 ();
 sg13g2_decap_8 FILLER_17_927 ();
 sg13g2_decap_8 FILLER_17_934 ();
 sg13g2_decap_8 FILLER_17_941 ();
 sg13g2_decap_8 FILLER_17_948 ();
 sg13g2_decap_8 FILLER_17_955 ();
 sg13g2_decap_8 FILLER_17_962 ();
 sg13g2_decap_8 FILLER_17_969 ();
 sg13g2_decap_8 FILLER_17_976 ();
 sg13g2_decap_8 FILLER_17_983 ();
 sg13g2_decap_8 FILLER_17_990 ();
 sg13g2_decap_8 FILLER_17_997 ();
 sg13g2_decap_8 FILLER_17_1004 ();
 sg13g2_decap_8 FILLER_17_1011 ();
 sg13g2_decap_8 FILLER_17_1018 ();
 sg13g2_decap_4 FILLER_17_1025 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_264 ();
 sg13g2_fill_2 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_430 ();
 sg13g2_fill_2 FILLER_18_473 ();
 sg13g2_decap_8 FILLER_18_502 ();
 sg13g2_decap_8 FILLER_18_509 ();
 sg13g2_decap_8 FILLER_18_516 ();
 sg13g2_decap_8 FILLER_18_523 ();
 sg13g2_decap_8 FILLER_18_530 ();
 sg13g2_decap_8 FILLER_18_537 ();
 sg13g2_decap_8 FILLER_18_544 ();
 sg13g2_decap_8 FILLER_18_551 ();
 sg13g2_decap_8 FILLER_18_558 ();
 sg13g2_decap_8 FILLER_18_565 ();
 sg13g2_decap_8 FILLER_18_572 ();
 sg13g2_decap_8 FILLER_18_579 ();
 sg13g2_decap_8 FILLER_18_586 ();
 sg13g2_decap_8 FILLER_18_593 ();
 sg13g2_decap_8 FILLER_18_600 ();
 sg13g2_decap_8 FILLER_18_607 ();
 sg13g2_decap_8 FILLER_18_614 ();
 sg13g2_decap_8 FILLER_18_621 ();
 sg13g2_decap_8 FILLER_18_628 ();
 sg13g2_decap_8 FILLER_18_635 ();
 sg13g2_decap_8 FILLER_18_642 ();
 sg13g2_decap_8 FILLER_18_649 ();
 sg13g2_decap_8 FILLER_18_656 ();
 sg13g2_decap_8 FILLER_18_663 ();
 sg13g2_decap_8 FILLER_18_670 ();
 sg13g2_decap_8 FILLER_18_677 ();
 sg13g2_decap_8 FILLER_18_684 ();
 sg13g2_decap_8 FILLER_18_691 ();
 sg13g2_decap_8 FILLER_18_698 ();
 sg13g2_decap_8 FILLER_18_705 ();
 sg13g2_decap_8 FILLER_18_712 ();
 sg13g2_decap_8 FILLER_18_719 ();
 sg13g2_decap_8 FILLER_18_726 ();
 sg13g2_decap_8 FILLER_18_733 ();
 sg13g2_decap_8 FILLER_18_740 ();
 sg13g2_decap_8 FILLER_18_747 ();
 sg13g2_decap_8 FILLER_18_754 ();
 sg13g2_decap_8 FILLER_18_761 ();
 sg13g2_decap_8 FILLER_18_768 ();
 sg13g2_decap_8 FILLER_18_775 ();
 sg13g2_decap_8 FILLER_18_782 ();
 sg13g2_decap_8 FILLER_18_789 ();
 sg13g2_decap_8 FILLER_18_796 ();
 sg13g2_decap_8 FILLER_18_803 ();
 sg13g2_decap_8 FILLER_18_810 ();
 sg13g2_decap_8 FILLER_18_817 ();
 sg13g2_decap_8 FILLER_18_824 ();
 sg13g2_decap_8 FILLER_18_831 ();
 sg13g2_decap_8 FILLER_18_838 ();
 sg13g2_decap_8 FILLER_18_845 ();
 sg13g2_decap_8 FILLER_18_852 ();
 sg13g2_decap_8 FILLER_18_859 ();
 sg13g2_decap_8 FILLER_18_866 ();
 sg13g2_decap_8 FILLER_18_873 ();
 sg13g2_decap_8 FILLER_18_880 ();
 sg13g2_decap_8 FILLER_18_887 ();
 sg13g2_decap_8 FILLER_18_894 ();
 sg13g2_decap_8 FILLER_18_901 ();
 sg13g2_decap_8 FILLER_18_908 ();
 sg13g2_decap_8 FILLER_18_915 ();
 sg13g2_decap_8 FILLER_18_922 ();
 sg13g2_decap_8 FILLER_18_929 ();
 sg13g2_decap_8 FILLER_18_936 ();
 sg13g2_decap_8 FILLER_18_943 ();
 sg13g2_decap_8 FILLER_18_950 ();
 sg13g2_decap_8 FILLER_18_957 ();
 sg13g2_decap_8 FILLER_18_964 ();
 sg13g2_decap_8 FILLER_18_971 ();
 sg13g2_decap_8 FILLER_18_978 ();
 sg13g2_decap_8 FILLER_18_985 ();
 sg13g2_decap_8 FILLER_18_992 ();
 sg13g2_decap_8 FILLER_18_999 ();
 sg13g2_decap_8 FILLER_18_1006 ();
 sg13g2_decap_8 FILLER_18_1013 ();
 sg13g2_decap_8 FILLER_18_1020 ();
 sg13g2_fill_2 FILLER_18_1027 ();
 sg13g2_fill_2 FILLER_19_76 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_decap_4 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_212 ();
 sg13g2_fill_2 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_392 ();
 sg13g2_fill_1 FILLER_19_424 ();
 sg13g2_fill_1 FILLER_19_461 ();
 sg13g2_decap_8 FILLER_19_488 ();
 sg13g2_decap_8 FILLER_19_495 ();
 sg13g2_decap_8 FILLER_19_502 ();
 sg13g2_decap_8 FILLER_19_509 ();
 sg13g2_decap_8 FILLER_19_516 ();
 sg13g2_decap_8 FILLER_19_523 ();
 sg13g2_decap_8 FILLER_19_530 ();
 sg13g2_decap_8 FILLER_19_537 ();
 sg13g2_decap_8 FILLER_19_544 ();
 sg13g2_decap_8 FILLER_19_551 ();
 sg13g2_decap_8 FILLER_19_558 ();
 sg13g2_decap_8 FILLER_19_565 ();
 sg13g2_decap_8 FILLER_19_572 ();
 sg13g2_decap_8 FILLER_19_579 ();
 sg13g2_decap_8 FILLER_19_586 ();
 sg13g2_decap_8 FILLER_19_593 ();
 sg13g2_decap_8 FILLER_19_600 ();
 sg13g2_decap_8 FILLER_19_607 ();
 sg13g2_decap_8 FILLER_19_614 ();
 sg13g2_decap_8 FILLER_19_621 ();
 sg13g2_decap_8 FILLER_19_628 ();
 sg13g2_decap_8 FILLER_19_635 ();
 sg13g2_decap_8 FILLER_19_642 ();
 sg13g2_decap_8 FILLER_19_649 ();
 sg13g2_decap_8 FILLER_19_656 ();
 sg13g2_decap_8 FILLER_19_663 ();
 sg13g2_decap_8 FILLER_19_670 ();
 sg13g2_decap_8 FILLER_19_677 ();
 sg13g2_decap_8 FILLER_19_684 ();
 sg13g2_decap_8 FILLER_19_691 ();
 sg13g2_decap_8 FILLER_19_698 ();
 sg13g2_decap_8 FILLER_19_705 ();
 sg13g2_decap_8 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_719 ();
 sg13g2_decap_8 FILLER_19_726 ();
 sg13g2_decap_8 FILLER_19_733 ();
 sg13g2_decap_8 FILLER_19_740 ();
 sg13g2_decap_8 FILLER_19_747 ();
 sg13g2_decap_8 FILLER_19_754 ();
 sg13g2_decap_8 FILLER_19_761 ();
 sg13g2_decap_8 FILLER_19_768 ();
 sg13g2_decap_8 FILLER_19_775 ();
 sg13g2_decap_8 FILLER_19_782 ();
 sg13g2_decap_8 FILLER_19_789 ();
 sg13g2_decap_8 FILLER_19_796 ();
 sg13g2_decap_8 FILLER_19_803 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_decap_8 FILLER_19_817 ();
 sg13g2_decap_8 FILLER_19_824 ();
 sg13g2_decap_8 FILLER_19_831 ();
 sg13g2_decap_8 FILLER_19_838 ();
 sg13g2_decap_8 FILLER_19_845 ();
 sg13g2_decap_8 FILLER_19_852 ();
 sg13g2_decap_8 FILLER_19_859 ();
 sg13g2_decap_8 FILLER_19_866 ();
 sg13g2_decap_8 FILLER_19_873 ();
 sg13g2_decap_8 FILLER_19_880 ();
 sg13g2_decap_8 FILLER_19_887 ();
 sg13g2_decap_8 FILLER_19_894 ();
 sg13g2_decap_8 FILLER_19_901 ();
 sg13g2_decap_8 FILLER_19_908 ();
 sg13g2_decap_8 FILLER_19_915 ();
 sg13g2_decap_8 FILLER_19_922 ();
 sg13g2_decap_8 FILLER_19_929 ();
 sg13g2_decap_8 FILLER_19_936 ();
 sg13g2_decap_8 FILLER_19_943 ();
 sg13g2_decap_8 FILLER_19_950 ();
 sg13g2_decap_8 FILLER_19_957 ();
 sg13g2_decap_8 FILLER_19_964 ();
 sg13g2_decap_8 FILLER_19_971 ();
 sg13g2_decap_8 FILLER_19_978 ();
 sg13g2_decap_8 FILLER_19_985 ();
 sg13g2_decap_8 FILLER_19_992 ();
 sg13g2_decap_8 FILLER_19_999 ();
 sg13g2_decap_8 FILLER_19_1006 ();
 sg13g2_decap_8 FILLER_19_1013 ();
 sg13g2_decap_8 FILLER_19_1020 ();
 sg13g2_fill_2 FILLER_19_1027 ();
 sg13g2_fill_2 FILLER_20_9 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_457 ();
 sg13g2_decap_8 FILLER_20_485 ();
 sg13g2_decap_8 FILLER_20_492 ();
 sg13g2_decap_8 FILLER_20_499 ();
 sg13g2_decap_8 FILLER_20_506 ();
 sg13g2_decap_8 FILLER_20_513 ();
 sg13g2_decap_8 FILLER_20_520 ();
 sg13g2_decap_8 FILLER_20_527 ();
 sg13g2_decap_8 FILLER_20_534 ();
 sg13g2_decap_8 FILLER_20_541 ();
 sg13g2_decap_8 FILLER_20_548 ();
 sg13g2_decap_8 FILLER_20_555 ();
 sg13g2_decap_8 FILLER_20_562 ();
 sg13g2_decap_8 FILLER_20_569 ();
 sg13g2_decap_8 FILLER_20_576 ();
 sg13g2_decap_8 FILLER_20_583 ();
 sg13g2_decap_8 FILLER_20_590 ();
 sg13g2_decap_8 FILLER_20_597 ();
 sg13g2_decap_8 FILLER_20_604 ();
 sg13g2_decap_8 FILLER_20_611 ();
 sg13g2_decap_8 FILLER_20_618 ();
 sg13g2_decap_8 FILLER_20_625 ();
 sg13g2_decap_8 FILLER_20_632 ();
 sg13g2_decap_8 FILLER_20_639 ();
 sg13g2_decap_8 FILLER_20_646 ();
 sg13g2_decap_8 FILLER_20_653 ();
 sg13g2_decap_8 FILLER_20_660 ();
 sg13g2_decap_8 FILLER_20_667 ();
 sg13g2_decap_8 FILLER_20_674 ();
 sg13g2_decap_8 FILLER_20_681 ();
 sg13g2_decap_8 FILLER_20_688 ();
 sg13g2_decap_8 FILLER_20_695 ();
 sg13g2_decap_8 FILLER_20_702 ();
 sg13g2_decap_8 FILLER_20_709 ();
 sg13g2_decap_8 FILLER_20_716 ();
 sg13g2_decap_8 FILLER_20_723 ();
 sg13g2_decap_8 FILLER_20_730 ();
 sg13g2_decap_8 FILLER_20_737 ();
 sg13g2_decap_8 FILLER_20_744 ();
 sg13g2_decap_8 FILLER_20_751 ();
 sg13g2_decap_8 FILLER_20_758 ();
 sg13g2_decap_8 FILLER_20_765 ();
 sg13g2_decap_8 FILLER_20_772 ();
 sg13g2_decap_8 FILLER_20_779 ();
 sg13g2_decap_8 FILLER_20_786 ();
 sg13g2_decap_8 FILLER_20_793 ();
 sg13g2_decap_8 FILLER_20_800 ();
 sg13g2_decap_8 FILLER_20_807 ();
 sg13g2_decap_8 FILLER_20_814 ();
 sg13g2_decap_8 FILLER_20_821 ();
 sg13g2_decap_8 FILLER_20_828 ();
 sg13g2_decap_8 FILLER_20_835 ();
 sg13g2_decap_8 FILLER_20_842 ();
 sg13g2_decap_8 FILLER_20_849 ();
 sg13g2_decap_8 FILLER_20_856 ();
 sg13g2_decap_8 FILLER_20_863 ();
 sg13g2_decap_8 FILLER_20_870 ();
 sg13g2_decap_8 FILLER_20_877 ();
 sg13g2_decap_8 FILLER_20_884 ();
 sg13g2_decap_8 FILLER_20_891 ();
 sg13g2_decap_8 FILLER_20_898 ();
 sg13g2_decap_8 FILLER_20_905 ();
 sg13g2_decap_8 FILLER_20_912 ();
 sg13g2_decap_8 FILLER_20_919 ();
 sg13g2_decap_8 FILLER_20_926 ();
 sg13g2_decap_8 FILLER_20_933 ();
 sg13g2_decap_8 FILLER_20_940 ();
 sg13g2_decap_8 FILLER_20_947 ();
 sg13g2_decap_8 FILLER_20_954 ();
 sg13g2_decap_8 FILLER_20_961 ();
 sg13g2_decap_8 FILLER_20_968 ();
 sg13g2_decap_8 FILLER_20_975 ();
 sg13g2_decap_8 FILLER_20_982 ();
 sg13g2_decap_8 FILLER_20_989 ();
 sg13g2_decap_8 FILLER_20_996 ();
 sg13g2_decap_8 FILLER_20_1003 ();
 sg13g2_decap_8 FILLER_20_1010 ();
 sg13g2_decap_8 FILLER_20_1017 ();
 sg13g2_decap_4 FILLER_20_1024 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_132 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_360 ();
 sg13g2_fill_2 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_376 ();
 sg13g2_fill_2 FILLER_21_421 ();
 sg13g2_decap_8 FILLER_21_478 ();
 sg13g2_decap_8 FILLER_21_485 ();
 sg13g2_decap_8 FILLER_21_492 ();
 sg13g2_decap_8 FILLER_21_499 ();
 sg13g2_decap_8 FILLER_21_506 ();
 sg13g2_decap_8 FILLER_21_513 ();
 sg13g2_decap_8 FILLER_21_520 ();
 sg13g2_decap_8 FILLER_21_527 ();
 sg13g2_decap_8 FILLER_21_534 ();
 sg13g2_decap_8 FILLER_21_541 ();
 sg13g2_decap_8 FILLER_21_548 ();
 sg13g2_decap_8 FILLER_21_555 ();
 sg13g2_decap_8 FILLER_21_562 ();
 sg13g2_decap_8 FILLER_21_569 ();
 sg13g2_decap_8 FILLER_21_576 ();
 sg13g2_decap_8 FILLER_21_583 ();
 sg13g2_decap_8 FILLER_21_590 ();
 sg13g2_decap_8 FILLER_21_597 ();
 sg13g2_decap_8 FILLER_21_604 ();
 sg13g2_decap_8 FILLER_21_611 ();
 sg13g2_decap_8 FILLER_21_618 ();
 sg13g2_decap_8 FILLER_21_625 ();
 sg13g2_decap_8 FILLER_21_632 ();
 sg13g2_decap_8 FILLER_21_639 ();
 sg13g2_decap_8 FILLER_21_646 ();
 sg13g2_decap_8 FILLER_21_653 ();
 sg13g2_decap_8 FILLER_21_660 ();
 sg13g2_decap_8 FILLER_21_667 ();
 sg13g2_decap_8 FILLER_21_674 ();
 sg13g2_decap_8 FILLER_21_681 ();
 sg13g2_decap_8 FILLER_21_688 ();
 sg13g2_decap_8 FILLER_21_695 ();
 sg13g2_decap_8 FILLER_21_702 ();
 sg13g2_decap_8 FILLER_21_709 ();
 sg13g2_decap_8 FILLER_21_716 ();
 sg13g2_decap_8 FILLER_21_723 ();
 sg13g2_decap_8 FILLER_21_730 ();
 sg13g2_decap_8 FILLER_21_737 ();
 sg13g2_decap_8 FILLER_21_744 ();
 sg13g2_decap_8 FILLER_21_751 ();
 sg13g2_decap_8 FILLER_21_758 ();
 sg13g2_decap_8 FILLER_21_765 ();
 sg13g2_decap_8 FILLER_21_772 ();
 sg13g2_decap_8 FILLER_21_779 ();
 sg13g2_decap_8 FILLER_21_786 ();
 sg13g2_decap_8 FILLER_21_793 ();
 sg13g2_decap_8 FILLER_21_800 ();
 sg13g2_decap_8 FILLER_21_807 ();
 sg13g2_decap_8 FILLER_21_814 ();
 sg13g2_decap_8 FILLER_21_821 ();
 sg13g2_decap_8 FILLER_21_828 ();
 sg13g2_decap_8 FILLER_21_835 ();
 sg13g2_decap_8 FILLER_21_842 ();
 sg13g2_decap_8 FILLER_21_849 ();
 sg13g2_decap_8 FILLER_21_856 ();
 sg13g2_decap_8 FILLER_21_863 ();
 sg13g2_decap_8 FILLER_21_870 ();
 sg13g2_decap_8 FILLER_21_877 ();
 sg13g2_decap_8 FILLER_21_884 ();
 sg13g2_decap_8 FILLER_21_891 ();
 sg13g2_decap_8 FILLER_21_898 ();
 sg13g2_decap_8 FILLER_21_905 ();
 sg13g2_decap_8 FILLER_21_912 ();
 sg13g2_decap_8 FILLER_21_919 ();
 sg13g2_decap_8 FILLER_21_926 ();
 sg13g2_decap_8 FILLER_21_933 ();
 sg13g2_decap_8 FILLER_21_940 ();
 sg13g2_decap_8 FILLER_21_947 ();
 sg13g2_decap_8 FILLER_21_954 ();
 sg13g2_decap_8 FILLER_21_961 ();
 sg13g2_decap_8 FILLER_21_968 ();
 sg13g2_decap_8 FILLER_21_975 ();
 sg13g2_decap_8 FILLER_21_982 ();
 sg13g2_decap_8 FILLER_21_989 ();
 sg13g2_decap_8 FILLER_21_996 ();
 sg13g2_decap_8 FILLER_21_1003 ();
 sg13g2_decap_8 FILLER_21_1010 ();
 sg13g2_decap_8 FILLER_21_1017 ();
 sg13g2_decap_4 FILLER_21_1024 ();
 sg13g2_fill_1 FILLER_21_1028 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_108 ();
 sg13g2_fill_2 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_158 ();
 sg13g2_fill_2 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_328 ();
 sg13g2_fill_1 FILLER_22_346 ();
 sg13g2_decap_4 FILLER_22_375 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_fill_1 FILLER_22_409 ();
 sg13g2_fill_2 FILLER_22_443 ();
 sg13g2_decap_8 FILLER_22_463 ();
 sg13g2_decap_8 FILLER_22_470 ();
 sg13g2_decap_8 FILLER_22_477 ();
 sg13g2_decap_8 FILLER_22_484 ();
 sg13g2_decap_8 FILLER_22_491 ();
 sg13g2_decap_8 FILLER_22_498 ();
 sg13g2_decap_8 FILLER_22_505 ();
 sg13g2_decap_8 FILLER_22_512 ();
 sg13g2_decap_8 FILLER_22_519 ();
 sg13g2_decap_8 FILLER_22_526 ();
 sg13g2_decap_8 FILLER_22_533 ();
 sg13g2_decap_8 FILLER_22_540 ();
 sg13g2_decap_8 FILLER_22_547 ();
 sg13g2_decap_8 FILLER_22_554 ();
 sg13g2_decap_8 FILLER_22_561 ();
 sg13g2_decap_8 FILLER_22_568 ();
 sg13g2_decap_8 FILLER_22_575 ();
 sg13g2_decap_8 FILLER_22_582 ();
 sg13g2_decap_8 FILLER_22_589 ();
 sg13g2_decap_8 FILLER_22_596 ();
 sg13g2_decap_8 FILLER_22_603 ();
 sg13g2_decap_8 FILLER_22_610 ();
 sg13g2_decap_8 FILLER_22_617 ();
 sg13g2_decap_8 FILLER_22_624 ();
 sg13g2_decap_8 FILLER_22_631 ();
 sg13g2_decap_8 FILLER_22_638 ();
 sg13g2_decap_8 FILLER_22_645 ();
 sg13g2_decap_8 FILLER_22_652 ();
 sg13g2_decap_8 FILLER_22_659 ();
 sg13g2_decap_8 FILLER_22_666 ();
 sg13g2_decap_8 FILLER_22_673 ();
 sg13g2_decap_8 FILLER_22_680 ();
 sg13g2_decap_8 FILLER_22_687 ();
 sg13g2_decap_8 FILLER_22_694 ();
 sg13g2_decap_8 FILLER_22_701 ();
 sg13g2_decap_8 FILLER_22_708 ();
 sg13g2_decap_8 FILLER_22_715 ();
 sg13g2_decap_8 FILLER_22_722 ();
 sg13g2_decap_8 FILLER_22_729 ();
 sg13g2_decap_8 FILLER_22_736 ();
 sg13g2_decap_8 FILLER_22_743 ();
 sg13g2_decap_8 FILLER_22_750 ();
 sg13g2_decap_8 FILLER_22_757 ();
 sg13g2_decap_8 FILLER_22_764 ();
 sg13g2_decap_8 FILLER_22_771 ();
 sg13g2_decap_8 FILLER_22_778 ();
 sg13g2_decap_8 FILLER_22_785 ();
 sg13g2_decap_8 FILLER_22_792 ();
 sg13g2_decap_8 FILLER_22_799 ();
 sg13g2_decap_8 FILLER_22_806 ();
 sg13g2_decap_8 FILLER_22_813 ();
 sg13g2_decap_8 FILLER_22_820 ();
 sg13g2_decap_8 FILLER_22_827 ();
 sg13g2_decap_8 FILLER_22_834 ();
 sg13g2_decap_8 FILLER_22_841 ();
 sg13g2_decap_8 FILLER_22_848 ();
 sg13g2_decap_8 FILLER_22_855 ();
 sg13g2_decap_8 FILLER_22_862 ();
 sg13g2_decap_8 FILLER_22_869 ();
 sg13g2_decap_8 FILLER_22_876 ();
 sg13g2_decap_8 FILLER_22_883 ();
 sg13g2_decap_8 FILLER_22_890 ();
 sg13g2_decap_8 FILLER_22_897 ();
 sg13g2_decap_8 FILLER_22_904 ();
 sg13g2_decap_8 FILLER_22_911 ();
 sg13g2_decap_8 FILLER_22_918 ();
 sg13g2_decap_8 FILLER_22_925 ();
 sg13g2_decap_8 FILLER_22_932 ();
 sg13g2_decap_8 FILLER_22_939 ();
 sg13g2_decap_8 FILLER_22_946 ();
 sg13g2_decap_8 FILLER_22_953 ();
 sg13g2_decap_8 FILLER_22_960 ();
 sg13g2_decap_8 FILLER_22_967 ();
 sg13g2_decap_8 FILLER_22_974 ();
 sg13g2_decap_8 FILLER_22_981 ();
 sg13g2_decap_8 FILLER_22_988 ();
 sg13g2_decap_8 FILLER_22_995 ();
 sg13g2_decap_8 FILLER_22_1002 ();
 sg13g2_decap_8 FILLER_22_1009 ();
 sg13g2_decap_8 FILLER_22_1016 ();
 sg13g2_decap_4 FILLER_22_1023 ();
 sg13g2_fill_2 FILLER_22_1027 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_fill_1 FILLER_23_33 ();
 sg13g2_fill_2 FILLER_23_39 ();
 sg13g2_fill_2 FILLER_23_52 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_151 ();
 sg13g2_decap_4 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_186 ();
 sg13g2_decap_4 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_282 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_fill_2 FILLER_23_311 ();
 sg13g2_decap_4 FILLER_23_374 ();
 sg13g2_decap_4 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_decap_4 FILLER_23_407 ();
 sg13g2_fill_2 FILLER_23_411 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_decap_8 FILLER_23_424 ();
 sg13g2_decap_8 FILLER_23_431 ();
 sg13g2_decap_8 FILLER_23_438 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_fill_2 FILLER_23_452 ();
 sg13g2_decap_8 FILLER_23_458 ();
 sg13g2_decap_8 FILLER_23_465 ();
 sg13g2_decap_8 FILLER_23_472 ();
 sg13g2_decap_8 FILLER_23_479 ();
 sg13g2_decap_8 FILLER_23_486 ();
 sg13g2_decap_8 FILLER_23_493 ();
 sg13g2_decap_8 FILLER_23_500 ();
 sg13g2_decap_8 FILLER_23_507 ();
 sg13g2_decap_8 FILLER_23_514 ();
 sg13g2_decap_8 FILLER_23_521 ();
 sg13g2_decap_8 FILLER_23_528 ();
 sg13g2_decap_8 FILLER_23_535 ();
 sg13g2_decap_8 FILLER_23_542 ();
 sg13g2_decap_8 FILLER_23_549 ();
 sg13g2_decap_8 FILLER_23_556 ();
 sg13g2_decap_8 FILLER_23_563 ();
 sg13g2_decap_8 FILLER_23_570 ();
 sg13g2_decap_8 FILLER_23_577 ();
 sg13g2_decap_8 FILLER_23_584 ();
 sg13g2_decap_8 FILLER_23_591 ();
 sg13g2_decap_8 FILLER_23_598 ();
 sg13g2_decap_8 FILLER_23_605 ();
 sg13g2_decap_8 FILLER_23_612 ();
 sg13g2_decap_8 FILLER_23_619 ();
 sg13g2_decap_8 FILLER_23_626 ();
 sg13g2_decap_8 FILLER_23_633 ();
 sg13g2_decap_8 FILLER_23_640 ();
 sg13g2_decap_8 FILLER_23_647 ();
 sg13g2_decap_8 FILLER_23_654 ();
 sg13g2_decap_8 FILLER_23_661 ();
 sg13g2_decap_8 FILLER_23_668 ();
 sg13g2_decap_8 FILLER_23_675 ();
 sg13g2_decap_8 FILLER_23_682 ();
 sg13g2_decap_8 FILLER_23_689 ();
 sg13g2_decap_8 FILLER_23_696 ();
 sg13g2_decap_8 FILLER_23_703 ();
 sg13g2_decap_8 FILLER_23_710 ();
 sg13g2_decap_8 FILLER_23_717 ();
 sg13g2_decap_8 FILLER_23_724 ();
 sg13g2_decap_8 FILLER_23_731 ();
 sg13g2_decap_8 FILLER_23_738 ();
 sg13g2_decap_8 FILLER_23_745 ();
 sg13g2_decap_8 FILLER_23_752 ();
 sg13g2_decap_8 FILLER_23_759 ();
 sg13g2_decap_8 FILLER_23_766 ();
 sg13g2_decap_8 FILLER_23_773 ();
 sg13g2_decap_8 FILLER_23_780 ();
 sg13g2_decap_8 FILLER_23_787 ();
 sg13g2_decap_8 FILLER_23_794 ();
 sg13g2_decap_8 FILLER_23_801 ();
 sg13g2_decap_8 FILLER_23_808 ();
 sg13g2_decap_8 FILLER_23_815 ();
 sg13g2_decap_8 FILLER_23_822 ();
 sg13g2_decap_8 FILLER_23_829 ();
 sg13g2_decap_8 FILLER_23_836 ();
 sg13g2_decap_8 FILLER_23_843 ();
 sg13g2_decap_8 FILLER_23_850 ();
 sg13g2_decap_8 FILLER_23_857 ();
 sg13g2_decap_8 FILLER_23_864 ();
 sg13g2_decap_8 FILLER_23_871 ();
 sg13g2_decap_8 FILLER_23_878 ();
 sg13g2_decap_8 FILLER_23_885 ();
 sg13g2_decap_8 FILLER_23_892 ();
 sg13g2_decap_8 FILLER_23_899 ();
 sg13g2_decap_8 FILLER_23_906 ();
 sg13g2_decap_8 FILLER_23_913 ();
 sg13g2_decap_8 FILLER_23_920 ();
 sg13g2_decap_8 FILLER_23_927 ();
 sg13g2_decap_8 FILLER_23_934 ();
 sg13g2_decap_8 FILLER_23_941 ();
 sg13g2_decap_8 FILLER_23_948 ();
 sg13g2_decap_8 FILLER_23_955 ();
 sg13g2_decap_8 FILLER_23_962 ();
 sg13g2_decap_8 FILLER_23_969 ();
 sg13g2_decap_8 FILLER_23_976 ();
 sg13g2_decap_8 FILLER_23_983 ();
 sg13g2_decap_8 FILLER_23_990 ();
 sg13g2_decap_8 FILLER_23_997 ();
 sg13g2_decap_8 FILLER_23_1004 ();
 sg13g2_decap_8 FILLER_23_1011 ();
 sg13g2_decap_8 FILLER_23_1018 ();
 sg13g2_decap_4 FILLER_23_1025 ();
 sg13g2_fill_1 FILLER_24_8 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_fill_2 FILLER_24_110 ();
 sg13g2_fill_1 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_181 ();
 sg13g2_decap_4 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_decap_8 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_24_414 ();
 sg13g2_decap_8 FILLER_24_421 ();
 sg13g2_decap_8 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_24_435 ();
 sg13g2_decap_8 FILLER_24_442 ();
 sg13g2_decap_8 FILLER_24_449 ();
 sg13g2_decap_8 FILLER_24_456 ();
 sg13g2_decap_8 FILLER_24_463 ();
 sg13g2_decap_8 FILLER_24_470 ();
 sg13g2_decap_8 FILLER_24_477 ();
 sg13g2_decap_8 FILLER_24_484 ();
 sg13g2_decap_8 FILLER_24_491 ();
 sg13g2_decap_8 FILLER_24_498 ();
 sg13g2_decap_8 FILLER_24_505 ();
 sg13g2_decap_8 FILLER_24_512 ();
 sg13g2_decap_8 FILLER_24_519 ();
 sg13g2_decap_8 FILLER_24_526 ();
 sg13g2_decap_8 FILLER_24_533 ();
 sg13g2_decap_8 FILLER_24_540 ();
 sg13g2_decap_8 FILLER_24_547 ();
 sg13g2_decap_8 FILLER_24_554 ();
 sg13g2_decap_8 FILLER_24_561 ();
 sg13g2_decap_8 FILLER_24_568 ();
 sg13g2_decap_8 FILLER_24_575 ();
 sg13g2_decap_8 FILLER_24_582 ();
 sg13g2_decap_8 FILLER_24_589 ();
 sg13g2_decap_8 FILLER_24_596 ();
 sg13g2_decap_8 FILLER_24_603 ();
 sg13g2_decap_8 FILLER_24_610 ();
 sg13g2_decap_8 FILLER_24_617 ();
 sg13g2_decap_8 FILLER_24_624 ();
 sg13g2_decap_8 FILLER_24_631 ();
 sg13g2_decap_8 FILLER_24_638 ();
 sg13g2_decap_8 FILLER_24_645 ();
 sg13g2_decap_8 FILLER_24_652 ();
 sg13g2_decap_8 FILLER_24_659 ();
 sg13g2_decap_8 FILLER_24_666 ();
 sg13g2_decap_8 FILLER_24_673 ();
 sg13g2_decap_8 FILLER_24_680 ();
 sg13g2_decap_8 FILLER_24_687 ();
 sg13g2_decap_8 FILLER_24_694 ();
 sg13g2_decap_8 FILLER_24_701 ();
 sg13g2_decap_8 FILLER_24_708 ();
 sg13g2_decap_8 FILLER_24_715 ();
 sg13g2_decap_8 FILLER_24_722 ();
 sg13g2_decap_8 FILLER_24_729 ();
 sg13g2_decap_8 FILLER_24_736 ();
 sg13g2_decap_8 FILLER_24_743 ();
 sg13g2_decap_8 FILLER_24_750 ();
 sg13g2_decap_8 FILLER_24_757 ();
 sg13g2_decap_8 FILLER_24_764 ();
 sg13g2_decap_8 FILLER_24_771 ();
 sg13g2_decap_8 FILLER_24_778 ();
 sg13g2_decap_8 FILLER_24_785 ();
 sg13g2_decap_8 FILLER_24_792 ();
 sg13g2_decap_8 FILLER_24_799 ();
 sg13g2_decap_8 FILLER_24_806 ();
 sg13g2_decap_8 FILLER_24_813 ();
 sg13g2_decap_8 FILLER_24_820 ();
 sg13g2_decap_8 FILLER_24_827 ();
 sg13g2_decap_8 FILLER_24_834 ();
 sg13g2_decap_8 FILLER_24_841 ();
 sg13g2_decap_8 FILLER_24_848 ();
 sg13g2_decap_8 FILLER_24_855 ();
 sg13g2_decap_8 FILLER_24_862 ();
 sg13g2_decap_8 FILLER_24_869 ();
 sg13g2_decap_8 FILLER_24_876 ();
 sg13g2_decap_8 FILLER_24_883 ();
 sg13g2_decap_8 FILLER_24_890 ();
 sg13g2_decap_8 FILLER_24_897 ();
 sg13g2_decap_8 FILLER_24_904 ();
 sg13g2_decap_8 FILLER_24_911 ();
 sg13g2_decap_8 FILLER_24_918 ();
 sg13g2_decap_8 FILLER_24_925 ();
 sg13g2_decap_8 FILLER_24_932 ();
 sg13g2_decap_8 FILLER_24_939 ();
 sg13g2_decap_8 FILLER_24_946 ();
 sg13g2_decap_8 FILLER_24_953 ();
 sg13g2_decap_8 FILLER_24_960 ();
 sg13g2_decap_8 FILLER_24_967 ();
 sg13g2_decap_8 FILLER_24_974 ();
 sg13g2_decap_8 FILLER_24_981 ();
 sg13g2_decap_8 FILLER_24_988 ();
 sg13g2_decap_8 FILLER_24_995 ();
 sg13g2_decap_8 FILLER_24_1002 ();
 sg13g2_decap_8 FILLER_24_1009 ();
 sg13g2_decap_8 FILLER_24_1016 ();
 sg13g2_decap_4 FILLER_24_1023 ();
 sg13g2_fill_2 FILLER_24_1027 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_1 FILLER_25_23 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_fill_2 FILLER_25_88 ();
 sg13g2_fill_2 FILLER_25_120 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_fill_1 FILLER_25_153 ();
 sg13g2_fill_2 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_179 ();
 sg13g2_fill_2 FILLER_25_205 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_2 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_fill_1 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_decap_8 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_decap_8 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_25_436 ();
 sg13g2_decap_8 FILLER_25_443 ();
 sg13g2_decap_8 FILLER_25_450 ();
 sg13g2_decap_8 FILLER_25_457 ();
 sg13g2_decap_8 FILLER_25_464 ();
 sg13g2_decap_8 FILLER_25_471 ();
 sg13g2_decap_8 FILLER_25_478 ();
 sg13g2_decap_8 FILLER_25_485 ();
 sg13g2_decap_8 FILLER_25_492 ();
 sg13g2_decap_8 FILLER_25_499 ();
 sg13g2_decap_8 FILLER_25_506 ();
 sg13g2_decap_8 FILLER_25_513 ();
 sg13g2_decap_8 FILLER_25_520 ();
 sg13g2_decap_8 FILLER_25_527 ();
 sg13g2_decap_8 FILLER_25_534 ();
 sg13g2_decap_8 FILLER_25_541 ();
 sg13g2_decap_8 FILLER_25_548 ();
 sg13g2_decap_8 FILLER_25_555 ();
 sg13g2_decap_8 FILLER_25_562 ();
 sg13g2_decap_8 FILLER_25_569 ();
 sg13g2_decap_8 FILLER_25_576 ();
 sg13g2_decap_8 FILLER_25_583 ();
 sg13g2_decap_8 FILLER_25_590 ();
 sg13g2_decap_8 FILLER_25_597 ();
 sg13g2_decap_8 FILLER_25_604 ();
 sg13g2_decap_8 FILLER_25_611 ();
 sg13g2_decap_8 FILLER_25_618 ();
 sg13g2_decap_8 FILLER_25_625 ();
 sg13g2_decap_8 FILLER_25_632 ();
 sg13g2_decap_8 FILLER_25_639 ();
 sg13g2_decap_8 FILLER_25_646 ();
 sg13g2_decap_8 FILLER_25_653 ();
 sg13g2_decap_8 FILLER_25_660 ();
 sg13g2_decap_8 FILLER_25_667 ();
 sg13g2_decap_8 FILLER_25_674 ();
 sg13g2_decap_8 FILLER_25_681 ();
 sg13g2_decap_8 FILLER_25_688 ();
 sg13g2_decap_8 FILLER_25_695 ();
 sg13g2_decap_8 FILLER_25_702 ();
 sg13g2_decap_8 FILLER_25_709 ();
 sg13g2_decap_8 FILLER_25_716 ();
 sg13g2_decap_8 FILLER_25_723 ();
 sg13g2_decap_8 FILLER_25_730 ();
 sg13g2_decap_8 FILLER_25_737 ();
 sg13g2_decap_8 FILLER_25_744 ();
 sg13g2_decap_8 FILLER_25_751 ();
 sg13g2_decap_8 FILLER_25_758 ();
 sg13g2_decap_8 FILLER_25_765 ();
 sg13g2_decap_8 FILLER_25_772 ();
 sg13g2_decap_8 FILLER_25_779 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_8 FILLER_25_856 ();
 sg13g2_decap_8 FILLER_25_863 ();
 sg13g2_decap_8 FILLER_25_870 ();
 sg13g2_decap_8 FILLER_25_877 ();
 sg13g2_decap_8 FILLER_25_884 ();
 sg13g2_decap_8 FILLER_25_891 ();
 sg13g2_decap_8 FILLER_25_898 ();
 sg13g2_decap_8 FILLER_25_905 ();
 sg13g2_decap_8 FILLER_25_912 ();
 sg13g2_decap_8 FILLER_25_919 ();
 sg13g2_decap_8 FILLER_25_926 ();
 sg13g2_decap_8 FILLER_25_933 ();
 sg13g2_decap_8 FILLER_25_940 ();
 sg13g2_decap_8 FILLER_25_947 ();
 sg13g2_decap_8 FILLER_25_954 ();
 sg13g2_decap_8 FILLER_25_961 ();
 sg13g2_decap_8 FILLER_25_968 ();
 sg13g2_decap_8 FILLER_25_975 ();
 sg13g2_decap_8 FILLER_25_982 ();
 sg13g2_decap_8 FILLER_25_989 ();
 sg13g2_decap_8 FILLER_25_996 ();
 sg13g2_decap_8 FILLER_25_1003 ();
 sg13g2_decap_8 FILLER_25_1010 ();
 sg13g2_decap_8 FILLER_25_1017 ();
 sg13g2_decap_4 FILLER_25_1024 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_29 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_2 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_2 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_decap_8 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_422 ();
 sg13g2_decap_8 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_26_436 ();
 sg13g2_decap_8 FILLER_26_443 ();
 sg13g2_decap_8 FILLER_26_450 ();
 sg13g2_decap_8 FILLER_26_457 ();
 sg13g2_decap_8 FILLER_26_464 ();
 sg13g2_decap_8 FILLER_26_471 ();
 sg13g2_decap_8 FILLER_26_478 ();
 sg13g2_decap_8 FILLER_26_485 ();
 sg13g2_decap_8 FILLER_26_492 ();
 sg13g2_decap_8 FILLER_26_499 ();
 sg13g2_decap_8 FILLER_26_506 ();
 sg13g2_decap_8 FILLER_26_513 ();
 sg13g2_decap_8 FILLER_26_520 ();
 sg13g2_decap_8 FILLER_26_527 ();
 sg13g2_decap_8 FILLER_26_534 ();
 sg13g2_decap_8 FILLER_26_541 ();
 sg13g2_decap_8 FILLER_26_548 ();
 sg13g2_decap_8 FILLER_26_555 ();
 sg13g2_decap_8 FILLER_26_562 ();
 sg13g2_decap_8 FILLER_26_569 ();
 sg13g2_decap_8 FILLER_26_576 ();
 sg13g2_decap_8 FILLER_26_583 ();
 sg13g2_decap_8 FILLER_26_590 ();
 sg13g2_decap_8 FILLER_26_597 ();
 sg13g2_decap_8 FILLER_26_604 ();
 sg13g2_decap_8 FILLER_26_611 ();
 sg13g2_decap_8 FILLER_26_618 ();
 sg13g2_decap_8 FILLER_26_625 ();
 sg13g2_decap_8 FILLER_26_632 ();
 sg13g2_decap_8 FILLER_26_639 ();
 sg13g2_decap_8 FILLER_26_646 ();
 sg13g2_decap_8 FILLER_26_653 ();
 sg13g2_decap_8 FILLER_26_660 ();
 sg13g2_decap_8 FILLER_26_667 ();
 sg13g2_decap_8 FILLER_26_674 ();
 sg13g2_decap_8 FILLER_26_681 ();
 sg13g2_decap_8 FILLER_26_688 ();
 sg13g2_decap_8 FILLER_26_695 ();
 sg13g2_decap_8 FILLER_26_702 ();
 sg13g2_decap_8 FILLER_26_709 ();
 sg13g2_decap_8 FILLER_26_716 ();
 sg13g2_decap_8 FILLER_26_723 ();
 sg13g2_decap_8 FILLER_26_730 ();
 sg13g2_decap_8 FILLER_26_737 ();
 sg13g2_decap_8 FILLER_26_744 ();
 sg13g2_decap_8 FILLER_26_751 ();
 sg13g2_decap_8 FILLER_26_758 ();
 sg13g2_decap_8 FILLER_26_765 ();
 sg13g2_decap_8 FILLER_26_772 ();
 sg13g2_decap_8 FILLER_26_779 ();
 sg13g2_decap_8 FILLER_26_786 ();
 sg13g2_decap_8 FILLER_26_793 ();
 sg13g2_decap_8 FILLER_26_800 ();
 sg13g2_decap_8 FILLER_26_807 ();
 sg13g2_decap_8 FILLER_26_814 ();
 sg13g2_decap_8 FILLER_26_821 ();
 sg13g2_decap_8 FILLER_26_828 ();
 sg13g2_decap_8 FILLER_26_835 ();
 sg13g2_decap_8 FILLER_26_842 ();
 sg13g2_decap_8 FILLER_26_849 ();
 sg13g2_decap_8 FILLER_26_856 ();
 sg13g2_decap_8 FILLER_26_863 ();
 sg13g2_decap_8 FILLER_26_870 ();
 sg13g2_decap_8 FILLER_26_877 ();
 sg13g2_decap_8 FILLER_26_884 ();
 sg13g2_decap_8 FILLER_26_891 ();
 sg13g2_decap_8 FILLER_26_898 ();
 sg13g2_decap_8 FILLER_26_905 ();
 sg13g2_decap_8 FILLER_26_912 ();
 sg13g2_decap_8 FILLER_26_919 ();
 sg13g2_decap_8 FILLER_26_926 ();
 sg13g2_decap_8 FILLER_26_933 ();
 sg13g2_decap_8 FILLER_26_940 ();
 sg13g2_decap_8 FILLER_26_947 ();
 sg13g2_decap_8 FILLER_26_954 ();
 sg13g2_decap_8 FILLER_26_961 ();
 sg13g2_decap_8 FILLER_26_968 ();
 sg13g2_decap_8 FILLER_26_975 ();
 sg13g2_decap_8 FILLER_26_982 ();
 sg13g2_decap_8 FILLER_26_989 ();
 sg13g2_decap_8 FILLER_26_996 ();
 sg13g2_decap_8 FILLER_26_1003 ();
 sg13g2_decap_8 FILLER_26_1010 ();
 sg13g2_decap_8 FILLER_26_1017 ();
 sg13g2_decap_4 FILLER_26_1024 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_fill_2 FILLER_27_22 ();
 sg13g2_fill_1 FILLER_27_48 ();
 sg13g2_fill_2 FILLER_27_59 ();
 sg13g2_fill_2 FILLER_27_79 ();
 sg13g2_fill_1 FILLER_27_81 ();
 sg13g2_fill_2 FILLER_27_121 ();
 sg13g2_fill_1 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_fill_2 FILLER_27_192 ();
 sg13g2_fill_2 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_decap_4 FILLER_27_401 ();
 sg13g2_fill_2 FILLER_27_419 ();
 sg13g2_fill_1 FILLER_27_421 ();
 sg13g2_decap_8 FILLER_27_431 ();
 sg13g2_decap_8 FILLER_27_438 ();
 sg13g2_decap_8 FILLER_27_445 ();
 sg13g2_decap_8 FILLER_27_452 ();
 sg13g2_decap_8 FILLER_27_459 ();
 sg13g2_decap_8 FILLER_27_466 ();
 sg13g2_decap_8 FILLER_27_473 ();
 sg13g2_decap_8 FILLER_27_480 ();
 sg13g2_decap_8 FILLER_27_487 ();
 sg13g2_decap_8 FILLER_27_494 ();
 sg13g2_decap_8 FILLER_27_501 ();
 sg13g2_decap_8 FILLER_27_508 ();
 sg13g2_decap_8 FILLER_27_515 ();
 sg13g2_decap_8 FILLER_27_522 ();
 sg13g2_decap_8 FILLER_27_529 ();
 sg13g2_decap_8 FILLER_27_536 ();
 sg13g2_decap_8 FILLER_27_543 ();
 sg13g2_decap_8 FILLER_27_550 ();
 sg13g2_decap_8 FILLER_27_557 ();
 sg13g2_decap_8 FILLER_27_564 ();
 sg13g2_decap_8 FILLER_27_571 ();
 sg13g2_decap_8 FILLER_27_578 ();
 sg13g2_decap_8 FILLER_27_585 ();
 sg13g2_decap_8 FILLER_27_592 ();
 sg13g2_decap_8 FILLER_27_599 ();
 sg13g2_decap_8 FILLER_27_606 ();
 sg13g2_decap_8 FILLER_27_613 ();
 sg13g2_decap_8 FILLER_27_620 ();
 sg13g2_decap_8 FILLER_27_627 ();
 sg13g2_decap_8 FILLER_27_634 ();
 sg13g2_decap_8 FILLER_27_641 ();
 sg13g2_decap_8 FILLER_27_648 ();
 sg13g2_decap_8 FILLER_27_655 ();
 sg13g2_decap_8 FILLER_27_662 ();
 sg13g2_decap_8 FILLER_27_669 ();
 sg13g2_decap_8 FILLER_27_676 ();
 sg13g2_decap_8 FILLER_27_683 ();
 sg13g2_decap_8 FILLER_27_690 ();
 sg13g2_decap_8 FILLER_27_697 ();
 sg13g2_decap_8 FILLER_27_704 ();
 sg13g2_decap_8 FILLER_27_711 ();
 sg13g2_decap_8 FILLER_27_718 ();
 sg13g2_decap_8 FILLER_27_725 ();
 sg13g2_decap_8 FILLER_27_732 ();
 sg13g2_decap_8 FILLER_27_739 ();
 sg13g2_decap_8 FILLER_27_746 ();
 sg13g2_decap_8 FILLER_27_753 ();
 sg13g2_decap_8 FILLER_27_760 ();
 sg13g2_decap_8 FILLER_27_767 ();
 sg13g2_decap_8 FILLER_27_774 ();
 sg13g2_decap_8 FILLER_27_781 ();
 sg13g2_decap_8 FILLER_27_788 ();
 sg13g2_decap_8 FILLER_27_795 ();
 sg13g2_decap_8 FILLER_27_802 ();
 sg13g2_decap_8 FILLER_27_809 ();
 sg13g2_decap_8 FILLER_27_816 ();
 sg13g2_decap_8 FILLER_27_823 ();
 sg13g2_decap_8 FILLER_27_830 ();
 sg13g2_decap_8 FILLER_27_837 ();
 sg13g2_decap_8 FILLER_27_844 ();
 sg13g2_decap_8 FILLER_27_851 ();
 sg13g2_decap_8 FILLER_27_858 ();
 sg13g2_decap_8 FILLER_27_865 ();
 sg13g2_decap_8 FILLER_27_872 ();
 sg13g2_decap_8 FILLER_27_879 ();
 sg13g2_decap_8 FILLER_27_886 ();
 sg13g2_decap_8 FILLER_27_893 ();
 sg13g2_decap_8 FILLER_27_900 ();
 sg13g2_decap_8 FILLER_27_907 ();
 sg13g2_decap_8 FILLER_27_914 ();
 sg13g2_decap_8 FILLER_27_921 ();
 sg13g2_decap_8 FILLER_27_928 ();
 sg13g2_decap_8 FILLER_27_935 ();
 sg13g2_decap_8 FILLER_27_942 ();
 sg13g2_decap_8 FILLER_27_949 ();
 sg13g2_decap_8 FILLER_27_956 ();
 sg13g2_decap_8 FILLER_27_963 ();
 sg13g2_decap_8 FILLER_27_970 ();
 sg13g2_decap_8 FILLER_27_977 ();
 sg13g2_decap_8 FILLER_27_984 ();
 sg13g2_decap_8 FILLER_27_991 ();
 sg13g2_decap_8 FILLER_27_998 ();
 sg13g2_decap_8 FILLER_27_1005 ();
 sg13g2_decap_8 FILLER_27_1012 ();
 sg13g2_decap_8 FILLER_27_1019 ();
 sg13g2_fill_2 FILLER_27_1026 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_fill_1 FILLER_28_164 ();
 sg13g2_fill_2 FILLER_28_199 ();
 sg13g2_fill_1 FILLER_28_229 ();
 sg13g2_decap_4 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_375 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_decap_8 FILLER_28_435 ();
 sg13g2_decap_8 FILLER_28_442 ();
 sg13g2_decap_8 FILLER_28_449 ();
 sg13g2_decap_8 FILLER_28_456 ();
 sg13g2_decap_8 FILLER_28_463 ();
 sg13g2_decap_8 FILLER_28_470 ();
 sg13g2_decap_8 FILLER_28_477 ();
 sg13g2_decap_8 FILLER_28_484 ();
 sg13g2_decap_8 FILLER_28_491 ();
 sg13g2_decap_8 FILLER_28_498 ();
 sg13g2_decap_8 FILLER_28_505 ();
 sg13g2_decap_8 FILLER_28_512 ();
 sg13g2_decap_8 FILLER_28_519 ();
 sg13g2_decap_8 FILLER_28_526 ();
 sg13g2_decap_8 FILLER_28_533 ();
 sg13g2_decap_8 FILLER_28_540 ();
 sg13g2_decap_8 FILLER_28_547 ();
 sg13g2_decap_8 FILLER_28_554 ();
 sg13g2_decap_8 FILLER_28_561 ();
 sg13g2_decap_8 FILLER_28_568 ();
 sg13g2_decap_8 FILLER_28_575 ();
 sg13g2_decap_8 FILLER_28_582 ();
 sg13g2_decap_8 FILLER_28_589 ();
 sg13g2_decap_8 FILLER_28_596 ();
 sg13g2_decap_8 FILLER_28_603 ();
 sg13g2_decap_8 FILLER_28_610 ();
 sg13g2_decap_8 FILLER_28_617 ();
 sg13g2_decap_8 FILLER_28_624 ();
 sg13g2_decap_8 FILLER_28_631 ();
 sg13g2_decap_8 FILLER_28_638 ();
 sg13g2_decap_8 FILLER_28_645 ();
 sg13g2_decap_8 FILLER_28_652 ();
 sg13g2_decap_8 FILLER_28_659 ();
 sg13g2_decap_8 FILLER_28_666 ();
 sg13g2_decap_8 FILLER_28_673 ();
 sg13g2_decap_8 FILLER_28_680 ();
 sg13g2_decap_8 FILLER_28_687 ();
 sg13g2_decap_8 FILLER_28_694 ();
 sg13g2_decap_8 FILLER_28_701 ();
 sg13g2_decap_8 FILLER_28_708 ();
 sg13g2_decap_8 FILLER_28_715 ();
 sg13g2_decap_8 FILLER_28_722 ();
 sg13g2_decap_8 FILLER_28_729 ();
 sg13g2_decap_8 FILLER_28_736 ();
 sg13g2_decap_8 FILLER_28_743 ();
 sg13g2_decap_8 FILLER_28_750 ();
 sg13g2_decap_8 FILLER_28_757 ();
 sg13g2_decap_8 FILLER_28_764 ();
 sg13g2_decap_8 FILLER_28_771 ();
 sg13g2_decap_8 FILLER_28_778 ();
 sg13g2_decap_8 FILLER_28_785 ();
 sg13g2_decap_8 FILLER_28_792 ();
 sg13g2_decap_8 FILLER_28_799 ();
 sg13g2_decap_8 FILLER_28_806 ();
 sg13g2_decap_8 FILLER_28_813 ();
 sg13g2_decap_8 FILLER_28_820 ();
 sg13g2_decap_8 FILLER_28_827 ();
 sg13g2_decap_8 FILLER_28_834 ();
 sg13g2_decap_8 FILLER_28_841 ();
 sg13g2_decap_8 FILLER_28_848 ();
 sg13g2_decap_8 FILLER_28_855 ();
 sg13g2_decap_8 FILLER_28_862 ();
 sg13g2_decap_8 FILLER_28_869 ();
 sg13g2_decap_8 FILLER_28_876 ();
 sg13g2_decap_8 FILLER_28_883 ();
 sg13g2_decap_8 FILLER_28_890 ();
 sg13g2_decap_8 FILLER_28_897 ();
 sg13g2_decap_8 FILLER_28_904 ();
 sg13g2_decap_8 FILLER_28_911 ();
 sg13g2_decap_8 FILLER_28_918 ();
 sg13g2_decap_8 FILLER_28_925 ();
 sg13g2_decap_8 FILLER_28_932 ();
 sg13g2_decap_8 FILLER_28_939 ();
 sg13g2_decap_8 FILLER_28_946 ();
 sg13g2_decap_8 FILLER_28_953 ();
 sg13g2_decap_8 FILLER_28_960 ();
 sg13g2_decap_8 FILLER_28_967 ();
 sg13g2_decap_8 FILLER_28_974 ();
 sg13g2_decap_8 FILLER_28_981 ();
 sg13g2_decap_8 FILLER_28_988 ();
 sg13g2_decap_8 FILLER_28_995 ();
 sg13g2_decap_8 FILLER_28_1002 ();
 sg13g2_decap_8 FILLER_28_1009 ();
 sg13g2_decap_8 FILLER_28_1016 ();
 sg13g2_decap_4 FILLER_28_1023 ();
 sg13g2_fill_2 FILLER_28_1027 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_53 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_fill_1 FILLER_29_100 ();
 sg13g2_fill_2 FILLER_29_128 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_fill_2 FILLER_29_355 ();
 sg13g2_decap_4 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_29_403 ();
 sg13g2_fill_1 FILLER_29_410 ();
 sg13g2_decap_8 FILLER_29_447 ();
 sg13g2_decap_8 FILLER_29_454 ();
 sg13g2_decap_8 FILLER_29_461 ();
 sg13g2_decap_8 FILLER_29_468 ();
 sg13g2_decap_8 FILLER_29_475 ();
 sg13g2_decap_8 FILLER_29_482 ();
 sg13g2_decap_8 FILLER_29_489 ();
 sg13g2_decap_8 FILLER_29_496 ();
 sg13g2_decap_8 FILLER_29_503 ();
 sg13g2_decap_8 FILLER_29_510 ();
 sg13g2_decap_8 FILLER_29_517 ();
 sg13g2_decap_8 FILLER_29_524 ();
 sg13g2_decap_8 FILLER_29_531 ();
 sg13g2_decap_8 FILLER_29_538 ();
 sg13g2_decap_8 FILLER_29_545 ();
 sg13g2_decap_8 FILLER_29_552 ();
 sg13g2_decap_8 FILLER_29_559 ();
 sg13g2_decap_8 FILLER_29_566 ();
 sg13g2_decap_8 FILLER_29_573 ();
 sg13g2_decap_8 FILLER_29_580 ();
 sg13g2_decap_8 FILLER_29_587 ();
 sg13g2_decap_8 FILLER_29_594 ();
 sg13g2_decap_8 FILLER_29_601 ();
 sg13g2_decap_8 FILLER_29_608 ();
 sg13g2_decap_8 FILLER_29_615 ();
 sg13g2_decap_8 FILLER_29_622 ();
 sg13g2_decap_8 FILLER_29_629 ();
 sg13g2_decap_8 FILLER_29_636 ();
 sg13g2_decap_8 FILLER_29_643 ();
 sg13g2_decap_8 FILLER_29_650 ();
 sg13g2_decap_8 FILLER_29_657 ();
 sg13g2_decap_8 FILLER_29_664 ();
 sg13g2_decap_8 FILLER_29_671 ();
 sg13g2_decap_8 FILLER_29_678 ();
 sg13g2_decap_8 FILLER_29_685 ();
 sg13g2_decap_8 FILLER_29_692 ();
 sg13g2_decap_8 FILLER_29_699 ();
 sg13g2_decap_8 FILLER_29_706 ();
 sg13g2_decap_8 FILLER_29_713 ();
 sg13g2_decap_8 FILLER_29_720 ();
 sg13g2_decap_8 FILLER_29_727 ();
 sg13g2_decap_8 FILLER_29_734 ();
 sg13g2_decap_8 FILLER_29_741 ();
 sg13g2_decap_8 FILLER_29_748 ();
 sg13g2_decap_8 FILLER_29_755 ();
 sg13g2_decap_8 FILLER_29_762 ();
 sg13g2_decap_8 FILLER_29_769 ();
 sg13g2_decap_8 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_783 ();
 sg13g2_decap_8 FILLER_29_790 ();
 sg13g2_decap_8 FILLER_29_797 ();
 sg13g2_decap_8 FILLER_29_804 ();
 sg13g2_decap_8 FILLER_29_811 ();
 sg13g2_decap_8 FILLER_29_818 ();
 sg13g2_decap_8 FILLER_29_825 ();
 sg13g2_decap_8 FILLER_29_832 ();
 sg13g2_decap_8 FILLER_29_839 ();
 sg13g2_decap_8 FILLER_29_846 ();
 sg13g2_decap_8 FILLER_29_853 ();
 sg13g2_decap_8 FILLER_29_860 ();
 sg13g2_decap_8 FILLER_29_867 ();
 sg13g2_decap_8 FILLER_29_874 ();
 sg13g2_decap_8 FILLER_29_881 ();
 sg13g2_decap_8 FILLER_29_888 ();
 sg13g2_decap_8 FILLER_29_895 ();
 sg13g2_decap_8 FILLER_29_902 ();
 sg13g2_decap_8 FILLER_29_909 ();
 sg13g2_decap_8 FILLER_29_916 ();
 sg13g2_decap_8 FILLER_29_923 ();
 sg13g2_decap_8 FILLER_29_930 ();
 sg13g2_decap_8 FILLER_29_937 ();
 sg13g2_decap_8 FILLER_29_944 ();
 sg13g2_decap_8 FILLER_29_951 ();
 sg13g2_decap_8 FILLER_29_958 ();
 sg13g2_decap_8 FILLER_29_965 ();
 sg13g2_decap_8 FILLER_29_972 ();
 sg13g2_decap_8 FILLER_29_979 ();
 sg13g2_decap_8 FILLER_29_986 ();
 sg13g2_decap_8 FILLER_29_993 ();
 sg13g2_decap_8 FILLER_29_1000 ();
 sg13g2_decap_8 FILLER_29_1007 ();
 sg13g2_decap_8 FILLER_29_1014 ();
 sg13g2_decap_8 FILLER_29_1021 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_40 ();
 sg13g2_fill_1 FILLER_30_95 ();
 sg13g2_fill_2 FILLER_30_128 ();
 sg13g2_fill_1 FILLER_30_130 ();
 sg13g2_fill_2 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_fill_2 FILLER_30_372 ();
 sg13g2_decap_4 FILLER_30_377 ();
 sg13g2_decap_4 FILLER_30_409 ();
 sg13g2_fill_1 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_444 ();
 sg13g2_fill_1 FILLER_30_451 ();
 sg13g2_decap_8 FILLER_30_465 ();
 sg13g2_decap_8 FILLER_30_472 ();
 sg13g2_decap_8 FILLER_30_479 ();
 sg13g2_decap_8 FILLER_30_486 ();
 sg13g2_decap_8 FILLER_30_493 ();
 sg13g2_decap_8 FILLER_30_500 ();
 sg13g2_decap_8 FILLER_30_507 ();
 sg13g2_decap_8 FILLER_30_514 ();
 sg13g2_decap_8 FILLER_30_521 ();
 sg13g2_decap_8 FILLER_30_528 ();
 sg13g2_decap_8 FILLER_30_535 ();
 sg13g2_decap_8 FILLER_30_542 ();
 sg13g2_decap_8 FILLER_30_549 ();
 sg13g2_decap_8 FILLER_30_556 ();
 sg13g2_decap_8 FILLER_30_563 ();
 sg13g2_decap_8 FILLER_30_570 ();
 sg13g2_decap_8 FILLER_30_577 ();
 sg13g2_decap_8 FILLER_30_584 ();
 sg13g2_decap_8 FILLER_30_591 ();
 sg13g2_decap_8 FILLER_30_598 ();
 sg13g2_decap_8 FILLER_30_605 ();
 sg13g2_decap_8 FILLER_30_612 ();
 sg13g2_decap_8 FILLER_30_619 ();
 sg13g2_decap_8 FILLER_30_626 ();
 sg13g2_decap_8 FILLER_30_633 ();
 sg13g2_decap_8 FILLER_30_640 ();
 sg13g2_decap_8 FILLER_30_647 ();
 sg13g2_decap_8 FILLER_30_654 ();
 sg13g2_decap_8 FILLER_30_661 ();
 sg13g2_decap_8 FILLER_30_668 ();
 sg13g2_decap_8 FILLER_30_675 ();
 sg13g2_decap_8 FILLER_30_682 ();
 sg13g2_decap_8 FILLER_30_689 ();
 sg13g2_decap_8 FILLER_30_696 ();
 sg13g2_decap_8 FILLER_30_703 ();
 sg13g2_decap_8 FILLER_30_710 ();
 sg13g2_decap_8 FILLER_30_717 ();
 sg13g2_decap_8 FILLER_30_724 ();
 sg13g2_decap_8 FILLER_30_731 ();
 sg13g2_decap_8 FILLER_30_738 ();
 sg13g2_decap_8 FILLER_30_745 ();
 sg13g2_decap_8 FILLER_30_752 ();
 sg13g2_decap_8 FILLER_30_759 ();
 sg13g2_decap_8 FILLER_30_766 ();
 sg13g2_decap_8 FILLER_30_773 ();
 sg13g2_decap_8 FILLER_30_780 ();
 sg13g2_decap_8 FILLER_30_787 ();
 sg13g2_decap_8 FILLER_30_794 ();
 sg13g2_decap_8 FILLER_30_801 ();
 sg13g2_decap_8 FILLER_30_808 ();
 sg13g2_decap_8 FILLER_30_815 ();
 sg13g2_decap_8 FILLER_30_822 ();
 sg13g2_decap_8 FILLER_30_829 ();
 sg13g2_decap_8 FILLER_30_836 ();
 sg13g2_decap_8 FILLER_30_843 ();
 sg13g2_decap_8 FILLER_30_850 ();
 sg13g2_decap_8 FILLER_30_857 ();
 sg13g2_decap_8 FILLER_30_864 ();
 sg13g2_decap_8 FILLER_30_871 ();
 sg13g2_decap_8 FILLER_30_878 ();
 sg13g2_decap_8 FILLER_30_885 ();
 sg13g2_decap_8 FILLER_30_892 ();
 sg13g2_decap_8 FILLER_30_899 ();
 sg13g2_decap_8 FILLER_30_906 ();
 sg13g2_decap_8 FILLER_30_913 ();
 sg13g2_decap_8 FILLER_30_920 ();
 sg13g2_decap_8 FILLER_30_927 ();
 sg13g2_decap_8 FILLER_30_934 ();
 sg13g2_decap_8 FILLER_30_941 ();
 sg13g2_decap_8 FILLER_30_948 ();
 sg13g2_decap_8 FILLER_30_955 ();
 sg13g2_decap_8 FILLER_30_962 ();
 sg13g2_decap_8 FILLER_30_969 ();
 sg13g2_decap_8 FILLER_30_976 ();
 sg13g2_decap_8 FILLER_30_983 ();
 sg13g2_decap_8 FILLER_30_990 ();
 sg13g2_decap_8 FILLER_30_997 ();
 sg13g2_decap_8 FILLER_30_1004 ();
 sg13g2_decap_8 FILLER_30_1011 ();
 sg13g2_decap_8 FILLER_30_1018 ();
 sg13g2_decap_4 FILLER_30_1025 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_48 ();
 sg13g2_fill_2 FILLER_31_76 ();
 sg13g2_fill_1 FILLER_31_91 ();
 sg13g2_fill_2 FILLER_31_106 ();
 sg13g2_fill_2 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_115 ();
 sg13g2_fill_1 FILLER_31_125 ();
 sg13g2_fill_2 FILLER_31_155 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_fill_2 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_256 ();
 sg13g2_fill_1 FILLER_31_258 ();
 sg13g2_fill_1 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_386 ();
 sg13g2_fill_2 FILLER_31_413 ();
 sg13g2_fill_2 FILLER_31_442 ();
 sg13g2_decap_8 FILLER_31_484 ();
 sg13g2_decap_8 FILLER_31_491 ();
 sg13g2_decap_8 FILLER_31_498 ();
 sg13g2_decap_8 FILLER_31_505 ();
 sg13g2_decap_8 FILLER_31_512 ();
 sg13g2_decap_8 FILLER_31_519 ();
 sg13g2_decap_8 FILLER_31_526 ();
 sg13g2_decap_8 FILLER_31_533 ();
 sg13g2_decap_8 FILLER_31_540 ();
 sg13g2_decap_8 FILLER_31_547 ();
 sg13g2_decap_8 FILLER_31_554 ();
 sg13g2_decap_8 FILLER_31_561 ();
 sg13g2_decap_8 FILLER_31_568 ();
 sg13g2_decap_8 FILLER_31_575 ();
 sg13g2_decap_8 FILLER_31_582 ();
 sg13g2_decap_8 FILLER_31_589 ();
 sg13g2_decap_8 FILLER_31_596 ();
 sg13g2_decap_8 FILLER_31_603 ();
 sg13g2_decap_8 FILLER_31_610 ();
 sg13g2_decap_8 FILLER_31_617 ();
 sg13g2_decap_8 FILLER_31_624 ();
 sg13g2_decap_8 FILLER_31_631 ();
 sg13g2_decap_8 FILLER_31_638 ();
 sg13g2_decap_8 FILLER_31_645 ();
 sg13g2_decap_8 FILLER_31_652 ();
 sg13g2_decap_8 FILLER_31_659 ();
 sg13g2_decap_8 FILLER_31_666 ();
 sg13g2_decap_8 FILLER_31_673 ();
 sg13g2_decap_8 FILLER_31_680 ();
 sg13g2_decap_8 FILLER_31_687 ();
 sg13g2_decap_8 FILLER_31_694 ();
 sg13g2_decap_8 FILLER_31_701 ();
 sg13g2_decap_8 FILLER_31_708 ();
 sg13g2_decap_8 FILLER_31_715 ();
 sg13g2_decap_8 FILLER_31_722 ();
 sg13g2_decap_8 FILLER_31_729 ();
 sg13g2_decap_8 FILLER_31_736 ();
 sg13g2_decap_8 FILLER_31_743 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_decap_8 FILLER_31_757 ();
 sg13g2_decap_8 FILLER_31_764 ();
 sg13g2_decap_8 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_778 ();
 sg13g2_decap_8 FILLER_31_785 ();
 sg13g2_decap_8 FILLER_31_792 ();
 sg13g2_decap_8 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_806 ();
 sg13g2_decap_8 FILLER_31_813 ();
 sg13g2_decap_8 FILLER_31_820 ();
 sg13g2_decap_8 FILLER_31_827 ();
 sg13g2_decap_8 FILLER_31_834 ();
 sg13g2_decap_8 FILLER_31_841 ();
 sg13g2_decap_8 FILLER_31_848 ();
 sg13g2_decap_8 FILLER_31_855 ();
 sg13g2_decap_8 FILLER_31_862 ();
 sg13g2_decap_8 FILLER_31_869 ();
 sg13g2_decap_8 FILLER_31_876 ();
 sg13g2_decap_8 FILLER_31_883 ();
 sg13g2_decap_8 FILLER_31_890 ();
 sg13g2_decap_8 FILLER_31_897 ();
 sg13g2_decap_8 FILLER_31_904 ();
 sg13g2_decap_8 FILLER_31_911 ();
 sg13g2_decap_8 FILLER_31_918 ();
 sg13g2_decap_8 FILLER_31_925 ();
 sg13g2_decap_8 FILLER_31_932 ();
 sg13g2_decap_8 FILLER_31_939 ();
 sg13g2_decap_8 FILLER_31_946 ();
 sg13g2_decap_8 FILLER_31_953 ();
 sg13g2_decap_8 FILLER_31_960 ();
 sg13g2_decap_8 FILLER_31_967 ();
 sg13g2_decap_8 FILLER_31_974 ();
 sg13g2_decap_8 FILLER_31_981 ();
 sg13g2_decap_8 FILLER_31_988 ();
 sg13g2_decap_8 FILLER_31_995 ();
 sg13g2_decap_8 FILLER_31_1002 ();
 sg13g2_decap_8 FILLER_31_1009 ();
 sg13g2_decap_8 FILLER_31_1016 ();
 sg13g2_decap_4 FILLER_31_1023 ();
 sg13g2_fill_2 FILLER_31_1027 ();
 sg13g2_fill_1 FILLER_32_27 ();
 sg13g2_fill_1 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_155 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_357 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_fill_2 FILLER_32_461 ();
 sg13g2_decap_8 FILLER_32_490 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_504 ();
 sg13g2_decap_8 FILLER_32_511 ();
 sg13g2_decap_8 FILLER_32_518 ();
 sg13g2_decap_8 FILLER_32_525 ();
 sg13g2_decap_8 FILLER_32_532 ();
 sg13g2_decap_8 FILLER_32_539 ();
 sg13g2_decap_8 FILLER_32_546 ();
 sg13g2_decap_8 FILLER_32_553 ();
 sg13g2_decap_8 FILLER_32_560 ();
 sg13g2_decap_8 FILLER_32_567 ();
 sg13g2_decap_8 FILLER_32_574 ();
 sg13g2_decap_8 FILLER_32_581 ();
 sg13g2_decap_8 FILLER_32_588 ();
 sg13g2_decap_8 FILLER_32_595 ();
 sg13g2_decap_8 FILLER_32_602 ();
 sg13g2_decap_8 FILLER_32_609 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_decap_8 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_637 ();
 sg13g2_decap_8 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_decap_8 FILLER_32_658 ();
 sg13g2_decap_8 FILLER_32_665 ();
 sg13g2_decap_8 FILLER_32_672 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_8 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_700 ();
 sg13g2_decap_8 FILLER_32_707 ();
 sg13g2_decap_8 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_decap_8 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_decap_8 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_32_868 ();
 sg13g2_decap_8 FILLER_32_875 ();
 sg13g2_decap_8 FILLER_32_882 ();
 sg13g2_decap_8 FILLER_32_889 ();
 sg13g2_decap_8 FILLER_32_896 ();
 sg13g2_decap_8 FILLER_32_903 ();
 sg13g2_decap_8 FILLER_32_910 ();
 sg13g2_decap_8 FILLER_32_917 ();
 sg13g2_decap_8 FILLER_32_924 ();
 sg13g2_decap_8 FILLER_32_931 ();
 sg13g2_decap_8 FILLER_32_938 ();
 sg13g2_decap_8 FILLER_32_945 ();
 sg13g2_decap_8 FILLER_32_952 ();
 sg13g2_decap_8 FILLER_32_959 ();
 sg13g2_decap_8 FILLER_32_966 ();
 sg13g2_decap_8 FILLER_32_973 ();
 sg13g2_decap_8 FILLER_32_980 ();
 sg13g2_decap_8 FILLER_32_987 ();
 sg13g2_decap_8 FILLER_32_994 ();
 sg13g2_decap_8 FILLER_32_1001 ();
 sg13g2_decap_8 FILLER_32_1008 ();
 sg13g2_decap_8 FILLER_32_1015 ();
 sg13g2_decap_8 FILLER_32_1022 ();
 sg13g2_fill_1 FILLER_33_8 ();
 sg13g2_fill_1 FILLER_33_62 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_fill_2 FILLER_33_269 ();
 sg13g2_fill_1 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_313 ();
 sg13g2_fill_1 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_33_435 ();
 sg13g2_fill_2 FILLER_33_459 ();
 sg13g2_decap_8 FILLER_33_501 ();
 sg13g2_decap_8 FILLER_33_508 ();
 sg13g2_decap_8 FILLER_33_515 ();
 sg13g2_decap_8 FILLER_33_522 ();
 sg13g2_decap_8 FILLER_33_529 ();
 sg13g2_decap_8 FILLER_33_536 ();
 sg13g2_decap_8 FILLER_33_543 ();
 sg13g2_decap_8 FILLER_33_550 ();
 sg13g2_decap_8 FILLER_33_557 ();
 sg13g2_decap_8 FILLER_33_564 ();
 sg13g2_decap_8 FILLER_33_571 ();
 sg13g2_decap_8 FILLER_33_578 ();
 sg13g2_decap_8 FILLER_33_585 ();
 sg13g2_decap_8 FILLER_33_592 ();
 sg13g2_decap_8 FILLER_33_599 ();
 sg13g2_decap_8 FILLER_33_606 ();
 sg13g2_decap_8 FILLER_33_613 ();
 sg13g2_decap_8 FILLER_33_620 ();
 sg13g2_decap_8 FILLER_33_627 ();
 sg13g2_decap_8 FILLER_33_634 ();
 sg13g2_decap_8 FILLER_33_641 ();
 sg13g2_decap_8 FILLER_33_648 ();
 sg13g2_decap_8 FILLER_33_655 ();
 sg13g2_decap_8 FILLER_33_662 ();
 sg13g2_decap_8 FILLER_33_669 ();
 sg13g2_decap_8 FILLER_33_676 ();
 sg13g2_decap_8 FILLER_33_683 ();
 sg13g2_decap_8 FILLER_33_690 ();
 sg13g2_decap_8 FILLER_33_697 ();
 sg13g2_decap_8 FILLER_33_704 ();
 sg13g2_decap_8 FILLER_33_711 ();
 sg13g2_decap_8 FILLER_33_718 ();
 sg13g2_decap_8 FILLER_33_725 ();
 sg13g2_decap_8 FILLER_33_732 ();
 sg13g2_decap_8 FILLER_33_739 ();
 sg13g2_decap_8 FILLER_33_746 ();
 sg13g2_decap_8 FILLER_33_753 ();
 sg13g2_decap_8 FILLER_33_760 ();
 sg13g2_decap_8 FILLER_33_767 ();
 sg13g2_decap_8 FILLER_33_774 ();
 sg13g2_decap_8 FILLER_33_781 ();
 sg13g2_decap_8 FILLER_33_788 ();
 sg13g2_decap_8 FILLER_33_795 ();
 sg13g2_decap_8 FILLER_33_802 ();
 sg13g2_decap_8 FILLER_33_809 ();
 sg13g2_decap_8 FILLER_33_816 ();
 sg13g2_decap_8 FILLER_33_823 ();
 sg13g2_decap_8 FILLER_33_830 ();
 sg13g2_decap_8 FILLER_33_837 ();
 sg13g2_decap_8 FILLER_33_844 ();
 sg13g2_decap_8 FILLER_33_851 ();
 sg13g2_decap_8 FILLER_33_858 ();
 sg13g2_decap_8 FILLER_33_865 ();
 sg13g2_decap_8 FILLER_33_872 ();
 sg13g2_decap_8 FILLER_33_879 ();
 sg13g2_decap_8 FILLER_33_886 ();
 sg13g2_decap_8 FILLER_33_893 ();
 sg13g2_decap_8 FILLER_33_900 ();
 sg13g2_decap_8 FILLER_33_907 ();
 sg13g2_decap_8 FILLER_33_914 ();
 sg13g2_decap_8 FILLER_33_921 ();
 sg13g2_decap_8 FILLER_33_928 ();
 sg13g2_decap_8 FILLER_33_935 ();
 sg13g2_decap_8 FILLER_33_942 ();
 sg13g2_decap_8 FILLER_33_949 ();
 sg13g2_decap_8 FILLER_33_956 ();
 sg13g2_decap_8 FILLER_33_963 ();
 sg13g2_decap_8 FILLER_33_970 ();
 sg13g2_decap_8 FILLER_33_977 ();
 sg13g2_decap_8 FILLER_33_984 ();
 sg13g2_decap_8 FILLER_33_991 ();
 sg13g2_decap_8 FILLER_33_998 ();
 sg13g2_decap_8 FILLER_33_1005 ();
 sg13g2_decap_8 FILLER_33_1012 ();
 sg13g2_decap_8 FILLER_33_1019 ();
 sg13g2_fill_2 FILLER_33_1026 ();
 sg13g2_fill_1 FILLER_33_1028 ();
 sg13g2_fill_2 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_fill_2 FILLER_34_345 ();
 sg13g2_fill_1 FILLER_34_347 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_34_416 ();
 sg13g2_fill_2 FILLER_34_460 ();
 sg13g2_fill_1 FILLER_34_471 ();
 sg13g2_decap_8 FILLER_34_494 ();
 sg13g2_decap_8 FILLER_34_501 ();
 sg13g2_decap_8 FILLER_34_508 ();
 sg13g2_decap_8 FILLER_34_515 ();
 sg13g2_decap_8 FILLER_34_522 ();
 sg13g2_decap_8 FILLER_34_529 ();
 sg13g2_decap_8 FILLER_34_536 ();
 sg13g2_decap_8 FILLER_34_543 ();
 sg13g2_decap_8 FILLER_34_550 ();
 sg13g2_decap_8 FILLER_34_557 ();
 sg13g2_decap_8 FILLER_34_564 ();
 sg13g2_decap_8 FILLER_34_571 ();
 sg13g2_decap_8 FILLER_34_578 ();
 sg13g2_decap_8 FILLER_34_585 ();
 sg13g2_decap_8 FILLER_34_592 ();
 sg13g2_decap_8 FILLER_34_599 ();
 sg13g2_decap_8 FILLER_34_606 ();
 sg13g2_decap_8 FILLER_34_613 ();
 sg13g2_decap_8 FILLER_34_620 ();
 sg13g2_decap_8 FILLER_34_627 ();
 sg13g2_decap_8 FILLER_34_634 ();
 sg13g2_decap_8 FILLER_34_641 ();
 sg13g2_decap_8 FILLER_34_648 ();
 sg13g2_decap_8 FILLER_34_655 ();
 sg13g2_decap_8 FILLER_34_662 ();
 sg13g2_decap_8 FILLER_34_669 ();
 sg13g2_decap_8 FILLER_34_676 ();
 sg13g2_decap_8 FILLER_34_683 ();
 sg13g2_decap_8 FILLER_34_690 ();
 sg13g2_decap_8 FILLER_34_697 ();
 sg13g2_decap_8 FILLER_34_704 ();
 sg13g2_decap_8 FILLER_34_711 ();
 sg13g2_decap_8 FILLER_34_718 ();
 sg13g2_decap_8 FILLER_34_725 ();
 sg13g2_decap_8 FILLER_34_732 ();
 sg13g2_decap_8 FILLER_34_739 ();
 sg13g2_decap_8 FILLER_34_746 ();
 sg13g2_decap_8 FILLER_34_753 ();
 sg13g2_decap_8 FILLER_34_760 ();
 sg13g2_decap_8 FILLER_34_767 ();
 sg13g2_decap_8 FILLER_34_774 ();
 sg13g2_decap_8 FILLER_34_781 ();
 sg13g2_decap_8 FILLER_34_788 ();
 sg13g2_decap_8 FILLER_34_795 ();
 sg13g2_decap_8 FILLER_34_802 ();
 sg13g2_decap_8 FILLER_34_809 ();
 sg13g2_decap_8 FILLER_34_816 ();
 sg13g2_decap_8 FILLER_34_823 ();
 sg13g2_decap_8 FILLER_34_830 ();
 sg13g2_decap_8 FILLER_34_837 ();
 sg13g2_decap_8 FILLER_34_844 ();
 sg13g2_decap_8 FILLER_34_851 ();
 sg13g2_decap_8 FILLER_34_858 ();
 sg13g2_decap_8 FILLER_34_865 ();
 sg13g2_decap_8 FILLER_34_872 ();
 sg13g2_decap_8 FILLER_34_879 ();
 sg13g2_decap_8 FILLER_34_886 ();
 sg13g2_decap_8 FILLER_34_893 ();
 sg13g2_decap_8 FILLER_34_900 ();
 sg13g2_decap_8 FILLER_34_907 ();
 sg13g2_decap_8 FILLER_34_914 ();
 sg13g2_decap_8 FILLER_34_921 ();
 sg13g2_decap_8 FILLER_34_928 ();
 sg13g2_decap_8 FILLER_34_935 ();
 sg13g2_decap_8 FILLER_34_942 ();
 sg13g2_decap_8 FILLER_34_949 ();
 sg13g2_decap_8 FILLER_34_956 ();
 sg13g2_decap_8 FILLER_34_963 ();
 sg13g2_decap_8 FILLER_34_970 ();
 sg13g2_decap_8 FILLER_34_977 ();
 sg13g2_decap_8 FILLER_34_984 ();
 sg13g2_decap_8 FILLER_34_991 ();
 sg13g2_decap_8 FILLER_34_998 ();
 sg13g2_decap_8 FILLER_34_1005 ();
 sg13g2_decap_8 FILLER_34_1012 ();
 sg13g2_decap_8 FILLER_34_1019 ();
 sg13g2_fill_2 FILLER_34_1026 ();
 sg13g2_fill_1 FILLER_34_1028 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_68 ();
 sg13g2_fill_1 FILLER_35_88 ();
 sg13g2_fill_2 FILLER_35_109 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_2 FILLER_35_245 ();
 sg13g2_fill_1 FILLER_35_247 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_fill_1 FILLER_35_321 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_fill_2 FILLER_35_457 ();
 sg13g2_fill_1 FILLER_35_459 ();
 sg13g2_decap_8 FILLER_35_492 ();
 sg13g2_decap_8 FILLER_35_499 ();
 sg13g2_decap_8 FILLER_35_506 ();
 sg13g2_decap_8 FILLER_35_513 ();
 sg13g2_decap_8 FILLER_35_520 ();
 sg13g2_decap_8 FILLER_35_527 ();
 sg13g2_decap_8 FILLER_35_534 ();
 sg13g2_decap_8 FILLER_35_541 ();
 sg13g2_decap_8 FILLER_35_548 ();
 sg13g2_decap_8 FILLER_35_555 ();
 sg13g2_decap_8 FILLER_35_562 ();
 sg13g2_decap_8 FILLER_35_569 ();
 sg13g2_decap_8 FILLER_35_576 ();
 sg13g2_decap_8 FILLER_35_583 ();
 sg13g2_decap_8 FILLER_35_590 ();
 sg13g2_decap_8 FILLER_35_597 ();
 sg13g2_decap_8 FILLER_35_604 ();
 sg13g2_decap_8 FILLER_35_611 ();
 sg13g2_decap_8 FILLER_35_618 ();
 sg13g2_decap_8 FILLER_35_625 ();
 sg13g2_decap_8 FILLER_35_632 ();
 sg13g2_decap_8 FILLER_35_639 ();
 sg13g2_decap_8 FILLER_35_646 ();
 sg13g2_decap_8 FILLER_35_653 ();
 sg13g2_decap_8 FILLER_35_660 ();
 sg13g2_decap_8 FILLER_35_667 ();
 sg13g2_decap_8 FILLER_35_674 ();
 sg13g2_decap_8 FILLER_35_681 ();
 sg13g2_decap_8 FILLER_35_688 ();
 sg13g2_decap_8 FILLER_35_695 ();
 sg13g2_decap_8 FILLER_35_702 ();
 sg13g2_decap_8 FILLER_35_709 ();
 sg13g2_decap_8 FILLER_35_716 ();
 sg13g2_decap_8 FILLER_35_723 ();
 sg13g2_decap_8 FILLER_35_730 ();
 sg13g2_decap_8 FILLER_35_737 ();
 sg13g2_decap_8 FILLER_35_744 ();
 sg13g2_decap_8 FILLER_35_751 ();
 sg13g2_decap_8 FILLER_35_758 ();
 sg13g2_decap_8 FILLER_35_765 ();
 sg13g2_decap_8 FILLER_35_772 ();
 sg13g2_decap_8 FILLER_35_779 ();
 sg13g2_decap_8 FILLER_35_786 ();
 sg13g2_decap_8 FILLER_35_793 ();
 sg13g2_decap_8 FILLER_35_800 ();
 sg13g2_decap_8 FILLER_35_807 ();
 sg13g2_decap_8 FILLER_35_814 ();
 sg13g2_decap_8 FILLER_35_821 ();
 sg13g2_decap_8 FILLER_35_828 ();
 sg13g2_decap_8 FILLER_35_835 ();
 sg13g2_decap_8 FILLER_35_842 ();
 sg13g2_decap_8 FILLER_35_849 ();
 sg13g2_decap_8 FILLER_35_856 ();
 sg13g2_decap_8 FILLER_35_863 ();
 sg13g2_decap_8 FILLER_35_870 ();
 sg13g2_decap_8 FILLER_35_877 ();
 sg13g2_decap_8 FILLER_35_884 ();
 sg13g2_decap_8 FILLER_35_891 ();
 sg13g2_decap_8 FILLER_35_898 ();
 sg13g2_decap_8 FILLER_35_905 ();
 sg13g2_decap_8 FILLER_35_912 ();
 sg13g2_decap_8 FILLER_35_919 ();
 sg13g2_decap_8 FILLER_35_926 ();
 sg13g2_decap_8 FILLER_35_933 ();
 sg13g2_decap_8 FILLER_35_940 ();
 sg13g2_decap_8 FILLER_35_947 ();
 sg13g2_decap_8 FILLER_35_954 ();
 sg13g2_decap_8 FILLER_35_961 ();
 sg13g2_decap_8 FILLER_35_968 ();
 sg13g2_decap_8 FILLER_35_975 ();
 sg13g2_decap_8 FILLER_35_982 ();
 sg13g2_decap_8 FILLER_35_989 ();
 sg13g2_decap_8 FILLER_35_996 ();
 sg13g2_decap_8 FILLER_35_1003 ();
 sg13g2_decap_8 FILLER_35_1010 ();
 sg13g2_decap_8 FILLER_35_1017 ();
 sg13g2_decap_4 FILLER_35_1024 ();
 sg13g2_fill_1 FILLER_35_1028 ();
 sg13g2_fill_1 FILLER_36_8 ();
 sg13g2_fill_2 FILLER_36_41 ();
 sg13g2_fill_2 FILLER_36_85 ();
 sg13g2_fill_1 FILLER_36_87 ();
 sg13g2_fill_1 FILLER_36_110 ();
 sg13g2_fill_2 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_fill_2 FILLER_36_437 ();
 sg13g2_decap_8 FILLER_36_493 ();
 sg13g2_decap_8 FILLER_36_500 ();
 sg13g2_decap_8 FILLER_36_507 ();
 sg13g2_decap_8 FILLER_36_514 ();
 sg13g2_decap_8 FILLER_36_521 ();
 sg13g2_decap_8 FILLER_36_528 ();
 sg13g2_decap_8 FILLER_36_535 ();
 sg13g2_decap_8 FILLER_36_542 ();
 sg13g2_decap_8 FILLER_36_549 ();
 sg13g2_decap_8 FILLER_36_556 ();
 sg13g2_decap_8 FILLER_36_563 ();
 sg13g2_decap_8 FILLER_36_570 ();
 sg13g2_decap_8 FILLER_36_577 ();
 sg13g2_decap_8 FILLER_36_584 ();
 sg13g2_decap_8 FILLER_36_591 ();
 sg13g2_decap_8 FILLER_36_598 ();
 sg13g2_decap_8 FILLER_36_605 ();
 sg13g2_decap_8 FILLER_36_612 ();
 sg13g2_decap_8 FILLER_36_619 ();
 sg13g2_decap_8 FILLER_36_626 ();
 sg13g2_decap_8 FILLER_36_633 ();
 sg13g2_decap_8 FILLER_36_640 ();
 sg13g2_decap_8 FILLER_36_647 ();
 sg13g2_decap_8 FILLER_36_654 ();
 sg13g2_decap_8 FILLER_36_661 ();
 sg13g2_decap_8 FILLER_36_668 ();
 sg13g2_decap_8 FILLER_36_675 ();
 sg13g2_decap_8 FILLER_36_682 ();
 sg13g2_decap_8 FILLER_36_689 ();
 sg13g2_decap_8 FILLER_36_696 ();
 sg13g2_decap_8 FILLER_36_703 ();
 sg13g2_decap_8 FILLER_36_710 ();
 sg13g2_decap_8 FILLER_36_717 ();
 sg13g2_decap_8 FILLER_36_724 ();
 sg13g2_decap_8 FILLER_36_731 ();
 sg13g2_decap_8 FILLER_36_738 ();
 sg13g2_decap_8 FILLER_36_745 ();
 sg13g2_decap_8 FILLER_36_752 ();
 sg13g2_decap_8 FILLER_36_759 ();
 sg13g2_decap_8 FILLER_36_766 ();
 sg13g2_decap_8 FILLER_36_773 ();
 sg13g2_decap_8 FILLER_36_780 ();
 sg13g2_decap_8 FILLER_36_787 ();
 sg13g2_decap_8 FILLER_36_794 ();
 sg13g2_decap_8 FILLER_36_801 ();
 sg13g2_decap_8 FILLER_36_808 ();
 sg13g2_decap_8 FILLER_36_815 ();
 sg13g2_decap_8 FILLER_36_822 ();
 sg13g2_decap_8 FILLER_36_829 ();
 sg13g2_decap_8 FILLER_36_836 ();
 sg13g2_decap_8 FILLER_36_843 ();
 sg13g2_decap_8 FILLER_36_850 ();
 sg13g2_decap_8 FILLER_36_857 ();
 sg13g2_decap_8 FILLER_36_864 ();
 sg13g2_decap_8 FILLER_36_871 ();
 sg13g2_decap_8 FILLER_36_878 ();
 sg13g2_decap_8 FILLER_36_885 ();
 sg13g2_decap_8 FILLER_36_892 ();
 sg13g2_decap_8 FILLER_36_899 ();
 sg13g2_decap_8 FILLER_36_906 ();
 sg13g2_decap_8 FILLER_36_913 ();
 sg13g2_decap_8 FILLER_36_920 ();
 sg13g2_decap_8 FILLER_36_927 ();
 sg13g2_decap_8 FILLER_36_934 ();
 sg13g2_decap_8 FILLER_36_941 ();
 sg13g2_decap_8 FILLER_36_948 ();
 sg13g2_decap_8 FILLER_36_955 ();
 sg13g2_decap_8 FILLER_36_962 ();
 sg13g2_decap_8 FILLER_36_969 ();
 sg13g2_decap_8 FILLER_36_976 ();
 sg13g2_decap_8 FILLER_36_983 ();
 sg13g2_decap_8 FILLER_36_990 ();
 sg13g2_decap_8 FILLER_36_997 ();
 sg13g2_decap_8 FILLER_36_1004 ();
 sg13g2_decap_8 FILLER_36_1011 ();
 sg13g2_decap_8 FILLER_36_1018 ();
 sg13g2_decap_4 FILLER_36_1025 ();
 sg13g2_fill_2 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_125 ();
 sg13g2_fill_2 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_174 ();
 sg13g2_fill_2 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_275 ();
 sg13g2_fill_1 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_437 ();
 sg13g2_decap_4 FILLER_37_473 ();
 sg13g2_decap_8 FILLER_37_499 ();
 sg13g2_decap_8 FILLER_37_506 ();
 sg13g2_decap_8 FILLER_37_513 ();
 sg13g2_decap_8 FILLER_37_520 ();
 sg13g2_decap_8 FILLER_37_527 ();
 sg13g2_decap_8 FILLER_37_534 ();
 sg13g2_decap_8 FILLER_37_541 ();
 sg13g2_decap_8 FILLER_37_548 ();
 sg13g2_decap_8 FILLER_37_555 ();
 sg13g2_decap_8 FILLER_37_562 ();
 sg13g2_decap_8 FILLER_37_569 ();
 sg13g2_decap_8 FILLER_37_576 ();
 sg13g2_decap_8 FILLER_37_583 ();
 sg13g2_decap_8 FILLER_37_590 ();
 sg13g2_decap_8 FILLER_37_597 ();
 sg13g2_decap_8 FILLER_37_604 ();
 sg13g2_decap_8 FILLER_37_611 ();
 sg13g2_decap_8 FILLER_37_618 ();
 sg13g2_decap_8 FILLER_37_625 ();
 sg13g2_decap_8 FILLER_37_632 ();
 sg13g2_decap_8 FILLER_37_639 ();
 sg13g2_decap_8 FILLER_37_646 ();
 sg13g2_decap_8 FILLER_37_653 ();
 sg13g2_decap_8 FILLER_37_660 ();
 sg13g2_decap_8 FILLER_37_667 ();
 sg13g2_decap_8 FILLER_37_674 ();
 sg13g2_decap_8 FILLER_37_681 ();
 sg13g2_decap_8 FILLER_37_688 ();
 sg13g2_decap_8 FILLER_37_695 ();
 sg13g2_decap_8 FILLER_37_702 ();
 sg13g2_decap_8 FILLER_37_709 ();
 sg13g2_decap_8 FILLER_37_716 ();
 sg13g2_decap_8 FILLER_37_723 ();
 sg13g2_decap_8 FILLER_37_730 ();
 sg13g2_decap_8 FILLER_37_737 ();
 sg13g2_decap_8 FILLER_37_744 ();
 sg13g2_decap_8 FILLER_37_751 ();
 sg13g2_decap_8 FILLER_37_758 ();
 sg13g2_decap_8 FILLER_37_765 ();
 sg13g2_decap_8 FILLER_37_772 ();
 sg13g2_decap_8 FILLER_37_779 ();
 sg13g2_decap_8 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_793 ();
 sg13g2_decap_8 FILLER_37_800 ();
 sg13g2_decap_8 FILLER_37_807 ();
 sg13g2_decap_8 FILLER_37_814 ();
 sg13g2_decap_8 FILLER_37_821 ();
 sg13g2_decap_8 FILLER_37_828 ();
 sg13g2_decap_8 FILLER_37_835 ();
 sg13g2_decap_8 FILLER_37_842 ();
 sg13g2_decap_8 FILLER_37_849 ();
 sg13g2_decap_8 FILLER_37_856 ();
 sg13g2_decap_8 FILLER_37_863 ();
 sg13g2_decap_8 FILLER_37_870 ();
 sg13g2_decap_8 FILLER_37_877 ();
 sg13g2_decap_8 FILLER_37_884 ();
 sg13g2_decap_8 FILLER_37_891 ();
 sg13g2_decap_8 FILLER_37_898 ();
 sg13g2_decap_8 FILLER_37_905 ();
 sg13g2_decap_8 FILLER_37_912 ();
 sg13g2_decap_8 FILLER_37_919 ();
 sg13g2_decap_8 FILLER_37_926 ();
 sg13g2_decap_8 FILLER_37_933 ();
 sg13g2_decap_8 FILLER_37_940 ();
 sg13g2_decap_8 FILLER_37_947 ();
 sg13g2_decap_8 FILLER_37_954 ();
 sg13g2_decap_8 FILLER_37_961 ();
 sg13g2_decap_8 FILLER_37_968 ();
 sg13g2_decap_8 FILLER_37_975 ();
 sg13g2_decap_8 FILLER_37_982 ();
 sg13g2_decap_8 FILLER_37_989 ();
 sg13g2_decap_8 FILLER_37_996 ();
 sg13g2_decap_8 FILLER_37_1003 ();
 sg13g2_decap_8 FILLER_37_1010 ();
 sg13g2_decap_8 FILLER_37_1017 ();
 sg13g2_decap_4 FILLER_37_1024 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_48 ();
 sg13g2_fill_2 FILLER_38_65 ();
 sg13g2_fill_2 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_86 ();
 sg13g2_fill_1 FILLER_38_88 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_1 FILLER_38_320 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_399 ();
 sg13g2_fill_1 FILLER_38_458 ();
 sg13g2_fill_2 FILLER_38_468 ();
 sg13g2_fill_1 FILLER_38_470 ();
 sg13g2_decap_8 FILLER_38_480 ();
 sg13g2_decap_8 FILLER_38_487 ();
 sg13g2_decap_8 FILLER_38_494 ();
 sg13g2_decap_8 FILLER_38_501 ();
 sg13g2_decap_8 FILLER_38_508 ();
 sg13g2_decap_8 FILLER_38_515 ();
 sg13g2_decap_8 FILLER_38_522 ();
 sg13g2_decap_8 FILLER_38_529 ();
 sg13g2_decap_8 FILLER_38_536 ();
 sg13g2_decap_8 FILLER_38_543 ();
 sg13g2_decap_8 FILLER_38_550 ();
 sg13g2_decap_8 FILLER_38_557 ();
 sg13g2_decap_8 FILLER_38_564 ();
 sg13g2_decap_8 FILLER_38_571 ();
 sg13g2_decap_8 FILLER_38_578 ();
 sg13g2_decap_8 FILLER_38_585 ();
 sg13g2_decap_8 FILLER_38_592 ();
 sg13g2_decap_8 FILLER_38_599 ();
 sg13g2_decap_8 FILLER_38_606 ();
 sg13g2_decap_8 FILLER_38_613 ();
 sg13g2_decap_8 FILLER_38_620 ();
 sg13g2_decap_8 FILLER_38_627 ();
 sg13g2_decap_8 FILLER_38_634 ();
 sg13g2_decap_8 FILLER_38_641 ();
 sg13g2_decap_8 FILLER_38_648 ();
 sg13g2_decap_8 FILLER_38_655 ();
 sg13g2_decap_8 FILLER_38_662 ();
 sg13g2_decap_8 FILLER_38_669 ();
 sg13g2_decap_8 FILLER_38_676 ();
 sg13g2_decap_8 FILLER_38_683 ();
 sg13g2_decap_8 FILLER_38_690 ();
 sg13g2_decap_8 FILLER_38_697 ();
 sg13g2_decap_8 FILLER_38_704 ();
 sg13g2_decap_8 FILLER_38_711 ();
 sg13g2_decap_8 FILLER_38_718 ();
 sg13g2_decap_8 FILLER_38_725 ();
 sg13g2_decap_8 FILLER_38_732 ();
 sg13g2_decap_8 FILLER_38_739 ();
 sg13g2_decap_8 FILLER_38_746 ();
 sg13g2_decap_8 FILLER_38_753 ();
 sg13g2_decap_8 FILLER_38_760 ();
 sg13g2_decap_8 FILLER_38_767 ();
 sg13g2_decap_8 FILLER_38_774 ();
 sg13g2_decap_8 FILLER_38_781 ();
 sg13g2_decap_8 FILLER_38_788 ();
 sg13g2_decap_8 FILLER_38_795 ();
 sg13g2_decap_8 FILLER_38_802 ();
 sg13g2_decap_8 FILLER_38_809 ();
 sg13g2_decap_8 FILLER_38_816 ();
 sg13g2_decap_8 FILLER_38_823 ();
 sg13g2_decap_8 FILLER_38_830 ();
 sg13g2_decap_8 FILLER_38_837 ();
 sg13g2_decap_8 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_decap_8 FILLER_38_858 ();
 sg13g2_decap_8 FILLER_38_865 ();
 sg13g2_decap_8 FILLER_38_872 ();
 sg13g2_decap_8 FILLER_38_879 ();
 sg13g2_decap_8 FILLER_38_886 ();
 sg13g2_decap_8 FILLER_38_893 ();
 sg13g2_decap_8 FILLER_38_900 ();
 sg13g2_decap_8 FILLER_38_907 ();
 sg13g2_decap_8 FILLER_38_914 ();
 sg13g2_decap_8 FILLER_38_921 ();
 sg13g2_decap_8 FILLER_38_928 ();
 sg13g2_decap_8 FILLER_38_935 ();
 sg13g2_decap_8 FILLER_38_942 ();
 sg13g2_decap_8 FILLER_38_949 ();
 sg13g2_decap_8 FILLER_38_956 ();
 sg13g2_decap_8 FILLER_38_963 ();
 sg13g2_decap_8 FILLER_38_970 ();
 sg13g2_decap_8 FILLER_38_977 ();
 sg13g2_decap_8 FILLER_38_984 ();
 sg13g2_decap_8 FILLER_38_991 ();
 sg13g2_decap_8 FILLER_38_998 ();
 sg13g2_decap_8 FILLER_38_1005 ();
 sg13g2_decap_8 FILLER_38_1012 ();
 sg13g2_decap_8 FILLER_38_1019 ();
 sg13g2_fill_2 FILLER_38_1026 ();
 sg13g2_fill_1 FILLER_38_1028 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_71 ();
 sg13g2_fill_1 FILLER_39_102 ();
 sg13g2_fill_2 FILLER_39_161 ();
 sg13g2_fill_2 FILLER_39_168 ();
 sg13g2_fill_2 FILLER_39_212 ();
 sg13g2_fill_1 FILLER_39_226 ();
 sg13g2_fill_2 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_332 ();
 sg13g2_fill_1 FILLER_39_361 ();
 sg13g2_fill_2 FILLER_39_367 ();
 sg13g2_fill_2 FILLER_39_397 ();
 sg13g2_decap_8 FILLER_39_467 ();
 sg13g2_decap_8 FILLER_39_474 ();
 sg13g2_decap_8 FILLER_39_481 ();
 sg13g2_decap_8 FILLER_39_488 ();
 sg13g2_decap_8 FILLER_39_495 ();
 sg13g2_decap_8 FILLER_39_502 ();
 sg13g2_decap_8 FILLER_39_509 ();
 sg13g2_decap_8 FILLER_39_516 ();
 sg13g2_decap_8 FILLER_39_523 ();
 sg13g2_decap_8 FILLER_39_530 ();
 sg13g2_decap_8 FILLER_39_537 ();
 sg13g2_decap_8 FILLER_39_544 ();
 sg13g2_decap_8 FILLER_39_551 ();
 sg13g2_decap_8 FILLER_39_558 ();
 sg13g2_decap_8 FILLER_39_565 ();
 sg13g2_decap_8 FILLER_39_572 ();
 sg13g2_decap_8 FILLER_39_579 ();
 sg13g2_decap_8 FILLER_39_586 ();
 sg13g2_decap_8 FILLER_39_593 ();
 sg13g2_decap_8 FILLER_39_600 ();
 sg13g2_decap_8 FILLER_39_607 ();
 sg13g2_decap_8 FILLER_39_614 ();
 sg13g2_decap_8 FILLER_39_621 ();
 sg13g2_decap_8 FILLER_39_628 ();
 sg13g2_decap_8 FILLER_39_635 ();
 sg13g2_decap_8 FILLER_39_642 ();
 sg13g2_decap_8 FILLER_39_649 ();
 sg13g2_decap_8 FILLER_39_656 ();
 sg13g2_decap_8 FILLER_39_663 ();
 sg13g2_decap_8 FILLER_39_670 ();
 sg13g2_decap_8 FILLER_39_677 ();
 sg13g2_decap_8 FILLER_39_684 ();
 sg13g2_decap_8 FILLER_39_691 ();
 sg13g2_decap_8 FILLER_39_698 ();
 sg13g2_decap_8 FILLER_39_705 ();
 sg13g2_decap_8 FILLER_39_712 ();
 sg13g2_decap_8 FILLER_39_719 ();
 sg13g2_decap_8 FILLER_39_726 ();
 sg13g2_decap_8 FILLER_39_733 ();
 sg13g2_decap_8 FILLER_39_740 ();
 sg13g2_decap_8 FILLER_39_747 ();
 sg13g2_decap_8 FILLER_39_754 ();
 sg13g2_decap_8 FILLER_39_761 ();
 sg13g2_decap_8 FILLER_39_768 ();
 sg13g2_decap_8 FILLER_39_775 ();
 sg13g2_decap_8 FILLER_39_782 ();
 sg13g2_decap_8 FILLER_39_789 ();
 sg13g2_decap_8 FILLER_39_796 ();
 sg13g2_decap_8 FILLER_39_803 ();
 sg13g2_decap_8 FILLER_39_810 ();
 sg13g2_decap_8 FILLER_39_817 ();
 sg13g2_decap_8 FILLER_39_824 ();
 sg13g2_decap_8 FILLER_39_831 ();
 sg13g2_decap_8 FILLER_39_838 ();
 sg13g2_decap_8 FILLER_39_845 ();
 sg13g2_decap_8 FILLER_39_852 ();
 sg13g2_decap_8 FILLER_39_859 ();
 sg13g2_decap_8 FILLER_39_866 ();
 sg13g2_decap_8 FILLER_39_873 ();
 sg13g2_decap_8 FILLER_39_880 ();
 sg13g2_decap_8 FILLER_39_887 ();
 sg13g2_decap_8 FILLER_39_894 ();
 sg13g2_decap_8 FILLER_39_901 ();
 sg13g2_decap_8 FILLER_39_908 ();
 sg13g2_decap_8 FILLER_39_915 ();
 sg13g2_decap_8 FILLER_39_922 ();
 sg13g2_decap_8 FILLER_39_929 ();
 sg13g2_decap_8 FILLER_39_936 ();
 sg13g2_decap_8 FILLER_39_943 ();
 sg13g2_decap_8 FILLER_39_950 ();
 sg13g2_decap_8 FILLER_39_957 ();
 sg13g2_decap_8 FILLER_39_964 ();
 sg13g2_decap_8 FILLER_39_971 ();
 sg13g2_decap_8 FILLER_39_978 ();
 sg13g2_decap_8 FILLER_39_985 ();
 sg13g2_decap_8 FILLER_39_992 ();
 sg13g2_decap_8 FILLER_39_999 ();
 sg13g2_decap_8 FILLER_39_1006 ();
 sg13g2_decap_8 FILLER_39_1013 ();
 sg13g2_decap_8 FILLER_39_1020 ();
 sg13g2_fill_2 FILLER_39_1027 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_35 ();
 sg13g2_fill_2 FILLER_40_47 ();
 sg13g2_fill_2 FILLER_40_89 ();
 sg13g2_fill_1 FILLER_40_107 ();
 sg13g2_fill_1 FILLER_40_132 ();
 sg13g2_fill_2 FILLER_40_146 ();
 sg13g2_fill_1 FILLER_40_148 ();
 sg13g2_fill_2 FILLER_40_176 ();
 sg13g2_fill_2 FILLER_40_202 ();
 sg13g2_fill_1 FILLER_40_226 ();
 sg13g2_fill_1 FILLER_40_276 ();
 sg13g2_fill_1 FILLER_40_291 ();
 sg13g2_decap_4 FILLER_40_297 ();
 sg13g2_fill_2 FILLER_40_301 ();
 sg13g2_fill_1 FILLER_40_357 ();
 sg13g2_fill_2 FILLER_40_441 ();
 sg13g2_fill_2 FILLER_40_453 ();
 sg13g2_decap_8 FILLER_40_459 ();
 sg13g2_decap_8 FILLER_40_466 ();
 sg13g2_decap_8 FILLER_40_473 ();
 sg13g2_decap_8 FILLER_40_480 ();
 sg13g2_decap_8 FILLER_40_487 ();
 sg13g2_decap_8 FILLER_40_494 ();
 sg13g2_decap_8 FILLER_40_501 ();
 sg13g2_decap_8 FILLER_40_508 ();
 sg13g2_decap_8 FILLER_40_515 ();
 sg13g2_decap_8 FILLER_40_522 ();
 sg13g2_decap_8 FILLER_40_529 ();
 sg13g2_decap_8 FILLER_40_536 ();
 sg13g2_decap_8 FILLER_40_543 ();
 sg13g2_decap_8 FILLER_40_550 ();
 sg13g2_decap_8 FILLER_40_557 ();
 sg13g2_decap_8 FILLER_40_564 ();
 sg13g2_decap_8 FILLER_40_571 ();
 sg13g2_decap_8 FILLER_40_578 ();
 sg13g2_decap_8 FILLER_40_585 ();
 sg13g2_decap_8 FILLER_40_592 ();
 sg13g2_decap_8 FILLER_40_599 ();
 sg13g2_decap_8 FILLER_40_606 ();
 sg13g2_decap_8 FILLER_40_613 ();
 sg13g2_decap_8 FILLER_40_620 ();
 sg13g2_decap_8 FILLER_40_627 ();
 sg13g2_decap_8 FILLER_40_634 ();
 sg13g2_decap_8 FILLER_40_641 ();
 sg13g2_decap_8 FILLER_40_648 ();
 sg13g2_decap_8 FILLER_40_655 ();
 sg13g2_decap_8 FILLER_40_662 ();
 sg13g2_decap_8 FILLER_40_669 ();
 sg13g2_decap_8 FILLER_40_676 ();
 sg13g2_decap_8 FILLER_40_683 ();
 sg13g2_decap_8 FILLER_40_690 ();
 sg13g2_decap_8 FILLER_40_697 ();
 sg13g2_decap_8 FILLER_40_704 ();
 sg13g2_decap_8 FILLER_40_711 ();
 sg13g2_decap_8 FILLER_40_718 ();
 sg13g2_decap_8 FILLER_40_725 ();
 sg13g2_decap_8 FILLER_40_732 ();
 sg13g2_decap_8 FILLER_40_739 ();
 sg13g2_decap_8 FILLER_40_746 ();
 sg13g2_decap_8 FILLER_40_753 ();
 sg13g2_decap_8 FILLER_40_760 ();
 sg13g2_decap_8 FILLER_40_767 ();
 sg13g2_decap_8 FILLER_40_774 ();
 sg13g2_decap_8 FILLER_40_781 ();
 sg13g2_decap_8 FILLER_40_788 ();
 sg13g2_decap_8 FILLER_40_795 ();
 sg13g2_decap_8 FILLER_40_802 ();
 sg13g2_decap_8 FILLER_40_809 ();
 sg13g2_decap_8 FILLER_40_816 ();
 sg13g2_decap_8 FILLER_40_823 ();
 sg13g2_decap_8 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_837 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_8 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_40_865 ();
 sg13g2_decap_8 FILLER_40_872 ();
 sg13g2_decap_8 FILLER_40_879 ();
 sg13g2_decap_8 FILLER_40_886 ();
 sg13g2_decap_8 FILLER_40_893 ();
 sg13g2_decap_8 FILLER_40_900 ();
 sg13g2_decap_8 FILLER_40_907 ();
 sg13g2_decap_8 FILLER_40_914 ();
 sg13g2_decap_8 FILLER_40_921 ();
 sg13g2_decap_8 FILLER_40_928 ();
 sg13g2_decap_8 FILLER_40_935 ();
 sg13g2_decap_8 FILLER_40_942 ();
 sg13g2_decap_8 FILLER_40_949 ();
 sg13g2_decap_8 FILLER_40_956 ();
 sg13g2_decap_8 FILLER_40_963 ();
 sg13g2_decap_8 FILLER_40_970 ();
 sg13g2_decap_8 FILLER_40_977 ();
 sg13g2_decap_8 FILLER_40_984 ();
 sg13g2_decap_8 FILLER_40_991 ();
 sg13g2_decap_8 FILLER_40_998 ();
 sg13g2_decap_8 FILLER_40_1005 ();
 sg13g2_decap_8 FILLER_40_1012 ();
 sg13g2_decap_8 FILLER_40_1019 ();
 sg13g2_fill_2 FILLER_40_1026 ();
 sg13g2_fill_1 FILLER_40_1028 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_80 ();
 sg13g2_fill_1 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_107 ();
 sg13g2_fill_2 FILLER_41_126 ();
 sg13g2_fill_2 FILLER_41_144 ();
 sg13g2_fill_1 FILLER_41_146 ();
 sg13g2_fill_1 FILLER_41_253 ();
 sg13g2_fill_2 FILLER_41_282 ();
 sg13g2_fill_1 FILLER_41_326 ();
 sg13g2_fill_1 FILLER_41_355 ();
 sg13g2_decap_4 FILLER_41_367 ();
 sg13g2_decap_4 FILLER_41_418 ();
 sg13g2_fill_2 FILLER_41_422 ();
 sg13g2_fill_2 FILLER_41_438 ();
 sg13g2_decap_8 FILLER_41_451 ();
 sg13g2_decap_8 FILLER_41_458 ();
 sg13g2_decap_8 FILLER_41_465 ();
 sg13g2_decap_8 FILLER_41_472 ();
 sg13g2_decap_8 FILLER_41_479 ();
 sg13g2_decap_8 FILLER_41_486 ();
 sg13g2_decap_8 FILLER_41_493 ();
 sg13g2_decap_8 FILLER_41_500 ();
 sg13g2_decap_8 FILLER_41_507 ();
 sg13g2_decap_8 FILLER_41_514 ();
 sg13g2_decap_8 FILLER_41_521 ();
 sg13g2_decap_8 FILLER_41_528 ();
 sg13g2_decap_8 FILLER_41_535 ();
 sg13g2_decap_8 FILLER_41_542 ();
 sg13g2_decap_8 FILLER_41_549 ();
 sg13g2_decap_8 FILLER_41_556 ();
 sg13g2_decap_8 FILLER_41_563 ();
 sg13g2_decap_8 FILLER_41_570 ();
 sg13g2_decap_8 FILLER_41_577 ();
 sg13g2_decap_8 FILLER_41_584 ();
 sg13g2_decap_8 FILLER_41_591 ();
 sg13g2_decap_8 FILLER_41_598 ();
 sg13g2_decap_8 FILLER_41_605 ();
 sg13g2_decap_8 FILLER_41_612 ();
 sg13g2_decap_8 FILLER_41_619 ();
 sg13g2_decap_8 FILLER_41_626 ();
 sg13g2_decap_8 FILLER_41_633 ();
 sg13g2_decap_8 FILLER_41_640 ();
 sg13g2_decap_8 FILLER_41_647 ();
 sg13g2_decap_8 FILLER_41_654 ();
 sg13g2_decap_8 FILLER_41_661 ();
 sg13g2_decap_8 FILLER_41_668 ();
 sg13g2_decap_8 FILLER_41_675 ();
 sg13g2_decap_8 FILLER_41_682 ();
 sg13g2_decap_8 FILLER_41_689 ();
 sg13g2_decap_8 FILLER_41_696 ();
 sg13g2_decap_8 FILLER_41_703 ();
 sg13g2_decap_8 FILLER_41_710 ();
 sg13g2_decap_8 FILLER_41_717 ();
 sg13g2_decap_8 FILLER_41_724 ();
 sg13g2_decap_8 FILLER_41_731 ();
 sg13g2_decap_8 FILLER_41_738 ();
 sg13g2_decap_8 FILLER_41_745 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_decap_8 FILLER_41_759 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_decap_8 FILLER_41_773 ();
 sg13g2_decap_8 FILLER_41_780 ();
 sg13g2_decap_8 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_794 ();
 sg13g2_decap_8 FILLER_41_801 ();
 sg13g2_decap_8 FILLER_41_808 ();
 sg13g2_decap_8 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_850 ();
 sg13g2_decap_8 FILLER_41_857 ();
 sg13g2_decap_8 FILLER_41_864 ();
 sg13g2_decap_8 FILLER_41_871 ();
 sg13g2_decap_8 FILLER_41_878 ();
 sg13g2_decap_8 FILLER_41_885 ();
 sg13g2_decap_8 FILLER_41_892 ();
 sg13g2_decap_8 FILLER_41_899 ();
 sg13g2_decap_8 FILLER_41_906 ();
 sg13g2_decap_8 FILLER_41_913 ();
 sg13g2_decap_8 FILLER_41_920 ();
 sg13g2_decap_8 FILLER_41_927 ();
 sg13g2_decap_8 FILLER_41_934 ();
 sg13g2_decap_8 FILLER_41_941 ();
 sg13g2_decap_8 FILLER_41_948 ();
 sg13g2_decap_8 FILLER_41_955 ();
 sg13g2_decap_8 FILLER_41_962 ();
 sg13g2_decap_8 FILLER_41_969 ();
 sg13g2_decap_8 FILLER_41_976 ();
 sg13g2_decap_8 FILLER_41_983 ();
 sg13g2_decap_8 FILLER_41_990 ();
 sg13g2_decap_8 FILLER_41_997 ();
 sg13g2_decap_8 FILLER_41_1004 ();
 sg13g2_decap_8 FILLER_41_1011 ();
 sg13g2_decap_8 FILLER_41_1018 ();
 sg13g2_decap_4 FILLER_41_1025 ();
 sg13g2_fill_2 FILLER_42_38 ();
 sg13g2_fill_2 FILLER_42_48 ();
 sg13g2_fill_1 FILLER_42_87 ();
 sg13g2_fill_1 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_129 ();
 sg13g2_fill_1 FILLER_42_131 ();
 sg13g2_fill_2 FILLER_42_155 ();
 sg13g2_fill_2 FILLER_42_250 ();
 sg13g2_fill_1 FILLER_42_252 ();
 sg13g2_fill_2 FILLER_42_317 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_fill_1 FILLER_42_351 ();
 sg13g2_fill_2 FILLER_42_395 ();
 sg13g2_fill_2 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_42_433 ();
 sg13g2_decap_8 FILLER_42_440 ();
 sg13g2_decap_8 FILLER_42_447 ();
 sg13g2_decap_8 FILLER_42_454 ();
 sg13g2_decap_8 FILLER_42_461 ();
 sg13g2_decap_8 FILLER_42_468 ();
 sg13g2_decap_8 FILLER_42_475 ();
 sg13g2_decap_8 FILLER_42_482 ();
 sg13g2_decap_8 FILLER_42_489 ();
 sg13g2_decap_8 FILLER_42_496 ();
 sg13g2_decap_8 FILLER_42_503 ();
 sg13g2_decap_8 FILLER_42_510 ();
 sg13g2_decap_8 FILLER_42_517 ();
 sg13g2_decap_8 FILLER_42_524 ();
 sg13g2_decap_8 FILLER_42_531 ();
 sg13g2_decap_8 FILLER_42_538 ();
 sg13g2_decap_8 FILLER_42_545 ();
 sg13g2_decap_8 FILLER_42_552 ();
 sg13g2_decap_8 FILLER_42_559 ();
 sg13g2_decap_8 FILLER_42_566 ();
 sg13g2_decap_8 FILLER_42_573 ();
 sg13g2_decap_8 FILLER_42_580 ();
 sg13g2_decap_8 FILLER_42_587 ();
 sg13g2_decap_8 FILLER_42_594 ();
 sg13g2_decap_8 FILLER_42_601 ();
 sg13g2_decap_8 FILLER_42_608 ();
 sg13g2_decap_8 FILLER_42_615 ();
 sg13g2_decap_8 FILLER_42_622 ();
 sg13g2_decap_8 FILLER_42_629 ();
 sg13g2_decap_8 FILLER_42_636 ();
 sg13g2_decap_8 FILLER_42_643 ();
 sg13g2_decap_8 FILLER_42_650 ();
 sg13g2_decap_8 FILLER_42_657 ();
 sg13g2_decap_8 FILLER_42_664 ();
 sg13g2_decap_8 FILLER_42_671 ();
 sg13g2_decap_8 FILLER_42_678 ();
 sg13g2_decap_8 FILLER_42_685 ();
 sg13g2_decap_8 FILLER_42_692 ();
 sg13g2_decap_8 FILLER_42_699 ();
 sg13g2_decap_8 FILLER_42_706 ();
 sg13g2_decap_8 FILLER_42_713 ();
 sg13g2_decap_8 FILLER_42_720 ();
 sg13g2_decap_8 FILLER_42_727 ();
 sg13g2_decap_8 FILLER_42_734 ();
 sg13g2_decap_8 FILLER_42_741 ();
 sg13g2_decap_8 FILLER_42_748 ();
 sg13g2_decap_8 FILLER_42_755 ();
 sg13g2_decap_8 FILLER_42_762 ();
 sg13g2_decap_8 FILLER_42_769 ();
 sg13g2_decap_8 FILLER_42_776 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_decap_8 FILLER_42_790 ();
 sg13g2_decap_8 FILLER_42_797 ();
 sg13g2_decap_8 FILLER_42_804 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_846 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_decap_8 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_42_867 ();
 sg13g2_decap_8 FILLER_42_874 ();
 sg13g2_decap_8 FILLER_42_881 ();
 sg13g2_decap_8 FILLER_42_888 ();
 sg13g2_decap_8 FILLER_42_895 ();
 sg13g2_decap_8 FILLER_42_902 ();
 sg13g2_decap_8 FILLER_42_909 ();
 sg13g2_decap_8 FILLER_42_916 ();
 sg13g2_decap_8 FILLER_42_923 ();
 sg13g2_decap_8 FILLER_42_930 ();
 sg13g2_decap_8 FILLER_42_937 ();
 sg13g2_decap_8 FILLER_42_944 ();
 sg13g2_decap_8 FILLER_42_951 ();
 sg13g2_decap_8 FILLER_42_958 ();
 sg13g2_decap_8 FILLER_42_965 ();
 sg13g2_decap_8 FILLER_42_972 ();
 sg13g2_decap_8 FILLER_42_979 ();
 sg13g2_decap_8 FILLER_42_986 ();
 sg13g2_decap_8 FILLER_42_993 ();
 sg13g2_decap_8 FILLER_42_1000 ();
 sg13g2_decap_8 FILLER_42_1007 ();
 sg13g2_decap_8 FILLER_42_1014 ();
 sg13g2_decap_8 FILLER_42_1021 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_105 ();
 sg13g2_fill_2 FILLER_43_128 ();
 sg13g2_fill_1 FILLER_43_298 ();
 sg13g2_decap_8 FILLER_43_404 ();
 sg13g2_decap_8 FILLER_43_411 ();
 sg13g2_decap_8 FILLER_43_418 ();
 sg13g2_decap_8 FILLER_43_425 ();
 sg13g2_decap_8 FILLER_43_432 ();
 sg13g2_decap_8 FILLER_43_439 ();
 sg13g2_decap_8 FILLER_43_446 ();
 sg13g2_decap_8 FILLER_43_453 ();
 sg13g2_decap_8 FILLER_43_460 ();
 sg13g2_decap_8 FILLER_43_467 ();
 sg13g2_decap_8 FILLER_43_474 ();
 sg13g2_decap_8 FILLER_43_481 ();
 sg13g2_decap_8 FILLER_43_488 ();
 sg13g2_decap_8 FILLER_43_495 ();
 sg13g2_decap_8 FILLER_43_502 ();
 sg13g2_decap_8 FILLER_43_509 ();
 sg13g2_decap_8 FILLER_43_516 ();
 sg13g2_decap_8 FILLER_43_523 ();
 sg13g2_decap_8 FILLER_43_530 ();
 sg13g2_decap_8 FILLER_43_537 ();
 sg13g2_decap_8 FILLER_43_544 ();
 sg13g2_decap_8 FILLER_43_551 ();
 sg13g2_decap_8 FILLER_43_558 ();
 sg13g2_decap_8 FILLER_43_565 ();
 sg13g2_decap_8 FILLER_43_572 ();
 sg13g2_decap_8 FILLER_43_579 ();
 sg13g2_decap_8 FILLER_43_586 ();
 sg13g2_decap_8 FILLER_43_593 ();
 sg13g2_decap_8 FILLER_43_600 ();
 sg13g2_decap_8 FILLER_43_607 ();
 sg13g2_decap_8 FILLER_43_614 ();
 sg13g2_decap_8 FILLER_43_621 ();
 sg13g2_decap_8 FILLER_43_628 ();
 sg13g2_decap_8 FILLER_43_635 ();
 sg13g2_decap_8 FILLER_43_642 ();
 sg13g2_decap_8 FILLER_43_649 ();
 sg13g2_decap_8 FILLER_43_656 ();
 sg13g2_decap_8 FILLER_43_663 ();
 sg13g2_decap_8 FILLER_43_670 ();
 sg13g2_decap_8 FILLER_43_677 ();
 sg13g2_decap_8 FILLER_43_684 ();
 sg13g2_decap_8 FILLER_43_691 ();
 sg13g2_decap_8 FILLER_43_698 ();
 sg13g2_decap_8 FILLER_43_705 ();
 sg13g2_decap_8 FILLER_43_712 ();
 sg13g2_decap_8 FILLER_43_719 ();
 sg13g2_decap_8 FILLER_43_726 ();
 sg13g2_decap_8 FILLER_43_733 ();
 sg13g2_decap_8 FILLER_43_740 ();
 sg13g2_decap_8 FILLER_43_747 ();
 sg13g2_decap_8 FILLER_43_754 ();
 sg13g2_decap_8 FILLER_43_761 ();
 sg13g2_decap_8 FILLER_43_768 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_8 FILLER_43_782 ();
 sg13g2_decap_8 FILLER_43_789 ();
 sg13g2_decap_8 FILLER_43_796 ();
 sg13g2_decap_8 FILLER_43_803 ();
 sg13g2_decap_8 FILLER_43_810 ();
 sg13g2_decap_8 FILLER_43_817 ();
 sg13g2_decap_8 FILLER_43_824 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_8 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_decap_8 FILLER_43_859 ();
 sg13g2_decap_8 FILLER_43_866 ();
 sg13g2_decap_8 FILLER_43_873 ();
 sg13g2_decap_8 FILLER_43_880 ();
 sg13g2_decap_8 FILLER_43_887 ();
 sg13g2_decap_8 FILLER_43_894 ();
 sg13g2_decap_8 FILLER_43_901 ();
 sg13g2_decap_8 FILLER_43_908 ();
 sg13g2_decap_8 FILLER_43_915 ();
 sg13g2_decap_8 FILLER_43_922 ();
 sg13g2_decap_8 FILLER_43_929 ();
 sg13g2_decap_8 FILLER_43_936 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_decap_8 FILLER_43_950 ();
 sg13g2_decap_8 FILLER_43_957 ();
 sg13g2_decap_8 FILLER_43_964 ();
 sg13g2_decap_8 FILLER_43_971 ();
 sg13g2_decap_8 FILLER_43_978 ();
 sg13g2_decap_8 FILLER_43_985 ();
 sg13g2_decap_8 FILLER_43_992 ();
 sg13g2_decap_8 FILLER_43_999 ();
 sg13g2_decap_8 FILLER_43_1006 ();
 sg13g2_decap_8 FILLER_43_1013 ();
 sg13g2_decap_8 FILLER_43_1020 ();
 sg13g2_fill_2 FILLER_43_1027 ();
 sg13g2_fill_1 FILLER_44_8 ();
 sg13g2_fill_2 FILLER_44_68 ();
 sg13g2_fill_2 FILLER_44_98 ();
 sg13g2_fill_1 FILLER_44_106 ();
 sg13g2_fill_2 FILLER_44_111 ();
 sg13g2_fill_1 FILLER_44_113 ();
 sg13g2_fill_2 FILLER_44_119 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_fill_2 FILLER_44_157 ();
 sg13g2_fill_2 FILLER_44_210 ();
 sg13g2_fill_2 FILLER_44_226 ();
 sg13g2_fill_2 FILLER_44_246 ();
 sg13g2_fill_2 FILLER_44_305 ();
 sg13g2_decap_4 FILLER_44_313 ();
 sg13g2_fill_2 FILLER_44_317 ();
 sg13g2_fill_2 FILLER_44_348 ();
 sg13g2_fill_1 FILLER_44_350 ();
 sg13g2_decap_4 FILLER_44_359 ();
 sg13g2_decap_4 FILLER_44_376 ();
 sg13g2_fill_2 FILLER_44_380 ();
 sg13g2_decap_8 FILLER_44_388 ();
 sg13g2_decap_8 FILLER_44_395 ();
 sg13g2_decap_8 FILLER_44_402 ();
 sg13g2_decap_8 FILLER_44_409 ();
 sg13g2_decap_8 FILLER_44_416 ();
 sg13g2_decap_8 FILLER_44_423 ();
 sg13g2_decap_8 FILLER_44_430 ();
 sg13g2_decap_8 FILLER_44_437 ();
 sg13g2_decap_8 FILLER_44_444 ();
 sg13g2_decap_8 FILLER_44_451 ();
 sg13g2_decap_8 FILLER_44_458 ();
 sg13g2_decap_8 FILLER_44_465 ();
 sg13g2_decap_8 FILLER_44_472 ();
 sg13g2_decap_8 FILLER_44_479 ();
 sg13g2_decap_8 FILLER_44_486 ();
 sg13g2_decap_8 FILLER_44_493 ();
 sg13g2_decap_8 FILLER_44_500 ();
 sg13g2_decap_8 FILLER_44_507 ();
 sg13g2_decap_8 FILLER_44_514 ();
 sg13g2_decap_8 FILLER_44_521 ();
 sg13g2_decap_8 FILLER_44_528 ();
 sg13g2_decap_8 FILLER_44_535 ();
 sg13g2_decap_8 FILLER_44_542 ();
 sg13g2_decap_8 FILLER_44_549 ();
 sg13g2_decap_8 FILLER_44_556 ();
 sg13g2_decap_8 FILLER_44_563 ();
 sg13g2_decap_8 FILLER_44_570 ();
 sg13g2_decap_8 FILLER_44_577 ();
 sg13g2_decap_8 FILLER_44_584 ();
 sg13g2_decap_8 FILLER_44_591 ();
 sg13g2_decap_8 FILLER_44_598 ();
 sg13g2_decap_8 FILLER_44_605 ();
 sg13g2_decap_8 FILLER_44_612 ();
 sg13g2_decap_8 FILLER_44_619 ();
 sg13g2_decap_8 FILLER_44_626 ();
 sg13g2_decap_8 FILLER_44_633 ();
 sg13g2_decap_8 FILLER_44_640 ();
 sg13g2_decap_8 FILLER_44_647 ();
 sg13g2_decap_8 FILLER_44_654 ();
 sg13g2_decap_8 FILLER_44_661 ();
 sg13g2_decap_8 FILLER_44_668 ();
 sg13g2_decap_8 FILLER_44_675 ();
 sg13g2_decap_8 FILLER_44_682 ();
 sg13g2_decap_8 FILLER_44_689 ();
 sg13g2_decap_8 FILLER_44_696 ();
 sg13g2_decap_8 FILLER_44_703 ();
 sg13g2_decap_8 FILLER_44_710 ();
 sg13g2_decap_8 FILLER_44_717 ();
 sg13g2_decap_8 FILLER_44_724 ();
 sg13g2_decap_8 FILLER_44_731 ();
 sg13g2_decap_8 FILLER_44_738 ();
 sg13g2_decap_8 FILLER_44_745 ();
 sg13g2_decap_8 FILLER_44_752 ();
 sg13g2_decap_8 FILLER_44_759 ();
 sg13g2_decap_8 FILLER_44_766 ();
 sg13g2_decap_8 FILLER_44_773 ();
 sg13g2_decap_8 FILLER_44_780 ();
 sg13g2_decap_8 FILLER_44_787 ();
 sg13g2_decap_8 FILLER_44_794 ();
 sg13g2_decap_8 FILLER_44_801 ();
 sg13g2_decap_8 FILLER_44_808 ();
 sg13g2_decap_8 FILLER_44_815 ();
 sg13g2_decap_8 FILLER_44_822 ();
 sg13g2_decap_8 FILLER_44_829 ();
 sg13g2_decap_8 FILLER_44_836 ();
 sg13g2_decap_8 FILLER_44_843 ();
 sg13g2_decap_8 FILLER_44_850 ();
 sg13g2_decap_8 FILLER_44_857 ();
 sg13g2_decap_8 FILLER_44_864 ();
 sg13g2_decap_8 FILLER_44_871 ();
 sg13g2_decap_8 FILLER_44_878 ();
 sg13g2_decap_8 FILLER_44_885 ();
 sg13g2_decap_8 FILLER_44_892 ();
 sg13g2_decap_8 FILLER_44_899 ();
 sg13g2_decap_8 FILLER_44_906 ();
 sg13g2_decap_8 FILLER_44_913 ();
 sg13g2_decap_8 FILLER_44_920 ();
 sg13g2_decap_8 FILLER_44_927 ();
 sg13g2_decap_8 FILLER_44_934 ();
 sg13g2_decap_8 FILLER_44_941 ();
 sg13g2_decap_8 FILLER_44_948 ();
 sg13g2_decap_8 FILLER_44_955 ();
 sg13g2_decap_8 FILLER_44_962 ();
 sg13g2_decap_8 FILLER_44_969 ();
 sg13g2_decap_8 FILLER_44_976 ();
 sg13g2_decap_8 FILLER_44_983 ();
 sg13g2_decap_8 FILLER_44_990 ();
 sg13g2_decap_8 FILLER_44_997 ();
 sg13g2_decap_8 FILLER_44_1004 ();
 sg13g2_decap_8 FILLER_44_1011 ();
 sg13g2_decap_8 FILLER_44_1018 ();
 sg13g2_decap_4 FILLER_44_1025 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_41 ();
 sg13g2_fill_2 FILLER_45_66 ();
 sg13g2_fill_2 FILLER_45_157 ();
 sg13g2_fill_1 FILLER_45_159 ();
 sg13g2_fill_1 FILLER_45_195 ();
 sg13g2_fill_1 FILLER_45_214 ();
 sg13g2_fill_2 FILLER_45_271 ();
 sg13g2_fill_1 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_fill_2 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_fill_1 FILLER_45_349 ();
 sg13g2_decap_8 FILLER_45_373 ();
 sg13g2_decap_8 FILLER_45_380 ();
 sg13g2_decap_8 FILLER_45_387 ();
 sg13g2_decap_8 FILLER_45_394 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_decap_8 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_45_415 ();
 sg13g2_decap_8 FILLER_45_422 ();
 sg13g2_decap_8 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_45_436 ();
 sg13g2_decap_8 FILLER_45_443 ();
 sg13g2_decap_8 FILLER_45_450 ();
 sg13g2_decap_8 FILLER_45_457 ();
 sg13g2_decap_8 FILLER_45_464 ();
 sg13g2_decap_8 FILLER_45_471 ();
 sg13g2_decap_8 FILLER_45_478 ();
 sg13g2_decap_8 FILLER_45_485 ();
 sg13g2_decap_8 FILLER_45_492 ();
 sg13g2_decap_8 FILLER_45_499 ();
 sg13g2_decap_8 FILLER_45_506 ();
 sg13g2_decap_8 FILLER_45_513 ();
 sg13g2_decap_8 FILLER_45_520 ();
 sg13g2_decap_8 FILLER_45_527 ();
 sg13g2_decap_8 FILLER_45_534 ();
 sg13g2_decap_8 FILLER_45_541 ();
 sg13g2_decap_8 FILLER_45_548 ();
 sg13g2_decap_8 FILLER_45_555 ();
 sg13g2_decap_8 FILLER_45_562 ();
 sg13g2_decap_8 FILLER_45_569 ();
 sg13g2_decap_8 FILLER_45_576 ();
 sg13g2_decap_8 FILLER_45_583 ();
 sg13g2_decap_8 FILLER_45_590 ();
 sg13g2_decap_8 FILLER_45_597 ();
 sg13g2_decap_8 FILLER_45_604 ();
 sg13g2_decap_8 FILLER_45_611 ();
 sg13g2_decap_8 FILLER_45_618 ();
 sg13g2_decap_8 FILLER_45_625 ();
 sg13g2_decap_8 FILLER_45_632 ();
 sg13g2_decap_8 FILLER_45_639 ();
 sg13g2_decap_8 FILLER_45_646 ();
 sg13g2_decap_8 FILLER_45_653 ();
 sg13g2_decap_8 FILLER_45_660 ();
 sg13g2_decap_8 FILLER_45_667 ();
 sg13g2_decap_8 FILLER_45_674 ();
 sg13g2_decap_8 FILLER_45_681 ();
 sg13g2_decap_8 FILLER_45_688 ();
 sg13g2_decap_8 FILLER_45_695 ();
 sg13g2_decap_8 FILLER_45_702 ();
 sg13g2_decap_8 FILLER_45_709 ();
 sg13g2_decap_8 FILLER_45_716 ();
 sg13g2_decap_8 FILLER_45_723 ();
 sg13g2_decap_8 FILLER_45_730 ();
 sg13g2_decap_8 FILLER_45_737 ();
 sg13g2_decap_8 FILLER_45_744 ();
 sg13g2_decap_8 FILLER_45_751 ();
 sg13g2_decap_8 FILLER_45_758 ();
 sg13g2_decap_8 FILLER_45_765 ();
 sg13g2_decap_8 FILLER_45_772 ();
 sg13g2_decap_8 FILLER_45_779 ();
 sg13g2_decap_8 FILLER_45_786 ();
 sg13g2_decap_8 FILLER_45_793 ();
 sg13g2_decap_8 FILLER_45_800 ();
 sg13g2_decap_8 FILLER_45_807 ();
 sg13g2_decap_8 FILLER_45_814 ();
 sg13g2_decap_8 FILLER_45_821 ();
 sg13g2_decap_8 FILLER_45_828 ();
 sg13g2_decap_8 FILLER_45_835 ();
 sg13g2_decap_8 FILLER_45_842 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_decap_8 FILLER_45_856 ();
 sg13g2_decap_8 FILLER_45_863 ();
 sg13g2_decap_8 FILLER_45_870 ();
 sg13g2_decap_8 FILLER_45_877 ();
 sg13g2_decap_8 FILLER_45_884 ();
 sg13g2_decap_8 FILLER_45_891 ();
 sg13g2_decap_8 FILLER_45_898 ();
 sg13g2_decap_8 FILLER_45_905 ();
 sg13g2_decap_8 FILLER_45_912 ();
 sg13g2_decap_8 FILLER_45_919 ();
 sg13g2_decap_8 FILLER_45_926 ();
 sg13g2_decap_8 FILLER_45_933 ();
 sg13g2_decap_8 FILLER_45_940 ();
 sg13g2_decap_8 FILLER_45_947 ();
 sg13g2_decap_8 FILLER_45_954 ();
 sg13g2_decap_8 FILLER_45_961 ();
 sg13g2_decap_8 FILLER_45_968 ();
 sg13g2_decap_8 FILLER_45_975 ();
 sg13g2_decap_8 FILLER_45_982 ();
 sg13g2_decap_8 FILLER_45_989 ();
 sg13g2_decap_8 FILLER_45_996 ();
 sg13g2_decap_8 FILLER_45_1003 ();
 sg13g2_decap_8 FILLER_45_1010 ();
 sg13g2_decap_8 FILLER_45_1017 ();
 sg13g2_decap_4 FILLER_45_1024 ();
 sg13g2_fill_1 FILLER_45_1028 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_1 FILLER_46_69 ();
 sg13g2_fill_1 FILLER_46_76 ();
 sg13g2_fill_2 FILLER_46_120 ();
 sg13g2_fill_1 FILLER_46_127 ();
 sg13g2_fill_1 FILLER_46_137 ();
 sg13g2_fill_2 FILLER_46_154 ();
 sg13g2_fill_2 FILLER_46_173 ();
 sg13g2_fill_2 FILLER_46_228 ();
 sg13g2_fill_2 FILLER_46_240 ();
 sg13g2_fill_2 FILLER_46_277 ();
 sg13g2_fill_2 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_344 ();
 sg13g2_decap_8 FILLER_46_351 ();
 sg13g2_decap_4 FILLER_46_358 ();
 sg13g2_decap_8 FILLER_46_367 ();
 sg13g2_decap_8 FILLER_46_374 ();
 sg13g2_decap_8 FILLER_46_381 ();
 sg13g2_decap_8 FILLER_46_388 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_decap_8 FILLER_46_409 ();
 sg13g2_decap_8 FILLER_46_416 ();
 sg13g2_decap_8 FILLER_46_423 ();
 sg13g2_decap_8 FILLER_46_430 ();
 sg13g2_decap_8 FILLER_46_437 ();
 sg13g2_decap_8 FILLER_46_444 ();
 sg13g2_decap_8 FILLER_46_451 ();
 sg13g2_decap_8 FILLER_46_458 ();
 sg13g2_decap_8 FILLER_46_465 ();
 sg13g2_decap_8 FILLER_46_472 ();
 sg13g2_decap_8 FILLER_46_479 ();
 sg13g2_decap_8 FILLER_46_486 ();
 sg13g2_decap_8 FILLER_46_493 ();
 sg13g2_decap_8 FILLER_46_500 ();
 sg13g2_decap_8 FILLER_46_507 ();
 sg13g2_decap_8 FILLER_46_514 ();
 sg13g2_decap_8 FILLER_46_521 ();
 sg13g2_decap_8 FILLER_46_528 ();
 sg13g2_decap_8 FILLER_46_535 ();
 sg13g2_decap_8 FILLER_46_542 ();
 sg13g2_decap_8 FILLER_46_549 ();
 sg13g2_decap_8 FILLER_46_556 ();
 sg13g2_decap_8 FILLER_46_563 ();
 sg13g2_decap_8 FILLER_46_570 ();
 sg13g2_decap_8 FILLER_46_577 ();
 sg13g2_decap_8 FILLER_46_584 ();
 sg13g2_decap_8 FILLER_46_591 ();
 sg13g2_decap_8 FILLER_46_598 ();
 sg13g2_decap_8 FILLER_46_605 ();
 sg13g2_decap_8 FILLER_46_612 ();
 sg13g2_decap_8 FILLER_46_619 ();
 sg13g2_decap_8 FILLER_46_626 ();
 sg13g2_decap_8 FILLER_46_633 ();
 sg13g2_decap_8 FILLER_46_640 ();
 sg13g2_decap_8 FILLER_46_647 ();
 sg13g2_decap_8 FILLER_46_654 ();
 sg13g2_decap_8 FILLER_46_661 ();
 sg13g2_decap_8 FILLER_46_668 ();
 sg13g2_decap_8 FILLER_46_675 ();
 sg13g2_decap_8 FILLER_46_682 ();
 sg13g2_decap_8 FILLER_46_689 ();
 sg13g2_decap_8 FILLER_46_696 ();
 sg13g2_decap_8 FILLER_46_703 ();
 sg13g2_decap_8 FILLER_46_710 ();
 sg13g2_decap_8 FILLER_46_717 ();
 sg13g2_decap_8 FILLER_46_724 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_738 ();
 sg13g2_decap_8 FILLER_46_745 ();
 sg13g2_decap_8 FILLER_46_752 ();
 sg13g2_decap_8 FILLER_46_759 ();
 sg13g2_decap_8 FILLER_46_766 ();
 sg13g2_decap_8 FILLER_46_773 ();
 sg13g2_decap_8 FILLER_46_780 ();
 sg13g2_decap_8 FILLER_46_787 ();
 sg13g2_decap_8 FILLER_46_794 ();
 sg13g2_decap_8 FILLER_46_801 ();
 sg13g2_decap_8 FILLER_46_808 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_8 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_8 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_843 ();
 sg13g2_decap_8 FILLER_46_850 ();
 sg13g2_decap_8 FILLER_46_857 ();
 sg13g2_decap_8 FILLER_46_864 ();
 sg13g2_decap_8 FILLER_46_871 ();
 sg13g2_decap_8 FILLER_46_878 ();
 sg13g2_decap_8 FILLER_46_885 ();
 sg13g2_decap_8 FILLER_46_892 ();
 sg13g2_decap_8 FILLER_46_899 ();
 sg13g2_decap_8 FILLER_46_906 ();
 sg13g2_decap_8 FILLER_46_913 ();
 sg13g2_decap_8 FILLER_46_920 ();
 sg13g2_decap_8 FILLER_46_927 ();
 sg13g2_decap_8 FILLER_46_934 ();
 sg13g2_decap_8 FILLER_46_941 ();
 sg13g2_decap_8 FILLER_46_948 ();
 sg13g2_decap_8 FILLER_46_955 ();
 sg13g2_decap_8 FILLER_46_962 ();
 sg13g2_decap_8 FILLER_46_969 ();
 sg13g2_decap_8 FILLER_46_976 ();
 sg13g2_decap_8 FILLER_46_983 ();
 sg13g2_decap_8 FILLER_46_990 ();
 sg13g2_decap_8 FILLER_46_997 ();
 sg13g2_decap_8 FILLER_46_1004 ();
 sg13g2_decap_8 FILLER_46_1011 ();
 sg13g2_decap_8 FILLER_46_1018 ();
 sg13g2_decap_4 FILLER_46_1025 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_9 ();
 sg13g2_fill_2 FILLER_47_27 ();
 sg13g2_fill_1 FILLER_47_46 ();
 sg13g2_fill_2 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_150 ();
 sg13g2_fill_1 FILLER_47_216 ();
 sg13g2_fill_2 FILLER_47_279 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_4 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_332 ();
 sg13g2_decap_8 FILLER_47_339 ();
 sg13g2_decap_8 FILLER_47_346 ();
 sg13g2_decap_8 FILLER_47_353 ();
 sg13g2_decap_8 FILLER_47_360 ();
 sg13g2_decap_8 FILLER_47_367 ();
 sg13g2_decap_8 FILLER_47_374 ();
 sg13g2_decap_8 FILLER_47_381 ();
 sg13g2_decap_8 FILLER_47_388 ();
 sg13g2_decap_8 FILLER_47_395 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_decap_8 FILLER_47_409 ();
 sg13g2_decap_8 FILLER_47_416 ();
 sg13g2_decap_8 FILLER_47_423 ();
 sg13g2_decap_8 FILLER_47_430 ();
 sg13g2_decap_8 FILLER_47_437 ();
 sg13g2_decap_8 FILLER_47_444 ();
 sg13g2_decap_8 FILLER_47_451 ();
 sg13g2_decap_8 FILLER_47_458 ();
 sg13g2_decap_8 FILLER_47_465 ();
 sg13g2_decap_8 FILLER_47_472 ();
 sg13g2_decap_8 FILLER_47_479 ();
 sg13g2_decap_8 FILLER_47_486 ();
 sg13g2_decap_8 FILLER_47_493 ();
 sg13g2_decap_8 FILLER_47_500 ();
 sg13g2_decap_8 FILLER_47_507 ();
 sg13g2_decap_8 FILLER_47_514 ();
 sg13g2_decap_8 FILLER_47_521 ();
 sg13g2_decap_8 FILLER_47_528 ();
 sg13g2_decap_8 FILLER_47_535 ();
 sg13g2_decap_8 FILLER_47_542 ();
 sg13g2_decap_8 FILLER_47_549 ();
 sg13g2_decap_8 FILLER_47_556 ();
 sg13g2_decap_8 FILLER_47_563 ();
 sg13g2_decap_8 FILLER_47_570 ();
 sg13g2_decap_8 FILLER_47_577 ();
 sg13g2_decap_8 FILLER_47_584 ();
 sg13g2_decap_8 FILLER_47_591 ();
 sg13g2_decap_8 FILLER_47_598 ();
 sg13g2_decap_8 FILLER_47_605 ();
 sg13g2_decap_8 FILLER_47_612 ();
 sg13g2_decap_8 FILLER_47_619 ();
 sg13g2_decap_8 FILLER_47_626 ();
 sg13g2_decap_8 FILLER_47_633 ();
 sg13g2_decap_8 FILLER_47_640 ();
 sg13g2_decap_8 FILLER_47_647 ();
 sg13g2_decap_8 FILLER_47_654 ();
 sg13g2_decap_8 FILLER_47_661 ();
 sg13g2_decap_8 FILLER_47_668 ();
 sg13g2_decap_8 FILLER_47_675 ();
 sg13g2_decap_8 FILLER_47_682 ();
 sg13g2_decap_8 FILLER_47_689 ();
 sg13g2_decap_8 FILLER_47_696 ();
 sg13g2_decap_8 FILLER_47_703 ();
 sg13g2_decap_8 FILLER_47_710 ();
 sg13g2_decap_8 FILLER_47_717 ();
 sg13g2_decap_8 FILLER_47_724 ();
 sg13g2_decap_8 FILLER_47_731 ();
 sg13g2_decap_8 FILLER_47_738 ();
 sg13g2_decap_8 FILLER_47_745 ();
 sg13g2_decap_8 FILLER_47_752 ();
 sg13g2_decap_8 FILLER_47_759 ();
 sg13g2_decap_8 FILLER_47_766 ();
 sg13g2_decap_8 FILLER_47_773 ();
 sg13g2_decap_8 FILLER_47_780 ();
 sg13g2_decap_8 FILLER_47_787 ();
 sg13g2_decap_8 FILLER_47_794 ();
 sg13g2_decap_8 FILLER_47_801 ();
 sg13g2_decap_8 FILLER_47_808 ();
 sg13g2_decap_8 FILLER_47_815 ();
 sg13g2_decap_8 FILLER_47_822 ();
 sg13g2_decap_8 FILLER_47_829 ();
 sg13g2_decap_8 FILLER_47_836 ();
 sg13g2_decap_8 FILLER_47_843 ();
 sg13g2_decap_8 FILLER_47_850 ();
 sg13g2_decap_8 FILLER_47_857 ();
 sg13g2_decap_8 FILLER_47_864 ();
 sg13g2_decap_8 FILLER_47_871 ();
 sg13g2_decap_8 FILLER_47_878 ();
 sg13g2_decap_8 FILLER_47_885 ();
 sg13g2_decap_8 FILLER_47_892 ();
 sg13g2_decap_8 FILLER_47_899 ();
 sg13g2_decap_8 FILLER_47_906 ();
 sg13g2_decap_8 FILLER_47_913 ();
 sg13g2_decap_8 FILLER_47_920 ();
 sg13g2_decap_8 FILLER_47_927 ();
 sg13g2_decap_8 FILLER_47_934 ();
 sg13g2_decap_8 FILLER_47_941 ();
 sg13g2_decap_8 FILLER_47_948 ();
 sg13g2_decap_8 FILLER_47_955 ();
 sg13g2_decap_8 FILLER_47_962 ();
 sg13g2_decap_8 FILLER_47_969 ();
 sg13g2_decap_8 FILLER_47_976 ();
 sg13g2_decap_8 FILLER_47_983 ();
 sg13g2_decap_8 FILLER_47_990 ();
 sg13g2_decap_8 FILLER_47_997 ();
 sg13g2_decap_8 FILLER_47_1004 ();
 sg13g2_decap_8 FILLER_47_1011 ();
 sg13g2_decap_8 FILLER_47_1018 ();
 sg13g2_decap_4 FILLER_47_1025 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_318 ();
 sg13g2_decap_8 FILLER_48_325 ();
 sg13g2_decap_8 FILLER_48_332 ();
 sg13g2_decap_8 FILLER_48_339 ();
 sg13g2_decap_8 FILLER_48_346 ();
 sg13g2_decap_8 FILLER_48_353 ();
 sg13g2_decap_8 FILLER_48_360 ();
 sg13g2_decap_8 FILLER_48_367 ();
 sg13g2_decap_8 FILLER_48_374 ();
 sg13g2_decap_8 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_48_388 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_48_409 ();
 sg13g2_decap_8 FILLER_48_416 ();
 sg13g2_decap_8 FILLER_48_423 ();
 sg13g2_decap_8 FILLER_48_430 ();
 sg13g2_decap_8 FILLER_48_437 ();
 sg13g2_decap_8 FILLER_48_444 ();
 sg13g2_decap_8 FILLER_48_451 ();
 sg13g2_decap_8 FILLER_48_458 ();
 sg13g2_decap_8 FILLER_48_465 ();
 sg13g2_decap_8 FILLER_48_472 ();
 sg13g2_decap_8 FILLER_48_479 ();
 sg13g2_decap_8 FILLER_48_486 ();
 sg13g2_decap_8 FILLER_48_493 ();
 sg13g2_decap_8 FILLER_48_500 ();
 sg13g2_decap_8 FILLER_48_507 ();
 sg13g2_decap_8 FILLER_48_514 ();
 sg13g2_decap_8 FILLER_48_521 ();
 sg13g2_decap_8 FILLER_48_528 ();
 sg13g2_decap_8 FILLER_48_535 ();
 sg13g2_decap_8 FILLER_48_542 ();
 sg13g2_decap_8 FILLER_48_549 ();
 sg13g2_decap_8 FILLER_48_556 ();
 sg13g2_decap_8 FILLER_48_563 ();
 sg13g2_decap_8 FILLER_48_570 ();
 sg13g2_decap_8 FILLER_48_577 ();
 sg13g2_decap_8 FILLER_48_584 ();
 sg13g2_decap_8 FILLER_48_591 ();
 sg13g2_decap_8 FILLER_48_598 ();
 sg13g2_decap_8 FILLER_48_605 ();
 sg13g2_decap_8 FILLER_48_612 ();
 sg13g2_decap_8 FILLER_48_619 ();
 sg13g2_decap_8 FILLER_48_626 ();
 sg13g2_decap_8 FILLER_48_633 ();
 sg13g2_decap_8 FILLER_48_640 ();
 sg13g2_decap_8 FILLER_48_647 ();
 sg13g2_decap_8 FILLER_48_654 ();
 sg13g2_decap_8 FILLER_48_661 ();
 sg13g2_decap_8 FILLER_48_668 ();
 sg13g2_decap_8 FILLER_48_675 ();
 sg13g2_decap_8 FILLER_48_682 ();
 sg13g2_decap_8 FILLER_48_689 ();
 sg13g2_decap_8 FILLER_48_696 ();
 sg13g2_decap_8 FILLER_48_703 ();
 sg13g2_decap_8 FILLER_48_710 ();
 sg13g2_decap_8 FILLER_48_717 ();
 sg13g2_decap_8 FILLER_48_724 ();
 sg13g2_decap_8 FILLER_48_731 ();
 sg13g2_decap_8 FILLER_48_738 ();
 sg13g2_decap_8 FILLER_48_745 ();
 sg13g2_decap_8 FILLER_48_752 ();
 sg13g2_decap_8 FILLER_48_759 ();
 sg13g2_decap_8 FILLER_48_766 ();
 sg13g2_decap_8 FILLER_48_773 ();
 sg13g2_decap_8 FILLER_48_780 ();
 sg13g2_decap_8 FILLER_48_787 ();
 sg13g2_decap_8 FILLER_48_794 ();
 sg13g2_decap_8 FILLER_48_801 ();
 sg13g2_decap_8 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_850 ();
 sg13g2_decap_8 FILLER_48_857 ();
 sg13g2_decap_8 FILLER_48_864 ();
 sg13g2_decap_8 FILLER_48_871 ();
 sg13g2_decap_8 FILLER_48_878 ();
 sg13g2_decap_8 FILLER_48_885 ();
 sg13g2_decap_8 FILLER_48_892 ();
 sg13g2_decap_8 FILLER_48_899 ();
 sg13g2_decap_8 FILLER_48_906 ();
 sg13g2_decap_8 FILLER_48_913 ();
 sg13g2_decap_8 FILLER_48_920 ();
 sg13g2_decap_8 FILLER_48_927 ();
 sg13g2_decap_8 FILLER_48_934 ();
 sg13g2_decap_8 FILLER_48_941 ();
 sg13g2_decap_8 FILLER_48_948 ();
 sg13g2_decap_8 FILLER_48_955 ();
 sg13g2_decap_8 FILLER_48_962 ();
 sg13g2_decap_8 FILLER_48_969 ();
 sg13g2_decap_8 FILLER_48_976 ();
 sg13g2_decap_8 FILLER_48_983 ();
 sg13g2_decap_8 FILLER_48_990 ();
 sg13g2_decap_8 FILLER_48_997 ();
 sg13g2_decap_8 FILLER_48_1004 ();
 sg13g2_decap_8 FILLER_48_1011 ();
 sg13g2_decap_8 FILLER_48_1018 ();
 sg13g2_decap_4 FILLER_48_1025 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_23 ();
 sg13g2_fill_2 FILLER_49_187 ();
 sg13g2_fill_1 FILLER_49_244 ();
 sg13g2_decap_4 FILLER_49_270 ();
 sg13g2_fill_2 FILLER_49_279 ();
 sg13g2_decap_8 FILLER_49_291 ();
 sg13g2_decap_8 FILLER_49_311 ();
 sg13g2_decap_8 FILLER_49_318 ();
 sg13g2_decap_8 FILLER_49_325 ();
 sg13g2_decap_8 FILLER_49_332 ();
 sg13g2_decap_8 FILLER_49_339 ();
 sg13g2_decap_8 FILLER_49_346 ();
 sg13g2_decap_8 FILLER_49_353 ();
 sg13g2_decap_8 FILLER_49_360 ();
 sg13g2_decap_8 FILLER_49_367 ();
 sg13g2_decap_8 FILLER_49_374 ();
 sg13g2_decap_8 FILLER_49_381 ();
 sg13g2_decap_8 FILLER_49_388 ();
 sg13g2_decap_8 FILLER_49_395 ();
 sg13g2_decap_8 FILLER_49_402 ();
 sg13g2_decap_8 FILLER_49_409 ();
 sg13g2_decap_8 FILLER_49_416 ();
 sg13g2_decap_8 FILLER_49_423 ();
 sg13g2_decap_8 FILLER_49_430 ();
 sg13g2_decap_8 FILLER_49_437 ();
 sg13g2_decap_8 FILLER_49_444 ();
 sg13g2_decap_8 FILLER_49_451 ();
 sg13g2_decap_8 FILLER_49_458 ();
 sg13g2_decap_8 FILLER_49_465 ();
 sg13g2_decap_8 FILLER_49_472 ();
 sg13g2_decap_8 FILLER_49_479 ();
 sg13g2_decap_8 FILLER_49_486 ();
 sg13g2_decap_8 FILLER_49_493 ();
 sg13g2_decap_8 FILLER_49_500 ();
 sg13g2_decap_8 FILLER_49_507 ();
 sg13g2_decap_8 FILLER_49_514 ();
 sg13g2_decap_8 FILLER_49_521 ();
 sg13g2_decap_8 FILLER_49_528 ();
 sg13g2_decap_8 FILLER_49_535 ();
 sg13g2_decap_8 FILLER_49_542 ();
 sg13g2_decap_8 FILLER_49_549 ();
 sg13g2_decap_8 FILLER_49_556 ();
 sg13g2_decap_8 FILLER_49_563 ();
 sg13g2_decap_8 FILLER_49_570 ();
 sg13g2_decap_8 FILLER_49_577 ();
 sg13g2_decap_8 FILLER_49_584 ();
 sg13g2_decap_8 FILLER_49_591 ();
 sg13g2_decap_8 FILLER_49_598 ();
 sg13g2_decap_8 FILLER_49_605 ();
 sg13g2_decap_8 FILLER_49_612 ();
 sg13g2_decap_8 FILLER_49_619 ();
 sg13g2_decap_8 FILLER_49_626 ();
 sg13g2_decap_8 FILLER_49_633 ();
 sg13g2_decap_8 FILLER_49_640 ();
 sg13g2_decap_8 FILLER_49_647 ();
 sg13g2_decap_8 FILLER_49_654 ();
 sg13g2_decap_8 FILLER_49_661 ();
 sg13g2_decap_8 FILLER_49_668 ();
 sg13g2_decap_8 FILLER_49_675 ();
 sg13g2_decap_8 FILLER_49_682 ();
 sg13g2_decap_8 FILLER_49_689 ();
 sg13g2_decap_8 FILLER_49_696 ();
 sg13g2_decap_8 FILLER_49_703 ();
 sg13g2_decap_8 FILLER_49_710 ();
 sg13g2_decap_8 FILLER_49_717 ();
 sg13g2_decap_8 FILLER_49_724 ();
 sg13g2_decap_8 FILLER_49_731 ();
 sg13g2_decap_8 FILLER_49_738 ();
 sg13g2_decap_8 FILLER_49_745 ();
 sg13g2_decap_8 FILLER_49_752 ();
 sg13g2_decap_8 FILLER_49_759 ();
 sg13g2_decap_8 FILLER_49_766 ();
 sg13g2_decap_8 FILLER_49_773 ();
 sg13g2_decap_8 FILLER_49_780 ();
 sg13g2_decap_8 FILLER_49_787 ();
 sg13g2_decap_8 FILLER_49_794 ();
 sg13g2_decap_8 FILLER_49_801 ();
 sg13g2_decap_8 FILLER_49_808 ();
 sg13g2_decap_8 FILLER_49_815 ();
 sg13g2_decap_8 FILLER_49_822 ();
 sg13g2_decap_8 FILLER_49_829 ();
 sg13g2_decap_8 FILLER_49_836 ();
 sg13g2_decap_8 FILLER_49_843 ();
 sg13g2_decap_8 FILLER_49_850 ();
 sg13g2_decap_8 FILLER_49_857 ();
 sg13g2_decap_8 FILLER_49_864 ();
 sg13g2_decap_8 FILLER_49_871 ();
 sg13g2_decap_8 FILLER_49_878 ();
 sg13g2_decap_8 FILLER_49_885 ();
 sg13g2_decap_8 FILLER_49_892 ();
 sg13g2_decap_8 FILLER_49_899 ();
 sg13g2_decap_8 FILLER_49_906 ();
 sg13g2_decap_8 FILLER_49_913 ();
 sg13g2_decap_8 FILLER_49_920 ();
 sg13g2_decap_8 FILLER_49_927 ();
 sg13g2_decap_8 FILLER_49_934 ();
 sg13g2_decap_8 FILLER_49_941 ();
 sg13g2_decap_8 FILLER_49_948 ();
 sg13g2_decap_8 FILLER_49_955 ();
 sg13g2_decap_8 FILLER_49_962 ();
 sg13g2_decap_8 FILLER_49_969 ();
 sg13g2_decap_8 FILLER_49_976 ();
 sg13g2_decap_8 FILLER_49_983 ();
 sg13g2_decap_8 FILLER_49_990 ();
 sg13g2_decap_8 FILLER_49_997 ();
 sg13g2_decap_8 FILLER_49_1004 ();
 sg13g2_decap_8 FILLER_49_1011 ();
 sg13g2_decap_8 FILLER_49_1018 ();
 sg13g2_decap_4 FILLER_49_1025 ();
 assign uo_out[6] = net33;
 assign uo_out[7] = net34;
endmodule
